//#;; Id7d2c4b2da7a6478426f10a28d9f9eba59a188d1bf2835798742825d32a11125 I8be3365cabaa6a0f90d2e64f03fa78268c135fe0b0758b576b447e9b2068d75d I18a0c098c7fb0098093fc0fd619c8032ae193215c5f695d7f5eaafa28aa64d70 I679eaac16659c013675081e715f7ef761bdd183f1d7f55d079eb46ad6e322ac5 I9ef2faffd23e7fdda264eeeb3114357fcb304142506cbb023c2894ac10f71654
/*Ic3f8d45b35548e4a4ee0b7181f1834df8a2e1aa0eea9b8c77323fcbf46bb42c8*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /I51a1f05af85e342e3c849b47d387086476282d5f50dc240c19216d6edfb1eb5a/I58466ebdd352f801198118e294e38715f864985fd87977f348bfcd7db62e7c76 -I54e67ab9c29a6cfd19408098a96b2a40ede7e06aadcf77336da0dd2b57f25ba7 *I4395dc236d13a1c9b88a791fd2e1275bbb97b927d52e9b8c38248a0d57259aea* *Ic7c59e97212940ba254bbb99e5f908fec3434155e0fbb2f0a3f2ab5a6b4ba2a1* ; If0c929a9e723bc62724e30c7e396e576019dfcb8cfd0a3f264ee5d72e64e49d1 I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.I3485639faf1591f3c16f295198e9389db5b33c949587ec48663597d4e00299d5 -If0c929a9e723bc62724e30c7e396e576019dfcb8cfd0a3f264ee5d72e64e49d1 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.sv > I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv ; Ia8d1cfa1fc63160715eed9e8f5f39538f4520ff839d850162536352ec0a5509c -Ic572272153455b732903e10d0db7356fb56fb5d0a6a9064766547a1304406c33 -I8c2574892063f995fdf756bce07f46c1a5193e54cd52837ed91e32008ccf41ac -I4e1de0094e501762cba645b8d4663534d3eee7dc7d8bc675574f6b130d9f5302 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv -Iacac86c0e609ca906f632b0e2dacccb2b77d22b0621f20ebece1a4835b93f6f0 I8803a3b234be60475d3d6498d388264bbc5edd49f43c780eee4753cddabfe052.1.I04ad2bfad8cbdb3afbf9a26ea1454ac0a07c0eebc856992b38114cdcb5098c47.sv.I836ff184e7b41b1e13cb5fd89fa1de98dbbab99e9d2918913ff43b86a5c7c213

 /*Ic3f8d45b35548e4a4ee0b7181f1834df8a2e1aa0eea9b8c77323fcbf46bb42c8*/

/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 Ib8a92ab2b5e2e68fc63a575fff1d62c25ec6d30209e164d82ec85f5576d9d940 I63985ce3eb57dbe35dec3a2e0dc38ffe14d2e2396edf773bd4f0298ce3ec7eff */

module  sntc_ldpc_decoder#(
// I168413ccee11e827c207105eecf061ecb7d6991383544364fda85556cdf96a57/I373a739f28b569ba97fa09dd5a21185f9bed4792859f1d9cc7fe4af7f6b9c7b7.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 


parameter SUM_NN         = $clog2(NN+1), // 8 : I47c35ffcd3135a74f03fef2155c1874927bc03c22812da0a352f40ca1d7339ea
parameter SUM_MM         = $clog2(MM+1), // 8 : Ifa20411ae2befe271235475378a99513a77cfe0a9614b7cba4d2d92a1f1168c3
parameter LEN            = MM,
parameter SUM_NN_WDTH    = $clog2(SUM_NN+2),
parameter SUM_MM_WDTH    = $clog2(SUM_MM+2),
`include "NR_2_0_4/sntc_LDPC_dec_param.sv"
parameter MAX_SUM_WDTH_LONG = MAX_SUM_WDTH +8 +1,
parameter SUM_LEN= 32
) (

input wire [NN-1:0]                  q0_0,
input wire [NN-1:0]                  q0_1,
output wire [NN-1:0]                 final_y_nr_dec,

input wire [MM-1:0]                  exp_syn,
input wire [MM-1:0]                  cur_syndrome,
input wire [31:0]                    percent_probability_int,


input wire  [SUM_LEN-1:0]            HamDist_sum_mm,
input wire  [SUM_LEN-1:0]            HamDist_loop,
input wire  [SUM_LEN-1:0]            HamDist_loop_max,
input wire  [SUM_LEN-1:0]            HamDist_loop_percentage,

output reg                           converged_loops_ended,
output reg                           converged_pass_fail,

output reg                           HamDist_cntr_inc_converged_valid,

input wire  [SUM_LEN-1:0]            HamDist_iir1,
input wire  [SUM_LEN-1:0]            HamDist_iir2,
input wire  [SUM_LEN-1:0]            HamDist_iir3,

input wire                           start_dec,
input wire                           iter_start_int,
output reg                           hamming_code_calc_out,
/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 Ib8a92ab2b5e2e68fc63a575fff1d62c25ec6d30209e164d82ec85f5576d9d940 I5fedfe54fddcdc5145ac6dd38b4c3dead65f127535af2e07a7b9790515afdb04 */
input wire                           clr,
/* I1e4d9aa7cb1ef438f80454b61c625f0c6aed19675cb2c2f865cbd2e2c3ef2ff7 I2f08a120cf6d1091827fd5d929bad0cbcaa5eff7ae0801098357ed0149cbc06e I5fedfe54fddcdc5145ac6dd38b4c3dead65f127535af2e07a7b9790515afdb04 */
input wire                           rstn,
input wire                           clk

);

wire [NN-1:0]           tmp_bit;
assign final_y_nr_dec = tmp_bit;
`ifdef ENCRYPT
`endif

reg [MAX_SUM_WDTH_LONG-1:0]                  I893355bf7ee2fbac8f9873385982e6b24128db3c9934e37db7bb8b576a4ac41e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb963323153058965c1bb1f6793ee1ed532b856329d971179c54c8172ba1b677;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic1d44b04503cdaccd5821f80e822659de6f6e305c3206e603ef6e23dd3dad3ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I623f2b3e99120e8f406c94a41831d851401dfcedfea86f4b34e5ee38b1273b14;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia02e90fa0c6b93819416a3059cf6adaaee9c396532e724c47648f414a16679b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e72afb03410a9a976620d722e3b11b93681ed53351a88a8fa3590f65bc2843c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43f540ed8151f48307326f27534afca5105989e179c37e992cc8516996b10bd8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8bade7cf8bdd5128caf2415690cff8ade1815c1a93e3d7519333c170fecd364b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d7d9699881b5d4d42cc19d1489f8116cf6f3eef7781b1fdc8cdedda72233a32;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1649cd92dddb73a78816076a829f1c12fb8877cae9ebd080a61259a1d2709c8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b0a3f720c3ed13e66b1c568162495031330a4369a4d0ddf65848c307e1d56e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2fd0a82f26ad0db034e9db0a2904a499de0ae72c5d12f6263aec7a213bf72335;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1927b4579e43362f62245cc1904e0deea9705e4427e3bbaeece21a3e36820df6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45c3eb9c92ff10381f7483843440f1f44e1bceac56ddee98e6bd46c1bd77a1e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia341cb94dc5268759917bc49586f20130d999dbbdcd5f1b34e576770d6d063bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a47b8dba409dae870aa2446c4c554596287cb31f07039a3c01ae78038ffcad9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I34d68a357aa2b44cf3a3b08384498af0e4cc195b0c725a67769d62e36877cb7f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24e4f15f94203d5d70544e5f8b146fcdb89e835acfb8937067299f0b440f7a34;
reg [MAX_SUM_WDTH_LONG-1:0]                  I48a2995df1784de9dc4a3b951d711905f920ed0b9fc0e20ee48f8838a3ba6502;
reg [MAX_SUM_WDTH_LONG-1:0]                  I32519f336568f17bae9f4135fd77eefd67f37ef3c5b6b624521209fc8a69ecdb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45e3ffea730c76c713d1e61276b644a026af54458af4d3894e44c4416f9e4867;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id6f531c71e2af56ad8f4d452827d89b82d866570bface8425648576edf2dc62f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I573b8edf32c67a0863b9e9ecb44ce7154a48ec67472c04821ffcb202bf3b28e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37d72f048ee656b44e4e465e7325741ce519f38a7c033cd596a312d8e12be42b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic2544a607bb965371402190fd2fe4afbd85977e8360b5f0091a6f11f885909c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie51bbbbf8e9ea4467e2c172d3855c3c783c8bc93166f414044020a5f7f45e7c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a641c18ed7edafaa7d5877ae724860b1d54fa6e6890510d1c7febf66944bc55;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id851fac0751063b14367885b08e771c57d9000f29e0e529be1106e6accfe4eb1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7301f67cfc0739e38aae8830e112df2193600d9581476251265730522284b6b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71ea9226d39bea8f66f1c13855318e475eca4a45fbcdfecb5b5bea94e9895019;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41ff59a42cce4bf7225d8f9296ec89aab75a0ec2dc10f0c341c696fc2461ce3a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4211635a82c1f604dfe16daddc0995754675f3d3059ad427ba374cea6f9e36fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I799ec6460c042feab5ece45c8877d0614bfea4ebd97b427e1bd00aaba217c1c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41e027c49a3c7e7075a937c21a58688cd46356ff9a8ecfd497cc216b1d8df456;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf5e207961c05c6ea8ee1cc657aa7bf8a0fd7827e4e550b65cb9cc20925f7536;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic090c90fe7246cfc964e807e465274744fde1c059c1a86c193a553def4295df6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ce1761a25063d6ca639d1aa9094a30899744186121a71229f255eaf3542b80a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I523b27aea266bed319f1eeb7acb39554b6d1129e3c850647d3d0a5f6b4ee87cc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa331e88bb390c67efa83efdb978b28023c3f4a74750928415242eff2a75326a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3585e76d77927b87fa2b357b5f3755404054e391f29839ba9c3a29c0a1084f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e5dd2b4a968c805518feeef59ac29c86d9c06c30446f8966bff4b169c65962a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icdb198ad2d4b3ffc14486474c17026ab6c9129e1783a62dfb7046874dc639667;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9663885f1f636653b6649709c8859bdf9e407c18311f63a0e6677f6671926884;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd4918d774147592104adca1c7b4abe2c20a82553bd5cdbae652d80335fb933a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9e8163c831756fc1d31bf9bb6e966a5c58738673504240801b73891e606845ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic935f15a1c1aa2ee20c06cccdc61d9b18929a70e43e44123bbc51e64bf29e1fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I211a4aa442cd695ebef8bfdd8734fca64e796eec6eaeae0f7c1c306d89ac50ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaaa7217330cfc4c43630903983e580f1ae9eff2fa7200e236b2055614a50531c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e3ac37a60fed64971c398ea5f48490f1a8ba9c0fe63583d4996ef4884aa0eea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76857068f374b6f47eda0c4192e95879ea55667a3d96b78003079f89c096843e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71f710555439b202404f08c784a66fffed0e12c7dad92ced1b83a6f28245a512;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife34f6a36501f7796b3321efdacf37a75e6cb15cc2276751fd20794654b3c515;
reg [MAX_SUM_WDTH_LONG-1:0]                  I458d537d6f291b854051834fc85511253dbd0054f1be7bde7ac2696c4e4424ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic269a154a2e6550cdc5270948790b9962936b7fe59e88379d1fb543fd7f9b8f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e27399b8d9e65418758d9dca1b1cfbcb4d908000611b218f4ad2097da556a51;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb1ef347bc6ea6aaed4c4763221f318e5b5db3997be4a4d107e338cc37e3a4bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38ef2b3fde182cebc6e8265c6e99d08e21e28d55b2eb1b7a161f13e385ac5b72;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d8215327a40c9b967e1a5dc8c9e9c390c37bf87f96114a7d81cd08285223c43;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f2d9a8f6ab682ae8c5fb31b30d5c11be65370398f373fda27a64bf6d718193c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id71a454e9889c6cf7e01d39d50bde9e8bc5850b88ccda4c91eb8266ef7e5a695;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie504e487c65a8cf270fcb907ff7a6f204c5afe50af53c0b0279719522b595c19;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib5228b88950d45370aa8a132d3824bd69b574875b1bd9d3783780b87edbc3ced;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7306fa7f8f192749aacf00bcfc3ee6266ad06e373f4075503bf8c7daa963f7b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2c860739a98a8e6052efa8701d70df89f34952d6249f7266956ad0a6d6701159;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica9704300b0989fb0bb8dd9ddc1807a4906458c6f7f487fb7d7e214e31458eb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I250cee6e4a22b9f9fe50b6acc67a25365520ec326130a11c9c68cce437e6f56f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic8e52a8db0d0cf4d90f46c2d5b5871d31db974cbd84b5e68f4d872ccb6fb9cf5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I805133cb6a397bf027d1985ca36380b66ae7d0b33ca30987f825dba8d803488d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I59ef74fe764da43c107f5eb1c48cc198be3cfce3b3c55e0eac3efe7c9af888a0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71c2e463b98044653ab94090116d3d5093fcaaf7ac48bbe2f5b2b26980af991c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib33fa9a97b26fc69be1d69ad97dcc345c1701bd9ca2fb0922d724237bd2cf8cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  If85b088f394e161ace940e64c404069e394099027a64365e447bebea842a0781;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc1655e6f13d450c6beb85bc81ffd4b765ed49cb361ddcae84e6e635e85513da;
reg [MAX_SUM_WDTH_LONG-1:0]                  I92da904919e10cc11e45847a0102a3b8cc6c52cdc4815d7de7a6c949a2024901;
reg [MAX_SUM_WDTH_LONG-1:0]                  I170b2f3df88d573e89dcd7abd2e33192d1e08eb33a333dab67be7795d2371e04;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3bd78d48b87d258733b0c2d0a166e6921566570e0131a68d8dc65eb28ca4a1c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia554b8c5dc66b7db32a935b99a2e41aa84c6c13fa944f2de90eed8c1d462d023;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3833bf9f2a4fc740f72874fec3b21e205b6fbdaaefca4942cee8751f170d55be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I60e54e7e8d975cee4bf0823ff91ce212f02e407e9e2064ea4ca882ba4961553f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62f9a8d7e8821466e48058b064f25fe8420acaf3a00a1eafc36103bdeded51c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4470cc46d92649aa472f4dce99afb05681b554782384542942fb243099cfc6de;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb8ea528ec3a42384215586669a0abeab4982d73d76a71c72e4c5c45ddb937c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f258a7197af9b66d573a49b5923adec1c8637c53af4c2073805fa31fef73dfe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib9a1b462db35f3d9d512995ddb639c3553c22f5020cc3fe7316a605096d8b8a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I52497162427ed0e9f305f509a79ddbdd02f12eebc337f57d63a9e477ce556e44;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie51c190c3c1827c2c707668d10923b176edee9736a17f532e7ed432af0544083;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d53fc143b190930a55ef8fcf893ea0b45d87abc54330c08bf4b4d5c67d4cbda;
reg [MAX_SUM_WDTH_LONG-1:0]                  I46ef2ced2e09d9ef212937cb037346d3309bba86efe06537a39a963d9debb65d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f819482e0a2454a58a949963a2600e43477da52fcac968f397cade6b69be570;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37b543101174150d8b288848968eb5974a06d0936975538caab590ec97366a1f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I551c9d548f30a033083c22bbd3fb8c0ad11c32fbbf66ccc8d0f6b7a177a49b39;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36fa36e23de34e375c1e39c129c8aa1f63ed250191e4bcc0cddeb9815fc1c717;
reg [MAX_SUM_WDTH_LONG-1:0]                  If00a6af912a327873844b41dfbbcb9b7383e07272e5eb09cdf9b4a4a827b4f1f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0cb9d359df8b98e0323b9bb85a1efa6ba10fd2478777accabfa9e658d8e02dbf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I770b9333cb3aebf6d60d58661bc3282c1fed64de0824268f9f7aaa2dad91efc7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie53bff4851def180b28f22f53a301b0e7c0e897bd637a0045221b0e969249ddf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27a121a528b8c373659d1b04c8b5eaf5856b441ddf1b24331855326f31bfc492;
reg [MAX_SUM_WDTH_LONG-1:0]                  I735d477462d8bc4faf83227feb6433daa37d331e95657535b4e8db091cf9b315;
reg [MAX_SUM_WDTH_LONG-1:0]                  I044870873609a6dc7acef74d59eaea493c553cbcc3eff5b580dfd6a8f176d987;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d907af9ccf3e40047d3c7e02550caa8588212f478714ba92e91482893944968;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1db3917cd01f808a2a2f4c78ef1ed3328ca804093065a1cfb9e15ef210bb8c93;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia588f9a4cffca8b6d433336ac4fdf52e81a27bdbeed8cf2a5d733183c7aa86f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idd38249645258d9f8ef1e5cfbda4f15a700ff3b6d78b9c202bfbeca278528f57;
reg [MAX_SUM_WDTH_LONG-1:0]                  I06e5c848aec73e10515e09f5e32ac2db3c5a972a8084519617121e18c27f4bbb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2757ee84c5d0e87b17c22db78eec37478ff53ed9383587a3afa0e3270afde8f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If809ec52b215e06373de8da5e7b6b16db8490684dab7ae07b39bc7440e19f4bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85ce012ac5bad111ae4ab945035baf1b2820c82822f28a7b7c314515345af8a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc9e721cab51c6460c44a26b6803f4cbd505fd11afe41341e3ec656fe2698779;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89db4b6e1da27586c9fb92f89e492af68c0497029c97adbcdd5e3facac07c213;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b55c5a4fc86bd53678cc688a8577a636d79a0d9b0f515135007234a4a807541;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3bdc9359c749bc85fb3a7fc68446c47edf3565e167d9a28caf4bf5010b95a575;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib378ca85da27dec3042e6f79bfea73ae2f099d548d5ea58fd3bf61c2ff85a4bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09a731c0252003cf8c9e4848c2e8ecb6a86e0bf4d76ed8fe028e3a609d639aaa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1bb76da4e4cc33ffa0f6f61ee985779f4f7a02f8e336f7ee969bf4b4d1599fc7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae3ca8fe4281bb23b5ed7e87317e7aea52a130420731529f44179ea0274a58f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1fb2ff888cbc4ad3ddee50de256240ef2be853fbe54f51092a1bfcf26ed4fcf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38f8f9e2731f858a15a6f2f3a375d0d29634c0da467767e21318213ae7beee7e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia03c4f3191a16f379150692d47660685ffb0b79d91fa4026b8410e2c02219dbb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01eae75c6d18bb06d82fd21bc1aaf1cb883bed514f5497fbc433fdc42d217535;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44aef1d958b6a776898fe8f0f0a8ebc867154b9d4605421433b66f6832c2be1b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5a56b54b520cb4b1b0e5509ed4b3fa804bfc0be8566ed98b455a29b7148d291;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1659da800cada125cbe3b104cf7d512523aa5616f7c9ce70ac7c72fd92403027;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a4b485210baac225fd3f32b36be68140468a6c307f3f91de4416553421e3db5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09149397adf0c3b57e577b66b5b3a58bd1396ade0ab7cb174692b182e52141d5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I172389b084abec531bf617713612fa0d8b27b0967bb62a6514aa873f609bb5b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I15d75a1d3038a54892de000a31379baa7cb9de5538a2823c1e52f64fb061b914;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff3e149eb4ce60c9f28638248c33ab96208976458886b1735785c2dba298121d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21909db4fda5a886100a19a744a9b172b3d171ccd1dddcb5c47b0d3488a48f6e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1bc8f647801308e33369cc5f2652781230a588ae772b1e53992f2124c17ad5d9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I668cba84a2aaea84945a6ebb1a72e6668cebbcec3d78bf88246f3872d78abb2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e3be7e07012df2e0a3bc90dcb0b4756a778cfcf9192e3722191ba8be32e7e14;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2bb5bd1737da6b4feec1bbd2245644956d6e825951368ab22e426f1662650a32;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c01e607e3f3ba8c06fa54e0ea9fdf0dea25c19c9eb317e51a670199ad40ea90;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a26f98f9f83ddae2958fe17b1b3f0d2f7dc64309a438e2fe1f4b8dc87e5d1f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38fa842b13449763b8db07a9f91ab3479670dbc6043c1b363df6c93f6d7011b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifd0ce5d7e19da5ad023cf65265ce2071eacda4cd9553f0823662bc9569ecf872;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie52aeb4c0ba45662d7f71f542630151f22c1801244258b9c8c20dcaed7f1472e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I91855e266ca0be3dab2b079bc241abd61a6724c1eae142ccc58d0a4b46fe2709;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie995e639d0338c10aaafa2dd930d57c74442bbde282aefcedcc9ac3b1eeee565;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a38f537a832431af9ac0e9070decc66ae16f850af8ac9349959011fdbf151f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b7705f03e900fd64d1b68f0b4036e5ef40c39722a2e6bc8ea6f22f91fb4b044;
reg [MAX_SUM_WDTH_LONG-1:0]                  I180662d06f4e8f2216950660d1078c52394ea152dbfff6443f6983f3493caa89;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4656f355712fef190fb3697699fda1c25bbe9f7577a4d1a95aab55550fd7bfbf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5093a95294be69b95d3d4e3cbcd6a93f482b9a77f5214ff42a003cfdb5bc34e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie53b7792c539fa6f2aac95f09dd4a489c9167cf9d6d749f498ab99380c2e694a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If6d7b3ad99d2259ce46cd080637bcf973f36b74bdf7b265d793f04aa27305ce7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie8270cd60cde73d16c5b65134dd393e02f413312f997a0344223cfe05d27985b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I298771c166c7b3809860fdc01e1ee8e865e1c5f2b6a4492af4a9f2dbb6b0e0a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53d82131f37765f57bd586de5a55e92a697f63f20f366913802549f9ce658e68;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2c03e9e66b771798f4ccfe5a9bebd633ac87eb38c9f211f1ce4d10950e5ef91;
reg [MAX_SUM_WDTH_LONG-1:0]                  I289dc39cab39ac30635179b9cd90bd31489a146c8c026138e1a1f9ef7a0ba30c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie15e789de7ea93b8fae0ec21d465a7c42518fee4af3e1f9584e08b3563488c1e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23d6a001aa9c80161e8b305bf34ef8d675247595457a8326a13fd348a02a1539;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6b05d841cdf5f0f96018c49f9a88d21f39875c8f8af17d0dfb16b0d12a670da;
reg [MAX_SUM_WDTH_LONG-1:0]                  I15c69e4ab6a25a44e8cb3ae11dfdf0e1dcf71c2cd63add1ab315e1d8a2d2043f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3c580027dfedf572f89eb6a3ad9f82877baf03f3d6ddba81a8d868dbab61d83;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36dcdce4926fb26d7d1b098549754fdfbc3b61a8947394227deedcb51ef1c374;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9edea5dd63fc137c4ea1044296f48581e5d5fc613cab5f0494a13a6241fa4b38;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic97aaa16a00e936ef8bd742c1c1c14696a72063ec283fcfd02962ffddc327cb5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I468b553f5f3c22cfd36667c1c4f5743c10bc1632ebb3581b3f5151e5f79c6a51;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia28ac0bd59dbf550e8f75ac42fa8618aef3a8323a0e0cd6bc6dccd79c71fe396;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5169c101f3b104ad3312dfa6e081e948c3354bc8a884861269c89dd7f8fe5e7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I70f499bcd8ce706da16f5d06d481e5197fda5d63b024d9850a34bdaf8f41c2cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie88edc9e0f743d11046dfe95865fce6327d2f63bba8fc4911fd93ceba76cb03b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7a936ed864922de2eca56a7a648d209cef422443181f89ebbbd6724f5bd0ee4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae0f73413a2fc8784aa61b30e9699da78e56fd7ba2fd8293e32cbc9dfe6bc114;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa54fad7897ca3a5db0d7fdf35cba73823e245f86c54af8a772f1d30f540247c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I68165edd77863351062c8e0a09c1efdd3d244841d10f66ed22b25236c10b84ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8c7c890f6f561a9a81130bf7ef4100851c3d86620903cb6b6d648746c0463b46;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6f3393df8a2c258b1c44d7ae93b7b9ebe39c27cecee6bc2acd3f5c191278d2ea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53795a7f407f9dd9d22f6483bbf9efb36313825abbc84c49e1885b01cb2724ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6189724f652320ab2c3d18de4f35ada1ebff4b32b2d3e86c66a3f2c74941172e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d28182f6270a0cad620a562c047b449c03bc2036e855d1842707337fbf007eb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib32260d6129253637588b8358e00892c493347f945a010d24fe897e6a9f2eae3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2837d4f41e5abdb0abe8c9282938afdd85015263ad60e9a187ee91944f18bd1a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idce2a9ec74e8909d7514e546c058c4adcd18ae2607f3490cc9918249ce38ceb4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I832e0057c56a4b0624a8ba7fc95565ff1322ef3b377d21b243c1fa69a9b83982;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8a985708ccedac94fd8d239571a6d5a2fe336ece2d15ee7d0abe9a79dc1e48c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81243c0fe8b8a3ab03ea4a07b48ae230b9783bc2b49006705893387b2eb0353b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic0ccbd30732da760b3a4fcf87c08c87c22cbf26d0cd50785f80ddd7682b1fdce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53e079434705c9ad3bf3e5cdf3f1d09bd1b0f7742fab2145a089e823e5c28f30;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6d7c4898670ee6aa4eb6fd97e1abacb7e4152c19d5e286e110420d2083a5412a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I77f3f1abf296aafc631f7b3d8bec79228071d4097f2083f70dfee8fa6ca52ba9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I48ec069746bb9dc6300ac6cacbcc382506e2c77773451d32f4d9fe4cdb43ba8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1704967bdd23aca028c7fd652f9a0efcc55a31662c9f9b65911b7c1241205d9c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94f08b3dab411dca5351bddf1de6f5e659685e48a5ef632fd7d4e52dc69d3dda;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia2313572dea3f44e7ec31d1474ed481064164548d3de394b69a6e99f60561388;
reg [MAX_SUM_WDTH_LONG-1:0]                  I80e179604c153f8ad75c1e75837fbd86beec291776ff5363e2302f962998776e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb8aee17be074ffae08bde14b025127c77773cdf482aa5fade629781c3488e18;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8608849b8538dae3f311153c3c70f026f5bce23c17237d20d192c838f0d890cc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b2da3ec326ef0ce2bd1ef54c04f06bb0c9c7fe6f0736613537206d5f5568ff9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I530532adc42fb00f7f781e6b1d108a4d2444cddb08da7c6d088ae9f3d6b7f265;
reg [MAX_SUM_WDTH_LONG-1:0]                  I475e873205aaae01975a2852b3d3d99aeb7ec9aa17759595012bf55fea91ff81;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia75f7e68c65cb713bde41f32c61fd9b320c8f4474fa8ce88598372c0fe14c930;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d7892388f5775db1b77de0b60b10ed4f40c44774e1ca7ffc723e5fad503c487;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icca7f4c8f454e356434907ebb02b97ee9f5bc1e7cf4860adb16a1dd6a6b709bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib459acc97fee8ddd325d7d8b18d5c339a3c1e03c919c750f88070ec8a4f8a0ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4214214ad8fd0512cbc2cdfcd1f1d11139d4a44c71628c5d2c1f00193b2dc777;
reg [MAX_SUM_WDTH_LONG-1:0]                  I25711c9c95cd06f19d25d01854fdb8290f4759c9133d1a0c9e88548b886050a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3151a9171bac0e6e2edf837e6bca27cffc3df8c9971c3b3a6873cd8169f34fda;
reg [MAX_SUM_WDTH_LONG-1:0]                  If9e2ce38db8f4cb30a3748fc7ee1244c98a4ef3c6dc840123405c585f6a867b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8249d9d116a929e5f3c900c84a36d456b162f7fcd71949c88fce1e080cdb72b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6b1a6a399505ffa0312c9c79ecca8d63de6c5a1c9f6c0590296cb316c22d114f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibce79851c8253df32d60965921c117f70bdd9b486aa72bb17bc3ad578bdee995;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5454f64581fced198aa8ed832feea4c5a3de221d45b8eb42ae5820d82e540931;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6a9121933f24798dc7d6c4671e05f959e4514a894f78f0e6ca37a9cfc0f7a53e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2235e43965f0eebff14c5c279ef56fc3e4055cc263c20f8d993756e7a5d9b2d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iab3c6e4766bca2055b7c11e462f459c0c69c45c76b11fd6aefe62006c7a1316d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72979b4880af333f9e67500779c23973ada097a3cd1e2d4dff0eed1c570f299f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib645fc54982c8fb5921b1dcc8ec4737c61a564e50d7195d4d9214b231fa4496e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d0c6d6a69f818fe0856050283b987099cd8c7f3c8c22fdc825a01734c4642bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7e0e378e8448fc365285c0651e01f06536e3adae7e9c95f309e7d9980d5035d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I811e21f3227b2bc3bd72e9b312edf9bf8e88261543c6bdb1bb09607f49b8206d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia325319a3b0f63d7d994b0e5ac83b8cab618c9f79ba7f60dfc0c32bb80c5c72c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e06a2f339c14dfd77c1d58f78598240d08a7fc156a785a8a3fcae2d2d6d0549;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2da0a6fb45c46249fce53133b82906b2668976ad484cce849bf7530b5c0420ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I167bb55e57f960522bce657a28f3a58bb6d82aec339cd46a3e8c4136ee023474;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e4f3c6c98d527ad3075a00ecc95decfa07785b7b0c5ff523ae53741ffe019b8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifde56fe010824d9eea62caa160db5bde8de47e31630cd6a8c5e0572df0fa0709;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4fb260b26ed5bd044dca51e17dc1b4a7902157d61ba92c823b47e375f9944bc0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b81ea9b142b222ca4b90724e3c4facaba82a4dea5c9b05c66032b06a459706e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e94b3f49feae361294ef10579f5ddf4cd4e7656029492a1598cd5cb01a85887;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e9361e7d30732f3e689391f56f9007c32c2368c9eb9d85b933f798babb0da68;
reg [MAX_SUM_WDTH_LONG-1:0]                  I54c78cf957f6d08b1ef46a35ec24b04b3400321d670b4137d64e89399cd3c370;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1774935be7ae799801f3b949e3a99707c4b32e7b1538e9f63cd8b940295ea6b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifcc80d9233cbe913ec2813cdf22e5da4f6a463f224ce7db93884c3b49e6a7a97;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia4f0bde88d8ea45e325a92c25209a97269d31e2e3999ffe83696236b611de74d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I30472f7544755b800fab38e17aa914eca481774221aa925e5fc526aa7431c05b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I30378eb921b9521d10fa2953f99f0f362b986bac12404a78a5f50619fe3b55fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2968bd466e64c0ebce5448acf7247671f5f669f88bff8cf1ed20b47e29a9f1f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I972ff0b38d85487454c289292e792035f568f072c33914f87e1f9c981da34370;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23dc7c83c84d15f94edcdac20ae49442bfe44709dffec43950a95b107b0521a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22ad40f4d98f11e2fc7b9a8d56e44092f6e319c4edb2a67c5d9dcacb6a038846;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40480c0b76e0574c82a8375bf6c3c255f6cd5e8d9f3c09c5ddcdae498d43e294;
reg [MAX_SUM_WDTH_LONG-1:0]                  If52bfa5da5e6508360b34b20a9607809dc732ad7d40860c8677bb6983d8c30a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idaf0d98b59e58bf2225f5790830f4162cfa3dc258f0bb9f84e81d33e2e2b097e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e9200c7443fa92d38415a8988c0a7ae2366612db06cfc84d9de4faf53d7d1c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia9202e23aadf215e5e8887fbe86fd5af4410c49d5dcd48ad38664a63e4a52a77;
reg [MAX_SUM_WDTH_LONG-1:0]                  If23a3c0642ef8cb4b2d375a21de5253ad97342b92d29b8b7417bbd9ad0fb2fd5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I911a22b33617a35907440f195ef34301e1abaef90df3cf6b455b7aab22aa7637;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b801d7872264ef55cc09008ded93c39bcf86fcd83e472ebc91d27c953520017;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8aceeead21c39681b7587f543140d493989947711214df2082211fddbe4467b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I727fdffb518b29e800d3761e94d33c96bf32b4006f248d8eeeb18a035a7c8abe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4a9ca51fe9e7ed20f97438fa441c48b74f2520d29c3c6f530f1317d014a4a09c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b5a25e13e61b54b754dbb201add03176d432d0c31f3ee1a4086797eec57cbd4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84b6567e6638ffe91637cb5c900fb87d964738c80c7a2bc3c02839e44c665bf8;
reg [MAX_SUM_WDTH_LONG-1:0]                  If4413af8c4f8f3dd1f90f00fb5067c95a240f9e3ba7271b134cfda0a1fad603b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8507dfdc1822c3c555877de0a703babb888342a1cd4a5345593c0eb99d72f5c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0640e35183fc639f884fbb98626d0d54556ba20b2a709c1b4eedad0d3e27ad12;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8bb5f8d242836821aa26e984a13318a5e507c6bca8479e9c2e3ef96bf24350b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79f29e0d9e4930c0e8eab1a5fa373778c2663402943ae843e94dc1d3ac60192a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic21b3ee91f7fd6945933b2d6aa6a8136c92b40340e6ce286cc5f592b6d585a1d;
reg [MAX_SUM_WDTH_LONG-1:0]                  If41e7a25c141c9a83ddd7dbf5bcbb72f579ba7d25231b25ab91ecdd1b8c50af0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41e581525a6f6f7decc5d6b1fb34553b16517fa79fe019d523dc0de19975dab0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iabb9a156ffea98c56dcbde6d29fd606deeb21debc4aa2629e41c035547d5a589;
reg [MAX_SUM_WDTH_LONG-1:0]                  I154a0c43cc16258a8b281935bb29839d099e65ee46bc98787be8aecdef9922e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I496dabb1a4608940824606478478a3050517d422cfb20c53c37523f34aa08a45;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifbd920d2032ef4cd599ba64059574352b60ae0734a6cbed208f65e8c04ab2efc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8bf71b880aa8654933f2008a17308e8366b6f6f22f52091e06364bd10004b891;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b8c17efb60e592f131daf550ffa3dc4a692cc5892ce1bc726f9024a5a714bb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1748e381924bfb743c1257d7830da580af261ef967ffdc1adfafee17c67693aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I12b9fcdf2336d8a724bb7131ee096233b51a61fb5150f5a622509303bf56d9ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7412e7d6cab6a1cdead2bfb425b79f89328cf155ce5e3b7e8593a4abc457d4aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3f507c6e543114ff388cd6b8eaa2ae808c46166e2b8badbadb1eaa37f0c04d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39fc2e50c10ec72f5df6ea43b36d62fae7c1c3cbf6f54e921133adc9d8ca884f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f46d67075a762da1edcdfcd9fecf3975109a4cc488f66687f81441a821bbabc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3be1c01d32bc2fd127d4c4b371fc566b3977bf6f5ecaf4fb7f662f7bdcb36ae;
reg [MAX_SUM_WDTH_LONG-1:0]                  I02c96d25df89a3bbd36a7aec220bc13566ead49f7fa02b64b96d46bb7cf8541a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic9bd71f61271b1ff2f37d36580487d70287b498a51770475819cbfe50d3e48e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I615191537e8873d55c3af429ce9e1019bda129cab124ff2dd1ca60465f185faa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5217a6046ea279ff9f6f40af49af30f0cdeb374e8c2543da9bb27ce89b08044a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33a3c95ff1b26a9158939189358494e93f924d9b8bc3a4032bbc53d5b7b241d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8c201e2467b255d627059eb66fab4ef48d0c235488dc0f7eb7c350a1d39467e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d8024a69b10baaf37cb9911eb275f1a827b75cc590c9830cfa90f1892ab1a87;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89de4a293c5da110f92bc9aa9b6ecc790b2fb3e1d282a6373d5ddaff63ef6518;
reg [MAX_SUM_WDTH_LONG-1:0]                  If683ab5a719cfcc8aea312c7be75e5fd3e2dae0d517ee14a136b1181209760cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66a3806824b2190f9af7e907d1b4e068fa12560233a9a67bcfc8835373d6d78e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3f9871ea280c6b53533e62c3927542a4c4dd28ff2c551ecd1166b9775315390;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia7af92f6f7d9e7629ea5a0dc73f90acb4cb2dd8694485491a528df10a2b00aea;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie07ac76b3131e7a779a284315a5adf27af7b970781350c076b5f5b6d74e7a45a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia0e8b0cadc0431f58baf6bd1e0fc4ea9babaadf97f47eea75ce07e41cd0e8822;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia9746cf96c8460169eb7c522565deb2322a9984aecdc1473193f1cf0ed5542b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c3df19631206eafab24135f4eff9ad9449c874e02c4fa9770d4fc4ede66b3f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4fb36b8d1dfb44eaa85b9445f8966900fcbe3e895daeb0451d5e23b9df6676de;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74ae8440b495f97712924217bb791b022bbfc59b228632b7f96649f2a2fa053e;
reg [MAX_SUM_WDTH_LONG-1:0]                  If922d63aac5ca5dafe88f6470303e1e0ba23c90de33d4bdc8432a3c81dae9fb9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia9c79734a6daa19386ecd68dad6da50274ac40a694cfd496dc40736cb4b33da7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I759f10838f0b7e3f75c8762cedfbc1cadbd61af8f7ab3a9e7d88bacde6dc9c40;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8d71dedf25220f16c883b67bc750a6e3c8886a6238f13693a22b41345296b0b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7541dae782ef8b038f2768096ba4fff06fa9fcc6bcb72ccd9b8fe5768ea28941;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieaea96e9413e940b5858f87f12dd18ef7c88b6e84caea900505a50fe657e21e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia13360e2c05d42edd07ecca114d163efa53ef77481588add80343fce0a426d24;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic8d159cee07bee92aa9171ca69177796c91fa7542a63970a29d785b3cac2f30c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I611d21feb8ebaeec639386a89b1cf2bf5144303d16d80b557265f9c66a00c1d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4aee30afbdf3dfb74a29ea9bc15aa1b0d200331984b528fade3be76c3249e3f3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b59fa34c611ba64fd61ffd1ba77f01508c0122f8e8b2e2aeeee753603349e2b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib48fdf999d6a37fee27e903a4581bf51bd4307f83a7a18c3d7fd5ff5e8490a4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4f44a415623a311f037559bed8d19a2cd306a1b12af2f9d015adbe009152908f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie581e7d5885d31995c15b699ff1c7f397dd32496d88a5a4c77d1c5bcda532212;
reg [MAX_SUM_WDTH_LONG-1:0]                  I65abc9fbfc8e631136259f0a5f47d007c810303995e55de1e7e9f7ccde035fad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I317cbed94b414a879715617065e78d4ac271816f7f331e5545ba55a46bcd9a5b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1f898aceb1ec1cc51f6b9f99e3f9d813eca57d9642b5e41ddf6175c6abe7740d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76b80ce969069fa14c6d7022d6c072434dfaed48bb2b30aae77035d134019afb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e2ec7ed430c3dc4cd717cc7a6961e5e7c636d451837ee16a456a1d04d6247cf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I732d56627c4f920af6fac9e623551f6c4c0e5e970b37e4d2f3b0dbc0d2491e29;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib9ff76d8c63a43b6873b5f305c93676bcd412530b04ebe4afbbbaa27a6b8f25c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c758d1653b4abf515df4c565803d4d5130fad01c8b46a5d447571d0fde55bb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3b55be9a317757f5c0144759a5adf67c44a5bb4afe4e60ebeb3be4ec94b1fc0;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8ee177b4825244aa2459f76ce3cfe5435b03e72d750c440474a42fee5009643;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3e25c67909179600ab8e63f0335fdb849cf0166472fb983fefe68e9f4f9df7f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibbffe343259cc28309085b16cf40fb046a0a7c9d5dcef49182ab8ba0a9acbb2a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iabafc2aaab132f1976385bb8e128f51ff86417dd26b96e57df8e56a2b7044d33;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ab2cbc5eeb87f6f79360ad8b27bcdf5daad4c85f829eaa00ed855099653be55;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic6492e40db63085730ca2ab4612ce1d9b385e004b467ac433bd9dee4b81990bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib928fe4e8b8da0fa26516833082019238c839091b1fb32c244e57a2aac417273;
reg [MAX_SUM_WDTH_LONG-1:0]                  I697243100d9508441bb98b0849280bf0d47509aa42f7f334968a19113ea5091b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib59d2666a9c62eea256e01a7e240af2a1c11a86a51058e6ed4034007a881acf1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b4daf5f5619a17e4bb744ddd92d5bb1a30a01e2928a200d796dfdb9f7594c1e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0eccf85cb5b32056038d4f13293549f535d994925067f49a8f1abb6253ed45be;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2534e75a32847d1999b520266575471effb319ae660aef5e38d0aaac66f83a8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c11c8d23929c41fd11d326b4535976b5e6ad33e2969128e4ec4ccfb0897a22c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc4f182435db6e718a7fde25165e26678a904f8d7372ecfcdacfff50c99c0f79;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c9db5ef7c22e9722e1811495675725bc9367c52f47417ac0127b2ece6c2b6d5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4927222cb1738667a383028851b08d20223cac5a89a663b6b443bb2ee77263a6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d113258d0831ee2590c286fb25bc418e5c1d0033cfa04428717bc3782db11a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1c743f39e92313845da6e20dafefce9dd80e43c11314962f5fba867c037687b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37fbc80705b247541af9b0468d3bb960bd4b8c1908084a570dc6435714c0f2eb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I580cb70e24ddeade0ded45cff406069ff648af95813a3d1ffe82fe9916894680;
reg [MAX_SUM_WDTH_LONG-1:0]                  I04ca88712e988bdef397bb8c4e680b6709f92094d54013e6d786aa459174baf5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id402959580cf99cd1d64f703a31be57b6a1b1eb883b8197096068729df11b293;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie8303e1d3cd1305166144c2a9c72da17dc5ff4c6afdb56ea458d2c017a90fcac;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e19af5e5f4b25b16be3d56eb0b7bd5261c3ca95a38576983db444d6655809a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c8296a684c3ac2e51841b13d88cf64656b4d2f7ac1625a77e0cbed908eb5f8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I87b00103000c17b5d537b5f7fb82eee037c57dc6b6a3a4cd43a19a92efd8b213;
reg [MAX_SUM_WDTH_LONG-1:0]                  I70b00c7b7fd70b24b225260cda2515d3d5df30d630e9fab4b9f85d810f441649;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57ee78ee192d7bc07ed64d3d42bbf209e954cb023f7725e15482335cbcf402a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I891eaf9692501bbe1df2bd2f2470be83664f12d9e6211b5523bd7500a1e9fc70;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibba300f2463e7761c495190751b83704f8a828f727ae23b274c153bd605c758e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I807e8a0a095e42d08f8682b77d262989f5440738b49f26eda30b3e70efc7a8e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I302b994f71bced52060f5016280bade3df63be8e6348e8137dbf09ea339b2ce0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24a328d80a0dd14fa15ad6101cafcef8008c5846474fcd62cfde858dd3d75461;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icdf358bc87f821358185d6b64ed28411a009602f1bf397ff98dee49cb851087a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8273973db378daf42a5ba6dc50c960e8433a2dcb5d17c30f95be6bf89ec0f0b8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia74859916985880396078b181652782883d5e69db172af2bd6b5abf5ca55da72;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7ecba0b25a70555c9243a99717462e9f43cacafcbb2ce9b03d34054858620493;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76b090fba89f431fd007a510b3d1be2527c10360521dfe032cb18928fe5e5e2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied4b1e4e915dc6bf15ce0f505d7ac9fa6c5b8cbcc5831cdf270791ea45402c8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie19a52435cba71b7b88711d46eb5d530a9f236e6a6a2a19c9213d0b527e90719;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b2b4121708eceb760e2854c76289daff432118cee2479045dcbd8ebe358e3cc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7541dea08da40dee1671fed651faf2225a9205f04627982312ea6d8eb94ae3db;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8eba7f46df1f21311e46e2657b38d61800060add0c96dccfa9c45fae66711d7d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I879436c6762d7a1f92f45aa9d70bcc63e0ca0957f69d2bd417c5a4410f4b24c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I587e2742d73f804efba3b90efacfca020ee8a5e13c2a490ec60ac494be39a275;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1c46edefc42352d5d7c429376d363db5a76ce8d5ddcc76e2da909f07c270a48e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4766de4b982a051c7546be035a94bb07bc822061d5bd46d9a4070d026b7a593;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icbda121f4b7c783c142a1034a6b893200c3a974ca08b153ee0ecd6baadd03099;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5ce28b3e49d61224902a9c1f675a4032351731bd0d14cf3bcab007b30d7e5c22;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib7a3b0d88758dcc368ea5aa65eb4c638502d363b70ebb303394e701e588d2a82;
reg [MAX_SUM_WDTH_LONG-1:0]                  I07afa69acae532add7b503ba1bf357b95ab120399bc63d32e65af6f61a369f15;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idd87b9bea69d81d0c6e4a3901c764fbae4fc8b0795bae1176b2f5b75ce571d04;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4c0f888abd9ba96ae660c5a3f6e9c627c5775611d7a2956fa3049c5574fde7df;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifda52cd13144d30d66a9a0fb8b6c68ceee044c33751a0f3864b564eff21bf815;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4bb74c7a5d5fa7f8a3bcc33e4aac51ace977350ac258b3af687b215c37407b49;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee4a4722007fd835cf2b8e7b244a8f72fd79b0f418fae3ef31a50b35769a3b0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia781a129677ad67c301dedf105bd58147a815283dd2c06d65ca7ada0aca7cc7e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97604434d22669367d9ace3fdacecd4f777dc9759b5940d5cff195fcb0881346;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieff7f5ac404485dc7719d026c898a08cddf9eac3289347c09da180a04400da13;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0c6a201e2d38ed7791d229f2df4ce0605197b5edb176ffd5369d85764de153a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idbea312fceb0d3b89f626dc27620dc564adf927f2587857f0c80926c0f323433;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69f0a9020d4480b3ab0eb58ec235ffa667587b7da910b3854f56cb49e9047d47;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1537778668b48b3115e7b1a3cde430a348b515e592a110c520b33226ecf7f47;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c2b1197b3d0c6879b675bf90f26c3a5ebd1cdfbf6f5eafc502ad622535df53e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d749601335050fe4f61b7b9280c1f83ae58f99216ee191f039f6b94b185e74c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I576f9c047b4db49719b8ef7ff32de3de609df2969827ec22e91d8b1c929abd99;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2a445ed5096a1929dc2ef74b28f3243c9e05c70b4e0aed9baedfe94c28d8e4ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22d7ba6fcb1a3830055bf29a53984fbb01f70b4f9c309f6dbf0a2cb493f39818;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae58883a74ef0111e20be8cc9df222d4e0e213d390b08244a5361328ba38895f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I16e5e8ec4564f64f3db568b15f064d343674e523b9f6ac2ffcdc1e64a3dcac44;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd5a78278d93327ec1527d2329cb8bdc601611fa5ee53fc37e64259d6bc217a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I240e73cf6faba62b6fd94d95cc67aa7703cc8e96875b5dab437e79e7a384ccf3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1f021d678d21318bd8881474b337f0b540c16dc97a33c4fc3abc12bb662f4a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c8e8025305283334b1155f2e020f3909d725f3d656a9209f357f396b345bf9a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id4d52f3a7303153d65a86d328d1e7e5dcdd602d284aba3e104ee0528d9b1d465;
reg [MAX_SUM_WDTH_LONG-1:0]                  I236740a734448318d6759a5e14178c1bfe93f1d1f793768577105ac5ee42d6f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I608fc1c1a500a0fd76e9a326afc6c5a26d1cd78f1b150d970f5ca74d1d7a3193;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4200e2460844e967c243fdd9ea3e3863aca3b8023d85311149c7b30e2d3ccc10;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7b2d4fe3f2c703eace8068da2810bc7bc190900ec3959bfc4a396e72ef5a8200;
reg [MAX_SUM_WDTH_LONG-1:0]                  I831a730b580c0d83322ab8cd6cf78e490b8e104fac72df3a67d75d029a18178e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72d8c9fea747adec725ada83bdebc85126870df2cd2cb9f88d2d043635bfdd84;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib33753185ecae290a3ff7193c21cb9f11014cd9ab59194b625bd9fb1ddf99413;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4f237165ee7800d1fd20968d90afd5a858b8ae73675c1a03b67be17159247ffa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I780dd1faa05c0ff00db1b222da69e706fa7d30b9522b0ec2b89f6b23c30366da;
reg [MAX_SUM_WDTH_LONG-1:0]                  I333abb8de54c2cdc50519fe091024d9862592e0191ef4acb0b6e1b7c45701234;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9cdd258f7d667c4be0a7f3eb13f79628e9bc1c12c8cd9febace271ff54191872;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ef7e70fed5f181598201b2c2c0002f1251010c752be38c1f229c337e4a66428;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5996255101f1029eab99365af8b51d34cd6ab7e8d3bdf19598c43c5fa910d513;
reg [MAX_SUM_WDTH_LONG-1:0]                  I75665f397a59da51376855f9b737164887c48da916cdadc4b4d1605f3d8e4071;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibfece5f844143052755772dc83b99eb3b78ef024232c0d1c1ca251da508d3516;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie81e5c2a20cacfd646fdc8795e265386030f32624e917b5877a38d9790ed93be;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3368641096566227d03c6778a2f243fdb3b21b67dc940542c24f4045931684a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9760a21471e149d0c56a22ba9a49f377439bba25562cdba484b355531562bd05;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ecfa55d807d1228b72f0ad1afd67133387e87cfa537cf8a7619fb887e86aaf4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9ad099032e87edfcc146b2b8fc401eb78cd1c370d99a7d87b96cffcb2bace7f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieab494ba47e97c3d84f264bf6017276cb149db18ad24479caadf0c8d24ec487c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I42d22931f7defa6032679880bb907c668d62e4c65343d359f7ee0679bb098ef2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief87170e911c48a4f8f1830ae52e6b34421df444bced0e8746e004999ff5f39f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d35fcce50496260be81878d7799638cbce05d2afe98817fe9c53a675ee5f98d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia1e1fad227b8e563997b52484713aec367521484f20e560a7dcb2780bf2e39b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0876112eaaac7d4bd5dda75039d334a15e6d500f29e0c471e8d6dd0ba6cf70e9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb4e9f7ca3ef03a86dc723495293aaa4ef9783f92a3b05b3344ec8468f9675dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I612926c7fd5a7811c91d55336a1ea5a427e4c28826227d05d2e08d501bb032d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I677395b9f313591599a7200d68572fa3eb1b30aa5a4bc4476ddd9fd840f29edb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4075a88832d68ad5005c73387153538516b97eb30d8d1bfc9f3d205cf338e042;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6001c8b3acc2e47f7beeda5c633fb76e0f191d6dce473637683c7f6efe4d3b7f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4471c46046bb6606ad97bff8b36a4a9c1643c861791e8b3bf97a41e8cb385220;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieff52577c0d3fdfd35282159bf2ce744dc12f879d290abdd6f38a0f8b5241dfe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee30715a934f261b8e1fb4814e196f3307e095ec0dbfcb10ac1fcaa1d1d16372;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9bbf9a8a49255908ad3f62b8c4a149837fde63060eaa2d01bb382fcf59e9edb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8b323499e4c61f57b164a287da64b2f1c933376dc7ec202d666ce57ccffc139f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ae8a856ac9eb44659cef37d3140bcef8b5253afff93a2b3e54eec5c88b6ebd6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic936076da3dcc6a7f335b0d3b428e8b01cfeb9240df6dd50bcfb2188cc37ae8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac850cacadce02a577a7ae8d4d48b52f43aeb883994730d170d89c9f6255c4af;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1cbbfb485fecaa90d26f81a89b89c0d778558fbc218268369c32c33117c33468;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic680429748da0cb695397674fbfe3bbd5f2b5496795b05051d9a62e0c7b38884;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5bd88b9b16b4fbeeecae426d343179b982f46fe09abc37e1db23e03a43157b89;
reg [MAX_SUM_WDTH_LONG-1:0]                  I617715b25070e943cf4b34892f49447ccca1e24e4182820b36e87194ca7edc1c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5fcf505c93f7902d4ed6f1877bf51599e910bbcc6002e122623c389e72e2600;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1eabd1ad44c5bacd15cba04670f5077da1ea3950e797f2ad5bfba62060a161a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2ed8f97504f1f2331d11107b05d538282eba6248d7d8fc3c9ccbb4a0cfd7e70;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd5dbd51229b1ffb3fbc33d4567e89a5b5767d759821c0b4761e8b1cba3fd021;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia2d0125fd752a306fa45115b7d888f2eb705d6f14d3e5d4f5191024ed7b1f746;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib59b40982a0fa0730bd4bc1b740c68166cd0db83909258e2d0db220140f7ade9;
reg [MAX_SUM_WDTH_LONG-1:0]                  If45da818944a7fc1d4baf55234b4a8299f0513f6db7e1e8cd87e7b57f72eb817;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3a3d8a238fcc1d5703240350b6f311213ce4d203c859b54a8ddfbc6af08e9a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I18d435d55c2e6ef05cdc85c7c5f1fc2e74307ca98333e485f5fcb8eb038dc3f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie1a01aa1296ed81d5b75478aa0ff85cd0866be9418bb8d44d257087fa4f6b345;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6b9155f4e226a633f272039c862d58cbce7e31a597a37e1be49eb81b0b72cf47;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01eaac160521c659f8be7398b4b66d448fdd6958d181bc148938a1aa3e3fd350;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7dce49639675176aa767ea6d5b2171e0c72deebe4e007b620860a1f8b177060;
reg [MAX_SUM_WDTH_LONG-1:0]                  I28e7f4c19cd1f47169d939f8c94bceb96e0801b0a66dad9dcb1d2c3a1e656d34;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8043c8446ed3aac742a14c3df20420bdd5f0e6561e15c32f4045e2ce8b6f3330;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic97e339e12a03eae013d5cd740b137561bde6188c1c9b31f5d39199bcf287b23;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb807bb8e9746d06de25556b579e51494e760b3a4312caa4862cbf2776acbccb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie83bcb1fe72e7583b427cb92e77a596a158312c89c2ddda3ca5ac113f7e8e58b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie1f84176002d4791b93729913c6021f1ffd76c58ad11593dc088cbcf2e4bc4c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e634f64bc4def7608286b21abd3f531fd18233e92626d134a8b986175008c38;
reg [MAX_SUM_WDTH_LONG-1:0]                  If56795023544f4a2942b0910b389ee77a220fffaf45786cb20c1806f3d76f76a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a3f32d46730431a4e8b755f34e45c99a2498f70b0a1a72e30247dc78e20e944;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic9d92acd0f4cc0aa5cf4bc5a5f14bb848cb4267dd6aec78011f70039bf4f7c8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ed20cd620c713a5aca6cc3a4b55daed825a10b3f9d779e6e83f4073130a5528;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83b87ecce5b21302ac79a58afdd995b617634440666c2a50df5ba1868c7f81c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I815ea11848fc8d4e5819cc19e041d9053b9f67a76ed786264b86c6d92c97464f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida44179080ae7121a94fa6ddc8d15e57d73d73f15c2007f200eb205bd6c0c63f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id78afeca7f85a7fd2eb3cbc54a726ab58c640d233f3b1f54a728f64ea1038fa2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0708b20a51af5c02051540c2de37aeeca5959bd958280e953a9cdf18c324d905;
reg [MAX_SUM_WDTH_LONG-1:0]                  I366b27c864334c4667735336cb00a70a99147206b5b080a90f7c73d36ff24f79;
reg [MAX_SUM_WDTH_LONG-1:0]                  I25510ca31a420de3078e0615a3a9f602e7a6f8698e6a79cb0d2688aa63f8e7cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36793dfe7c63681d4c68b218eaed75db71f018b3b9a1902c95a586f9a040e60f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief493235efee1fdb4705ae4a1a0244c57346ff2b56b269552c6b5d64595056ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f23f925a53b7246e36a09e80472df08b155e259db2d0ced8963692d36f85c84;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a5ffd7c103836e4867f6819fab3096c582f2ce1db2c303bfebf50104b7d496b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45bd49dc6c406523eda6bab5c72af5615d2a052f7f43502665d95c616383950c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife97a26fdf22e53aaf139436dd732d1fc8cd6cb4957269b6d0666495a0873c4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I17013aa37e8e70e1e6cee9d90e8a3d4b07b1ff9122b2ad8c3b4c99deab9e6952;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2bb55e3fbb0c342fd0434fbb00b85eae3c5f4075979e290f3d22673c392e3a60;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7506221ee4a6d544aac3f4da89b28ab6fa9d4ea68075210db51d8c6c0d486af0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7dbeb05d89d3fea39368b48237973c682e796d24aba3438109147cc316b96ba2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc7ef4ff5d5e894f81ff8cd7b641624a6a898281185b77a1e2ecaa556312dba6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e863b3eb7ba8e7ad90945ec76c695330de32ae32b69ae2a03091d1ef0142670;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94f547c68a6f0daca7dd1152b5c9440fb76b34a3a133c8947cf8e1ec151cf3cc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib13a4de6ca8fc3856fdeaa543ff8aae727f62ebff652acce5e23c6c121ee740a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I80b8de6095d16eb257b9da8adcb999d08ca7412d77b70d50bbf75ad9ceb0ee02;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22692863c63315b86c8a72a902c88573f4af6aa3b1691f68ed588a38ac77f7c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife51a94dad3ebb020992018db5c1e1884eef8a8afa5487a3365594fdabcda2e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f18a4d6ae6bbfa53e26a0aa169b1cd1c40ff544f7fd42b9ac493729ffa90ce3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I71fe587ddc1cfb6d7ddd3b8471786134d761d3987128e249992f460a0fabf1a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c4daf848487e7de6d8f95704179a300218ae460e56dbe71d33805739ea61144;
reg [MAX_SUM_WDTH_LONG-1:0]                  I693f23e6d443e1a19036a40851f82c92837e7bc1db7efa4913fd4f4354e88471;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94386cfbe9c6f26a678c961cdb0f15d314fc3e6bd04edc61d5596107adc68969;
reg [MAX_SUM_WDTH_LONG-1:0]                  I43594a967fc4ae5970a0ea8821dc6b91e5de451cd6a5bee90fe8be18dd172caf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icbf8ff1f03b79fbbdd3d73ba2d399ba98a814ca4db6f6541ce67d8e5558d0eb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62053bc27431d9b3e1615fbf5ede27d633603a9bbdde1e6df0eb795ad9a00d07;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia69053f259b67f0fd728ca4fcd2bd39802adb86be01404890b17989eb74240db;
reg [MAX_SUM_WDTH_LONG-1:0]                  I108b6619ec88853b35b010ac5ab6a5c649973073d8523fbe5503a6ce91a78534;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id372f6f6b6b8b583699e8af0deba407a85b166caf3110f896594d222f0114cb8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I719ca66a3b30047457c24a43119751ee15bd686df9a03f81885e3d8b2cbd07f8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9b0a59eec0b8ceb485b7dafbff07051b5bd44c8b9ee4c3fda3773cef4450e78;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a9a7a98aafa77a8d0eac55b80e3c9a4dbc6b79d4a714c249193062b14ab5695;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic0563f05659ac941778904304c02575d9c9f2125ee05515ffd05749e20880d90;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifaa8161798b18d4d55533a337ff4bbfcba6a94e4f92c99d728f1b9e0a9afd72e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81590f464fadabf1667af046de2f41172c36389854de1ad410e32cbe3b719ced;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic2f50a4dad9dc0ec10f13868d7a117a26e43b501da77693b309eee3c9c713b1f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2f85bbcac9533694e4da81d1e86313ed14510ac8a37929a6158c888ba9cdb0c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I92edc25de8e424524b27a64e0970c549d2ee4d232fea857eeb0b9a391fd8a03c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6128d022628a70641f03bc8d1508dc00be5665cbb426ab6b2befa774ad124efc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09572043800626670079ecc4ff74ee7ff644d70879ed7598d124a0d5e847b288;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9eb8c67587f031f7dd6668286278ec62c632eebd218d4b5fca188e6447de8cff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b3e88dd84be91d43898b83141459d2ecaa7f53424793691b357a4153fbe885c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I930d8c08531d026f47ecb265d741cbd6a41286e3898d547ec9770fe114da36a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5947b18a468bba37f977f0c09103b82cda7962015feff03f0f7259f29d77d3b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7401c9a97f13630805f89ca9767771302df865505689963bf68db913a151a1bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e2ad7d4039c25bbd7c09ac2d55efdb8a8660f4949c64c3ddc3729f253ffd9f3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0533ded3a5c68b582fb4785c33ad5742da4947c904b1a52e05c80a3645f3fef1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf297726d3ad1a4e50327cce6585b2b5449e95ba1c222311ce9d2fa03c74dd88;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2616f37126555e344d3b2f904a46af3f8a5fcfd59fcbf0677377f16cd59f3be5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2118c0ebdd9baa8fcfd921632fb1fc58d995fc55e506507087ed673f52693ec0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia049b06c7b1e457c3ee5643e87fc729a409f2fa943275ce5dda083fb1253c2eb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica997f542c175790baa0650ff204f09e387d1e1119096ae7f1bf9b6a683c6b80;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6d785370057273f67048d3cda9ebfb0c8bc43fc5f34af47935e45302ed66e021;
reg [MAX_SUM_WDTH_LONG-1:0]                  I49b78fc64683b38b3318a903923a2523aa1fd7e2f3e13bfb26709a93fd8ed772;
reg [MAX_SUM_WDTH_LONG-1:0]                  If668ac9edc8047d257ed4f162d07f8f326c0c3ffed244595bc249275f04f02b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2965e4d3241186a43f93eeb83b4ec8d7e25faf3502c42556448bcca049d1add7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ecda1185b64bb196b1281095a7e3bf01377e6fbc7ec9cb20a3700f458944fa9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I883f00e2f9f6d78ae17d150f6305fed3e16ab0da7c8b4ccea0b9aae62672cce8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4b6ef863f3c19600f1325225dfeba21b5e9333dff55ddcf9f0cd8e8ec3581a32;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4611a21e5c71e60d5cbf9d62950215aee3679907ef0c908ba375182103b06375;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2cfed4bfd244233c8d85a9ebd9edd2c03f3bbbeddb7c7a32de444794e9c44e17;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58f661e6c3018394127a3cf6fb03e6993ca641adb970d8a7c0c2fe2547a36c94;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7e91102c5105c0ecfc871fce4bfb86900fbfc837d6f06f3229d362d20e51ae0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a660d35184450970491123819f2a1ac18ae2eb7132339cd57e564cff1dceac4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7643b1d4690f708c2c0d93adf0c5ac9ef99fe85eedc024e505edc74208d0f94f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93aaae3307747b620bdc3ad1ef6bd872c1b4fa81e99664494ff00b4357f1675f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I78f713264010c545a0147149b2fa2efaa92985405649e4c4313a0832e8222787;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1efa5f2029f0dba2f9a46aeafb6ad51afc192458717939428f80359d159e00f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6fc297df8d4527160ce05230a017f3710f7c026c6b11d64babe81959156f3462;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib4e74743b49becf72add5b8e28261cfde3acda86de12ad6d7ee855668c1c79f8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3e13531d22eb604e4a351dce5ee5512894170b3dd6f87962756c534438688ea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8aed9a4d4cda2feddfa8b481712f5723cd792e834384343bede45a150ec1b12e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I10312c661b621655f99ef4c729f81bfd1c6aabf28b2f3372264d69d6d177d475;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5f5d06e01de5ae4ba52dc9f61ddb507f1e34bdd36dceca20c19df859460eda6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic4b994b93547d46c87ce7cd1fff323144f9de0ff6e79ef0ce9ecc1db89340e6b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia1f7010c7618800ab0201f331741ab58055c31cd72fdd0e3db900aa455703ad0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I38340f75bcbf775a9e070a528d926355b818091cd8e5c1792450d2713ae436bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idba5ae25e3ea830381b3dadc351ea69d0e7b2bae1370ecc24dec6d408e7f0e3a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iad0e03f141449cf08d3cfdfcd976e4b5a8401179533f5aa4f8216198b749a4e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc06285b311fcba47b9670c971839fa401cb4c74f3da347961786337621bc629;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc82061cbb8fc5b88d39b5b714381ff331de2b2877376cb96a32d6742f3cac6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4332a72ae402f4043459e290fc47700a896e6eef5e383e720847ff34ef1cb150;
reg [MAX_SUM_WDTH_LONG-1:0]                  I49af7bf73e330c26c437d8f0447a930c63d4677498d07a28ff9b2b25860258d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I937131c2de1f55c3990b577d63b44282462abde126ef6a5fbe5ea962d48479e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e977efb6007fb448a0cd05362289e5bbace24ff868e4fb623ba54135e53fc82;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83e04a31ba3a09afcd0f223722c2852e314c79d93374a673cfd952bbe94fa816;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98233f63b47681b1d8b5e3decd1ab8ad783734a17e2b27c88234f00b23fa30cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7258f6d3dbef6e7ae01af1761728fc7b034158f1e7f26b13b21b500e1bf3e189;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58660674a5ad4c7022a05e5cfcd03fdc7161e65e8050cc59ae6fefc404b6b310;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3d284053eea1d128eb2703e23589b78e03e04e2b5219696ee3b70b3645c0267c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9612c348b28222bc7559977c8bd902d73267c977bfbe179506c88be746830331;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia14eb5936f779af58b044db01b8d6d6f89557eaa5deb1b16ddc8f7400351b6de;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifea5f415406637bbe581d11e57aaab23cecc2dc1957f45152f03d3006334d24c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7a3f69cd5191d002a2b8428d09a32b0572981dfa535a5fe1d4406ff3c5193797;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie56c2e96de8be01add59d3005f52661524c2193f6bd0fae2a759d4afe9607388;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a2e691f96157814ff15983f1dc0c522dfeccac15ebe1fa25bcacaa461170b15;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1744ca88c13acb5d2afa42ffe0ee5823eab5e32cbcf3248db4faffd6fe9e2537;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifef7ad6de75a930ef9a0fd7a22e35afa498ad3ae74dbf41596b9bd952bb82be2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2646e32dd3a69da746d970611fa0a89f96286df22ebdcef1ab746d70c4db4331;
reg [MAX_SUM_WDTH_LONG-1:0]                  I680a7b47f68662a83f4298c9110d5e5a04eb459ef379b69a53e7f90d371084a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4c7da80c76f8d8ad9ed1199810aaa919460f955b2745ae54cdea9276ad5e2491;
reg [MAX_SUM_WDTH_LONG-1:0]                  I343f02bd7da57ace84d1a265307da810c9ef6a56ada6ca3f1e102c8e4d53d89f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e411a908fa94c50629647023bf56aaf275299c8c49933fe67ccf00d3ed68d7b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83858f36d2e66e2bb6f4357e978909888d598c4ae084d87a74d06f3ab7c334c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia06978f4049096a298ffcdf526e89060e8f27418076fa351962ec6f407576753;
reg [MAX_SUM_WDTH_LONG-1:0]                  If9bcfc0a82ffb81925d5e0fb3b8bd0ebd910b079c271c352751e38dbe327f634;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93695abbc93c5e195bbc5a1fee05aa7ceb4c58b273ed67ec6f28538aef0843e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie08a9d45e117e5fad39310981ed379f876f4330ccc7674752b26bfd2547adcac;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81b17367c5766001911129ae2370c1dc7b3509565fe78fa6e552b7ef936da360;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice7416e3625bcb882a0caa84958b2d20b2a6901ef7a7c748ada330c86ea41763;
reg [MAX_SUM_WDTH_LONG-1:0]                  I189d5a40f26a8b2893b53242a4ec7613797831a4a2192289df09283c7da753d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba6cd77ac5adf667b7d229aeec4f15eb6112ab90e4b51c09bcd7c64912cbdeb7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I15429bf02bcaf6ac17ed02efb1e65c5c37254aedb9ef6181c2731c3f7e2a829d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib6cd4feec46af9df7727d5febf22dfe6059c43712e65fc7d982d1a6bcfeeba61;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1807ee521c06cb799faa136864a31c00869398289b0e3b185e702f42cb0e7412;
reg [MAX_SUM_WDTH_LONG-1:0]                  I65b7c3c6e73e0f305942123f4ce97d6765b7bf86e61a3388774c36aabda5a491;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id4ff3dcea8b6c38c5288cac263296941b841255967f2f58fa97a49fadb2fd2c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3525fe2422d10480b4caa9b5a6fda0228ffa3bcef28a2592f1eda3194cf30bc5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3856054a7ed02c524f8816bd8ba22a48935b393ced40e98c693416364ff512b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id78e42777220c16c860f907907256a6b28e2c5bb9cd011c71943ada87d30a9a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I358ca9d90eebc0e19c434a7d1070a69b3c20b4f8152adcc45c0b73e8cf2c9902;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c427f570b0c040928fa6aa62250920306e19e3031494e8933e30766f0c782a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e60aaae452f97c016f3f3929c33637509d02988bea72048f7901a440232a85a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id55c37de3455c6ed8da5c25f25a98b0ced5787638a4ac262c1bca6fafab7240d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I312753748b2d173f2dde21bfad8dcf880f5fae94cd73fea4dbedb01c43c99b43;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7049605331e013c95aa5eae16577637a3e8c80f5e4c325675654dcbbed1b613;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6f210ff43165afc5b4c3a9a22dab74940c409a5fbdf9c47b9eaa68fa08918f23;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb9c4b9e280f7dd8b4c34242a9e58352a23799e10c7abf9c3448e8a28af55e33;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3422d7c29697052f1d70152dce7d92858081099a7bd19bcb2a48add3d660ef12;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3f33ea5e4ff428c3f59701f77e6f288293231923203fdc140d147d7ec769295;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90ed9972249e176fb13ac19818b591acc7f7048588409d394fbbb79ac26b3519;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieee64ec5ee871ab61afdf8c73149bb2fa68fcdc0050d80179dd9645b4f14a201;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee565a93d37ce096492969d59077dd347ffeabe00c447298bd22adb6f66926dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8cab52d76008f7803024c4d66307e41aa48256ae1e9d364c354b4b3e405e5c8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ef1e4ffe1fdc795a0b74f93f87b834e26e14a3a6cf78496df39c9cbdc70a819;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7acd9d954e3db160301869bcb6aedd5652613816ae8340f271aa4f90b9ca4658;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7bcdd7375cc16a2a91d81c5608f9953d21293d5121600dc475a15b190967b143;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e3bcd83962abb7b063abe3da76e0bc387b63894a47a4f50f9ae7abce8b944f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I75bab5d1e71ba5ad182fb01cfa39d37572ab33f5f848dd0775e3358154e4644f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I60f85c5d32cf353d7191d12cc29773a42aea456697214a1249353a6c2d7463c9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f17ac4c0a37a850db6a1d3c1a5b2483c0f3afd684853df30d66933c8c593d03;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia9665e417120a907ca7c884c26250701f6c61f0e97c21fc62160f80c74ff05db;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6f8e6ce3128ce55b822fddcc664d0340c940bc85adbb5c93acff37548e3018fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5de5cb17db6bcb69528e636b4248c6995caf3e9f30dd363ac514f8f68d651ebb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3234faedbd9c50f29c09060c3f7ad76e44648841500b09c499875ea77aad9537;
reg [MAX_SUM_WDTH_LONG-1:0]                  I20647c051506a783956d48236b4a5097f9484e404c42e9176d52d59c8efe6c5f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74189716f0b6628c0d75d54cd0815cd8fa65b9047c3f51c5218fa0ba7b7fc47f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I898c9cd15d2ccc181e81531a379b969a0bcc87d38b0f3a9f9c413606bab42b15;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icaffca7436caceaf13fa42e9e496c7b149d5931e08057ec92a73fbeb9e610648;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie75a482f66bf63ff96fb92dfaff210e0e43f91de86567ac2bd323fb0017a9f62;
reg [MAX_SUM_WDTH_LONG-1:0]                  I13009f7de199aa969d82e233d26476e44aa1bfbb7d8a4fbfa0fe4f1f1e7579ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I67d64752ba4f83a2592c0a83a7ff2773e71e84453dc882c23f8aec987abb6731;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8c7ca4914849b513537d3688dc1b76461348ca06e80e489afb60a2a082e905bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37387450a3e4f68a3f1fb2cd428d54ffa4098528dce70e0a1fe3870830602efd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9117209a7cbd232356943389578d67bb7d6c217e7e40bdbb904fb46fb00e9385;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7db05f66d2fad420c57a7205c5a1b9d9036f088c64b58031e6fa82617923544e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f16d6ab2d87cb715b071b05ad14fc6be271b1d7966b71c80795894643e6fc91;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62c3f28235cae0fcbc04a55e0e578258ec501e25bcdef661063661346cba651b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9fe8ab2f590451df0986a4f7a74194c27699bdfae0f182440f4c1875633cfcf3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib230966e790f9859c0c85bef2949dd2fb9fdaab81865b0b294036d12648fede0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57876d51522e735eff337a69dc597cdcbb100bb3d3e0e541aad4428637f34e26;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94c80b77b7ee413cd168e55905cfc4beb26ae2f6cbbb944ef335f47cf424086a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9fc6ec0055cf4788a1f382e41d1bd50b2ee07f2cdacf368e2075fdeef55f53b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ffff1f75581c6409c82505e1ad4216ff385151e7d592f1d59a1d983eedcbf82;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib2ce92509ff0447a434264639ad96df47b161136cea1535b3e802c0c4ebc32e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I979f67eb071e28ab1fea67ea8e52910bd67827cf1dd23c07768c0c237703e23d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I20b66d31e195a0db14cc87da1f6d8810b5f1056c2250bd5cfcb02fb4edc9dd0e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I39e3942d2695061c6bffca3b7cbbbcd0c973e8412976c07d2387e9b05d75246e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7595f637907686de85c9038415609949a80fee8bbb0c4e9f3873225ae6c56bc;
reg [MAX_SUM_WDTH_LONG-1:0]                  If17d9a9ece84d9cfc9fcc430d453155458b6c8a7a3ecaad974c8f29d71b7d440;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6d41031fb10896690dda6067df08ad914896baaa5f83c46b4051cd5a02f3baef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia3496c8ef63a7e37f4836fd3f0bec02370cc7614a22a1756e61fa1a536f942fc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc6c8bd2a37e01dec18007c8fa763941f7016bf299e3cebbbbee3066d4bf8c7b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79473cb7e5feaef4d80685528a576e134e739af85c92bfc85278f949ae938a96;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac1565ee006c23dca041f0aaff4dd7023b8a22cb72c9f206170be661a66d4732;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib6f1e860bf50cfc54de5c515cb40c392f0fd1f02c325d52c5e28cb5d3a811a48;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7318d295676d4cc0682f246020963a6411be5cfc2fa525dd7af0f2e651b4f9f8;
reg [MAX_SUM_WDTH_LONG-1:0]                  If9f2c8dcaceff8232ed4bdc9261d1ee5adc0291873452c335748d5bcca9435a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I596ee6206f54965079551ffb23aa3c1948f6fbcd48659c4e30b205dd06de79f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic215b986ae9a8ff5c760e17d5e71da08756ba48d0f8874e35766d0f8fc18b061;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7c8c24bd3806dbea5552d386a7363828eb5a822bb292fa0c14ba407a1937d11d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic945b809e46ac7f930479330040e1b167e8f5b96a0583a39713a34261e764ffe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib7690a963a38d899184e89d3e51ac5cd99cc0ea9b2fca1c2e36e51ea65b893ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  If6a91bef840a62f8234c19c7783b8ec5d1910ffcc05eae66cf63c1bd541c5caf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie55d9e9e5c4a66363393994597d9138fccd6c11a2a6c939768b63d9cf933ae1a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd9c2cc79d2377baf6c47290fb8b0671bebedb2aa72b90f8d9fe98d0acfad39e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2a5a1513f2b8c1f000f58640c3650ae03d4d56205a8cbd04742be5b91c8c594;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic655dcfe5a7d40fcf2eb0e61961010434f0098e4cb08794fa7963797c764bac2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a2e9ef69e2c24fdb342d3334d2b71a1bebf10ffe1518dc5f3ebd5ff34dc719a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I302186a080a24d93f21320fc1165055fc1a2cdfb86171f35cc5fa8ee98f0e1b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8052be48c5148738c00fa7e5be66ac6898d51e7fca2e5905ef028d897d47b236;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia3900ae4b178203e8a6aab20f112207ecbe30e66c7fbdff63d82e1bc1c9ef760;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc4766e0c1913ae910a794a3de1155638a9352251d646b270e3aba4eac09aa31;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4734d2e489a9d1d0d797602f00bbd0e63d76f1ab0bbc514401ab815d5ebeabaa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2322db4da4e5112d362e202ee964c08830d852a01c92f802c1c8bc2978ba25e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d325e738820d37fcdc02fddf7899f4e910dc410218c77432a6e47f1f9a956f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  If29e3e5b3c3425bf0fd40a98d32046f215032a8ae181688dff1c4a253b0460ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I66cfe3b553e345d01602cf9440774c8383b14922fb66580046e0819ce297b0f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I51e9d69995015664cbb95900d25d26d386de1f49fa7b7d612964802060fd7a8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I00c3f248f180ba740d0d97e10760d76e4d9033a2e4125b04ff783a554db09b1e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2af69278f44ee2d81c64b9447b85bd09d2ce2a8dc86bacb9a175b33f72d4f851;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9954c6247025cfb8b0264906e6dc6a703b9dc8d3c4f2736930fe68d278dad962;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib82fbfc182e6598a7a8dbae45ea083d2922e3f10e781ac40e1c89f79097f1f23;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc519e00af8bd07f427774d04fc48f95781295dfe970673d84feca42e324b583;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3180a2d7f37d66f9895c1de89329e69ef7e88d0808fce147b25636e639efdd5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida260241e2192ba6e2a1d15acbfabfce6023278ca1f2be17943bf48d0b95d045;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb545544cfc26097f08bb8236d489536608fd3ef900015de2da0a8a5dfcd44ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief91e723aebbfa64c457be6ccd3ed8e2faa4703c627ae36bf868d8d970bc315a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90ba4bf676fa4d1eb6132a37c0b4a580ef39ac1cc44d6111b84d6c7b907922b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53a559b412f643abf84ed01e98377ed96246560bb003bd28eedf2164de2c2db4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie66d53b4bed43cf8037cd1937f7562e7bdd6cac54cfc8313572b853088528a0f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie685d62aec7093c42c2c432f32fb1bca42a9af0ceff50f2ff2ffe57f0d98af75;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id812808edf2372138b1569ea1a2ae0583ef70eaad98a941b8394d5d9efeb44c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaa2f1dc17d04b53a43d7435ff62012f950453b06af95243f1e1fae92885e9480;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6b9daca681053a70322aec979459e65099a78668854de86dd3f51ad58c5dced5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie74bccfd27d7ef80fd7b51b8e57ade889188901b44e7236766861e8e9601fed5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieafce3772abd32b8004981fe3f3d102d629075a15b6dfff65169984219911dd9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d27f6db1cba68a36e75da65709b30702412affd297564d2b4e563e41db875f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I279bb276ee61f29e0c143251191c161862c9d95cf0bf3a3fdcb6b3d6acaee983;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0fd6ce3dc520f3fb4fc9a66c0abe0c05b943610bb0bd11b7f9dd10befd5c0b99;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife98dd3babdd2b2db4edbc673874d3f8f184f531c9d96b1a89b68ba60a9a57d1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7a11ca0ad51e87c9eae3a026eaaf462f9f4757831277dccbd25881de07202e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I038f11e434287c1e184cece6178f4ce26889bc2ea583aba8889b8953306e2e60;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9abd971b53c2f6c0d24fd41004554d3175db4b8fd63b38c7667ff78272cb26ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I25c61073e64c8149ae96f3157045d317349321841e21a3d69b3baf3bd70bbd03;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24d9c2b238ea5964b3c4bb358f301815fa15836cade3b5ab5ceb0e81a6d3a6bb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id156956a3b93d6a741a81c5a94e057e054ad7d4467a54a691bbd147afb30ead7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia755a5da1132f62cc35903f93050e9743df11befaba728cfa055601606c0caa5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4eea240addf4997dde0e268e6404bea936a04629cd4d244a101a6a38e6ec03e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4646084cb89b559ecb864051cae61dc568e6b9c6db4f1030904a572f7e58a22a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I536f7bfebdfdbdfef2f9b530022a63e1a70a1ef0b344d7f34ef956bed72fc94b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58754d218860b8400d1e6ffc21c817a447bb64d182e74f0d162abd70e15c5db6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53a83ec9af418aeb6869bf9db2b0ce128564fcf62d2a16506906303025076ca3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3a8f1a1dfbdbc1705527f0e6f864ae594bdb100ee8b14a349147d98da860f09;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4644d5f1dfb72ca4669b26a415cb9aeb54051fe8d28a6461d696f00bdf6c930a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If36c8f00155dc15627d5005ff98abb7a6eebcfa62de82fdfa50d86fc6e7cc166;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie02a7d9471f0915572b8db6797d0ea1f2fa380d96a4e02a5783e584800e6676b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id97692b9a9b0e7edbdf517b47ed0b87d007cca8fafa703956ffc2686b727ca9f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f39af323e102d03f5089838b2b6576c03169135defb533f54e57d8450f1130e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3391de01ebddc6f92c31c74e3b3ce12ae2081b56b461ce9e890a0fef3d14fadc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaaee3c7078bf1bcda85bade0d66984c675177a0f1c66c58f47e3775916797a57;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5f3145a0720b745a384e157d352823fe10bb6436875a5c52ad6c81c882d9e9e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifcc101725d905f243fff4a458ab8da67311d5563911d69daad960072e1927054;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f807b6151726e387854a9a6c778b3b069ed5ab61b41aef6541f3c2330b71673;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5e789a890f931a53acd095741f7a5936f15da9e0007b159a3a3762ec13223f8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6bb8ab1ec9d2824241e526c7aad88002dd83769fe53a79caed88f4f25929dc8e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7fa79c98c1eda80a19d8475857fb44ab41c53596b0b59806fa776d4c4ad02f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5637f02c1a3f8b9ac950dd6a246e2721f9e4d30906ec3662975bb3528e3d7170;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c1edf3d3971f7ab6f93e50a9500cd37fa3bb42d75c70d236f514e4c15a61f2b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f381294ee877c6e693fc57e804a48a9efe7e3289f2967a006a7da1659cfaa3b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3234b24482f57a12d4db307382a5591bd66ceb0dd4bb120eadc7ab2770d003d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib31ed62a3528251d6f00b4c346c776a8d5c3906b66e951288449677cc9865773;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icaa9abc6adde275d5c5011fc8cf6ead11032cc1bfc286b3a392ec507e4ff0d4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  If6073191b5a616ca29300286d02c0ea3f8eb57da345d41625650caac734bae9b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc444a5134bbeeda6005a847d5ce4e180e6c809776e32d1ac709c3827d1d84b4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ac115af593010e9556a2ce7fe8e479b1d1d15b34750a8084c442b1be7a181df;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41fff62fe024b1bc1071aae30dd931c1dabf2e12d0d1cdc295bbbbd946d63358;
reg [MAX_SUM_WDTH_LONG-1:0]                  I306ef55d92e069bbb7dcaaa61fd648d31d246928bed83dd8b2764f94de45356d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ef6ca3a27d76c9635bc942fcfb21cae619dc5b7bc842952e2a29f7f2915e62b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I915bb804d2926482383b55712d495d9d5a5df9ef4621a5ff8a2a4d5bfc882c09;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ec8e7e460c616e3d6459dd35f82ebcebdc1bd7f9680c38489e292be831ada10;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6cdb31ece4d35306b0d4aea87dff3b178f6664744c85f6307e1c1d6153d74c72;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c396eafe78ef3a7c94cae71c86a808a9fc88960e7519256fb1c0b54bc865334;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4282e3203fc14bbe70311010f6132cef075c94dc8fe22dd1f115e58e560c2652;
reg [MAX_SUM_WDTH_LONG-1:0]                  I78382168abd43ba48f24ad5e574782b47afeeffe0632ae5b4aeff07ebedabf4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98cf027b8e2ef347c03bcff057b551436e1b053e2439164297c60094d957f760;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55de212bade4801bfd54acbc885f19f7f43fc63874f6a531f8289cccb06c81a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8a156bf85802162d32801b45b639076f8ba98827cf96d3e1cb48a5a3b774b491;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia4c73e87649527da20616919420137fa4c1c8cfb4c85f4728a8441109168c6ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia9058e9aec6d06a5fa6d715e681719f75ca9938f6fecbce752a4d166fb9f2bca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I04eb84d9339dab27e5615403aad9f09e40f6b123c73c8c8fd6c27f8e91ed4af6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2db4e765057361b39c8d20e87f89051b0016f067baa15cf01865623088a9b984;
reg [MAX_SUM_WDTH_LONG-1:0]                  I49fac311626d99832accfdbaf5db0e3da11e0d89693c843295ada1310a5d8f84;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4203cf0a99cde14acce3ce3c04a6405aef0edfda7026924b1491de1d42089051;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic15cf2e839052d47aa87202bae190c69e5410914d9e00120099307d6f7a663c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie8a61b138cd654efb72fb596046bc9d2b50c97e34d4a27a1d457261b4f8a9fc6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74677cda9719646b1c842acbed5d3b13462ef153d0a8907019b2553c808f84c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied33aea50e5d0112a854d4877d3bbcb4bc21b4ef75e4b120c0104770d83aeec1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e0c405b4f7107ae7d9a35eff8fc48672c1ff35ede5dcbaa4340926c9d9e65d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac16fa27063df4a80f23e3757dd21e3116aa16f591d7e80e7079571e2f2ab6b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1db1a5d4e476af4fb7bbf80331760238438096833616b30904a4b6fbe0057e63;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd7c491a614817929db2d44117b8bdd384f7d9387d4bca021959efbc58fb7b3d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I083b6e833d8b3bda9d56f159a5e297305e44fad9f2024a3204c6e5b7afca9405;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9114e7211d58cd46c3e15d782c0822ef34b1436c74a1842a8af9abddb2117c7c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I410bc8d9b13d79713c47cab785cae1ee4db55ba3e7a207519bdbc646dfa815dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8fb26cd47b8f0da1d89b9818685edf5f9c9776e0df5beab4ebddd0e3c616c7e2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iab1ad3fda6ef48c15a116045600ab96f057c4e2769b1736742ece54e049a9884;
reg [MAX_SUM_WDTH_LONG-1:0]                  I207e7042b2c0cdcf57378c651ebe265368b8b922f54a33e5b327d55548833526;
reg [MAX_SUM_WDTH_LONG-1:0]                  If01282d291c85bcab01b47104be9ed13915609c85c61d979b60b02847a685e4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3a032b15228b0da60d25deecdfa1ec1898c483d70e6d08be8f89248292b2fb1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2c3551c0a960cbdcab2b802148c759ca7c8dc401d98b251d9ea21d6de16d3bf8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida75a6cb83f408b8efb2b6a75c221c6d3ec50c673bad1265d400a39da9eadfee;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7977549066f72a2e4c0d91c592a5d93a2a64fd1ac48cafd6f0f4600912f3fc1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d246b2101b98789f6c8b328fb0184f6d02065d04c6935ef49dd5baf259c1e54;
reg [MAX_SUM_WDTH_LONG-1:0]                  I08c54adda4326fbc5985605f17f5b1c47ce821476ba25053aaa7449a571bf33c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf193fba82d63a518161b53b8a23b3fbd93fbdda529aa080fe932edbea6fc57c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74a65dbb33c6088646be4339ced1e6167ed3c67fe3f520e10d4fb2c96358ce62;
reg [MAX_SUM_WDTH_LONG-1:0]                  I351f23377572c7cc4bcab051aeda29360f51b89eb290bac8e484fe05adc29065;
reg [MAX_SUM_WDTH_LONG-1:0]                  I378dc69acacc690da268354f08a9f1fd08b11a899cd2253c2cca3c979245a06b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id85a42323f6615cb44efeb003b9a3bf7309bc463bfe55bbab0aac732f99c975c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8519733c2d4de3643ecf515bc788e665d7661c947a6532dcefce59b255fc05c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I77385a4a50aa8eead5b897d5c076357ef507c90dbfec7d442ff728bc20b90048;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b3f1cb9e25ac68c67abdee581e7dbb74b039b9f1f04459e3a4049769f27c474;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ac9c9564bd70c4a8c9a6a76450dae9f55e8008338bb7d9f85f52e06b17ba7fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id79e7da27c2a195d433419bcc0481ffe12155390f0a10ac6be75723cf2ad53f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I02325f467c1fa16e231a42dbb8e973427b2a4c081fdb336e3f3838d5f7a7061b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9aa3880979a20743da2aa753686d0ecaf0702008920d80af34d834ef1e2249be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I389ed2df5d3890d3c2f628edb1a043d51a972de9cb338f32389788f5acd90028;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie591b9c2c777632b671f8aa86f6befb3d02e16c23329cbc7c07438588aea4c9b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9e38d40473faaf687741f97150071792a45a4926ec46762a3d1729e7b1d7111;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibaccfedeb751c2506a2342df2f75fe492accc5c68614fcb90b4f5c332c088808;
reg [MAX_SUM_WDTH_LONG-1:0]                  I49092cce392bbf2662076c5d86322bf8c9c77a778ef3893fb58e9b08396f2d24;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa134df77ff670a0cb559c384c786af4de916cea66ca13147d43f4030d474d0f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5b1f9cbdb5bf4a096a6c8bcb4db57912d6cad99055ec47831516d612f7129dd2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib378be3532348ccba868d918209ee3f013c1844044c8a93467a93c3463f7a36c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81a866e481435399f8705efd8f264d7419c1acdc086298638158f4d75202b567;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib85e84ee2add613edb76e2321f7a5d6b4de3be9b1ab97905b5980277ed273dd1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44c742e7ad2e3e18153ce9b645fc21efb4e3016f063b05a8bc1825b05a303374;
reg [MAX_SUM_WDTH_LONG-1:0]                  I10ee9fd16ea681268e4bcdcc30b515d990dc30d3fd41e059e9f1dcc80042ae1f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff70805870814e2f1b8de2513c56a30b9e6194298cb863c87a6e75221c8ef1db;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic33e33bdd936748553ff29221e983dc115121fc84bd1a2799a3da8120be82c04;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6188d9b90b4bb155ad464258b5d3ae28e757f4b3ca73453ac4ab3d6cfa8e6643;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0705a3be469f22a69c0c4d2366fd0eaee02065685349db5abd81049530fbf842;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2603a3570f686ace17fc46e9c5190f79e2cb32b4e6d3c39c26265951b22dc00;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic0edcffe7bf2caf311b42675297cde79af81c022f660757cdbed53dbf5c04eaf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97a0471ea526aac1fb508c6cf38c387c6afd71b9089e63470279445f4ac8f7a0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I600367d873f901e6b7f92a4f9c0ac92c9f8efa6da1d6e6945f83b863e8bb8519;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia2ebfd7cea041d6ce3b26d85588f2113701cf7f6970206eb4ea2001c3ab0f52c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e30a7f3eb36b84c9df9d59f6164c757c8612fb12567ddfd03c32388af750bb6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41854c843f5042d94267a6b9d374dd0f5c46fcb45df0f40b587aca943f7bb396;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8d123ed314ee10c10f04151727cd5ce1e836c01f0f8143285b54425633591008;
reg [MAX_SUM_WDTH_LONG-1:0]                  I542e912b5cd0969a23f6d60abd1923cf0d333b3f20df92061570f156f395d756;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0ae31ee6a1c597ec90ca13dd69a651079d801c279292523953428af55188ddea;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib49bc31787442badfaedc737b3e1e4014bbd7818595fcf9cf42f23dafe03fa9c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7bbfdff59068ad7e527ada31d96fd47cb737e6b7ba56b1b2b9e522fe3a63a954;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3069d559ed47e3e17dfd391829deba4bec9932d5ceaee52ba24e585c3ca750c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I09001eb04237069c413098f07bb41538c6d39b0ac000f175d61ee3c0b47cfae2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74beac54df2553b0529872dab3dc06224f214ce3e1028033e9830a31dbc6b036;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iddcd6e6693d5f625ba82ec2cdb0a93ca1826dca4989d19221c8127513648eab2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2213f69a2b20b811c1ffe8ddc5b7a0c31df06430e2d02679663fe31305bb6c87;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89df294963327dee66a931b858b05dddd97e3fe4d048ecbfaa9c15e28c57602e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85dd7ff4d35dc1bfbca02c07a3f89560d8b9f8f10c9f28ed1709e4e00583b5d7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1f0110f45df674628a1a02cf01dc58577628dd88049b93ebf02b5c4143781ade;
reg [MAX_SUM_WDTH_LONG-1:0]                  I385ea910caf7d0563d1214dbd983b37fd5cceeae24015a0b4cc253612b316c22;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0995588ac28564326a4dec88344ddd733075750fab9f4f8fec64cc91b3b48e2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c1a4f9167a1ddf22a7642545eb95954fe17112c630b62d9e95f899783de734b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a2ddd5962242d66fa4b8bca39a81765dfbc6c0b6b012ee42329dcdfc12ae9b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I231bdd513a7d05321aa7ee4d1bfc4b59edcc82ae92b1e27403f0773bdea92e92;
reg [MAX_SUM_WDTH_LONG-1:0]                  I83cd839beef638f212312a0093595ec3d71dc80e240aba892f6404de6d614bec;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0b5d2604bb5b289b82f24f9e91c4669cbbc04d0e3d79aa18ebe3dd27374837d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3420837ce14103293c9ee75848088cd144ed5b975add2adfd479ad10eff552ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44a2a1b5e4fefb27d702cad5d65609674fef85f845b8cc0da1c6122c867d9317;
reg [MAX_SUM_WDTH_LONG-1:0]                  I641204b71e0368d174adf904e08c12465fc7a18e1adf1372e1649efad206ba0a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic3e639bd8b640b9a08515fb88cb35f8d263c8b4bba6612a800b303bb21974a4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I10bd3ad7827da7bbb0e1170d7e495b88ab6ac55e0421b4f208f5c1ccd722198d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85f4e180cb842542efe4294bad76481afdab9af7982dbc049af943d3fb23787b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee26e4077668d0e7329068693c4279480b26e4f16adb0161c8e7f87de802a14a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2d2a89c4664389a9d5615140b32a9a994b150385e23a1ba81bf0823ae34ff5b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8e573753ddee4fe18b1f9fbafcd135efc7fb7e7eec52e45b5148b0dcf346050;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idff2c2e52bd3a5b88eb4da782cd2bfcf9621c26033b6643a8ab96749a80c9fe6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie8e89070910f06608a4df5951936faf465b4f235d92b3cf8a3820d03bcaa83ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I13ca4018c147e25a38463d2fa98d04240b46a846f1b8b13f69b99942a4b2539c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1a0b36a215887b4419ebcfbddb0ab8b4b9b21c4643051db135c9d9ee53c6bb3e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45e1276a5f5af744327fb6f85b50f8aa50bb442469cbda4ba869adf5a8d0fcbf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84694b26e240bcc3e7c9b224ce3c2f5891fb546a4fc11e4597819fd9827c3105;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie63f997e6206a536a5e45901da6593c5c49645e6cef643846980c4e2070091b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie69f3ad2e3dcb172e525302a533963ab9a2a08af8d1ec71e07d0946d393c056f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I275a2a54f37e000edfcc6f35cbdf2ab6c2a28604ce2e6dc31d6430693c2ddd4a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e0e1c5361317aa91a6e54e23fe2585744a1ec47fcb2412ed152b660781c7832;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5848db5ea2fd0385e583946224dbe078419a4c9684d15157ec460537baa30d91;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia338a53ab734049efb28655e209908f1fd2c5d19f8056463d711cc1e50dde602;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic0dbeca58e8f490493dc5672f4aeea9b98fb9aa4aedb922714f3aa21a4836223;
reg [MAX_SUM_WDTH_LONG-1:0]                  If63dbf3e3c6000184af28e72b5f2960f6a376f509d5693a96d2ab9f92ae7b237;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7363f53cc60b20a744ae33ca65adb0345b104fbedfc2ddb5bb00b1dd50bc13d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib89d5800576f979f189d88e7976f8d49b8470bcbf6b365f7cc6031735e3adb4a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8ae67d7680689c7007d27eb5af9c5bc1277025b9ca78c804632ce105d41fb08;
reg [MAX_SUM_WDTH_LONG-1:0]                  I622321198c6f868e554b595d1e1616dd63ad46a80c33bbe896df9b6558418ccc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f21d46e9cf807c74d37e3d383186daf9288e68431e128ddf72f9f448f671ad5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iafcf26b8f2df7719a0b660b41de28c5a325e50d75382579e53aa9d065bd81cbf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9f2f5a180ba3e3b29c209d7e3c735224fab3c309f2dc627046d864a58f42897;
reg [MAX_SUM_WDTH_LONG-1:0]                  I859639da611c77242efe899343358a650652277ea45277d9792b619196c66a1a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6dfe9c7c9935ceb07f55d4fcf7feea54e13050347b5991fca21d79ad74608aa1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2899ec4e420edc766050ec0042965f87c79455271a54ba7c947e94d37450a033;
reg [MAX_SUM_WDTH_LONG-1:0]                  I65290aca857afa1ad9b6aa754dfaaa0671d173c7b3d9fab7cee9ebb973b32862;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibb256fb3d4bbe6ddc65378ced36e01255d8164d29755891e06fbd4caf2a290cf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8748f772ce4e677c9220c1fb10521d69acb830ffb623c0490c1410b515445dbc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I60f4bae66121b814e2faa564c162bccbd2ef0a73bcaf10c3c78e30ff2edcde4a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id6123d9000c37cf18ad9bee82fef91900b7ee165a1841b5a4d23af27bcd0fbbe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac70da997560fcd3949fde686e6f8a3dc834a2ab7ff2beaeedf7614710bbfaff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e43798e3391bdb6c6a9a6ad85e51c960fe4bba982ae765cecfb287b0573e5ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie32e4f67efcbea2f033a66104b3315b46a1c857781ac63283f4d955384bcdd4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8b3199a20ef98c9f204d2a8686fa71d5094b2e701c6f84b7630ddcce89c77c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4720d84525310ad5428da40677f1cd99365d1467c29d214ab4ae300277322cbe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I916b56be359d608276fb2fe1be1c65df20d635e00211fdba107a1d6f9c0f0a36;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia1f10017528e76925426be916c558186f2196a0c4d7520e57e0895e14e7c1d53;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0b3cca386cb4a6627354dc8fcb01c27aebb58435b78d7df234937d5aa2bc457;
reg [MAX_SUM_WDTH_LONG-1:0]                  I46a3710c0e472a92b83354b668ac21c775b2c4e3dceadc49dc0cb712c08c319e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I72ad7a4f024406e89bfc87296a9c0456459b729b9e4adb046d703069cc9ed1fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I594b73c43f22c1cc15daf1eb602be4366502100a0ad3a3bad7b7992c9839dbbb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I725f7893c803b548e668b87cdd368f2b26e58193cca109b618d87e949b8b0d25;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id6264ccfced253e14f1f9be10f967d475695838c367808b97abbd7578447179a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d49190282814ee6220a4a003e2f4879a2e37459fb2c3a1e1ffecc35f57c26ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied0e2037bbb2f2b7d0cef3d7d3f5b7123c006255cb7f2297df7e1a1eb03dee16;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iebcafdf2cd96dc5a859f7087ad96383f07d57818696f1522555720021c3fa8c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ica6a39f57caae5761078aaf00587554f1acef5d9b2e1fb73931f5715ebc762dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8b5082d5099ba65d612d86118ba3489888d375a6d8dc1816ca6c4338150b98d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0fe26cc77a5b117d82b8f0da27f4cc5e9465360eba32d35aeefc16ff600ad5f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia11ca5043541c5c51fba4205915afd0b4e97bc70d10317e9d3b952138dd15572;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8bfbee6346d016ff8cd0ef681e0efdf28d0f27b3e887397fa1aff647739e25a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iefe655d513457dbbd05f22922accc5bebfc22843447254ee0d6eb4b48056884b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57f07e2955da5218122f614720d5890af9d7b5ac4f033e9d1c10db08e7ad1882;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e23dd0658534242ac135a6b401ee146d0ba48841d3464a8c58def92970d50aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c71f3f968f3265215ce730a5f922db81aa408218fc76de3b64ee4f9396d3f78;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4190e8ea4ed62c9f3512e102be78d80de31e05fdb31f39bbecec25c5fe4838c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3afdbbfca5c952e1800c1e15ca629173eac62810b6bf8097421addeae979ca81;
reg [MAX_SUM_WDTH_LONG-1:0]                  I22800d7bf254d48f28f9d0e56af31271b20bd989575a3ae510dc64f592b1e08a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9d906bda89623d793bc65968cd86bd0c63458c7a6b12fd38f7054069dfcd132;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4bfc7db23a7b268d945c751ac989718287b1730e8ec35d623ea7636b6946d554;
reg [MAX_SUM_WDTH_LONG-1:0]                  I969b9fa05c651f6e2f2dc426e35c43864f9b5c6d4f6278b0f7ec4e7c5e872eec;
reg [MAX_SUM_WDTH_LONG-1:0]                  If4a3f6ad253dd104911b6d1a09ae4a3ece88afedd537e8f7fdfa8735aac88fc2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I436c98ccee6d1a138f1c47ef4e5b7ac39db15122b2b134828b257dd629e310a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ec9f763c06f61ba0e1a2669b6ee19aa5be8a80a6ce04c0355956dabdad55e9b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ide4ad5678bce6a696f0c6cb163eaf670c47c2506acf7977c1031c6ec03e03a58;
reg [MAX_SUM_WDTH_LONG-1:0]                  I280472596040e145f7bf9d23aac7c569dea951975e67e53b2677fca092dc4fa6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I043258a364cd91821e9bb3e9c46441ac7d330c706e4b0b7e29c4b92f7c5ce562;
reg [MAX_SUM_WDTH_LONG-1:0]                  I593137c88d2dc13a0bf028b949e6ec556b7787557f6a5c72f0d1161db6b096fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f639b76b1afd86d9ba4d07d54f5b45df8cb99d7bc58cafd0c1a9a9001842260;
reg [MAX_SUM_WDTH_LONG-1:0]                  I331fc2f98c551ea5b177eb3f3c1072371f7f7a02e45d4ae3fb41bdb96cf7426d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1dd0421d7e31a316541c339f8b4f1e3afbe37ce09254ed825c1b6086a0c0f3f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic5a2e5d00e362ead90ecd9182e61b0e3a99a7756994cd358bfdecf8ffd957491;
reg [MAX_SUM_WDTH_LONG-1:0]                  I50ccddac87e61ba10dd9410a224c74ca88b521dfed962bf601c38ae78299384f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I15f2b29740b5d1a9a5412db4a0bf09bacbde963b08c243ebfbb4740dac56349f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5fd9960aaa562ff70e5d0e913dd4d88aac1b73a95c41ba903c0b7fc4dd4d93b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iab45b41ab7c1056072ef64483afe800af63354919bd1a7ec95cd3d9219ab0301;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icdff2336860758127c20c1d45d5723511fa42577417bf4f77d0c770abcbb175b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I96c8864be45f3a0501bcfbccd5bc984738c1e05cf6834d8aad47468465908abf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9351e784be3825e94dcf67151cf38c9fddcf244bf5512db57dcc612882b449ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic01034eb6c2ef07602777d1a6ce7195524d4d1e3093d15966e36f45fd58d5bb6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23f7465a60acd0fb198e753834d30932ddab8939bb2df2172f54c7bdbe02e154;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaabcf58807b565d00812cdda849cdc45a34b1e0019a539ddfcc9aa957814de19;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40687a0e9fee803f38df7cf7dbc3d3107b859b4e80822bc59a157fdc606416b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5cac542afddc74aa26163f65fddc7689b04bc5f3bf1fda74a7557cb4dea506d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I807d8cd303e5c8c8379a9a2954804c606d897fc06412c924a89f3dc9e29909bd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3fd692bcb65a1508f7a095a74ff2159e97a3c5c14ddd8b2c96a7a2bfe43d07e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1244d935c6db7b5441533aab87f518ea215aa6f5903b071f2ee8cb3359b3bcb2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0fdc11587841ff68e0606d5e9924388a5822c1f6f5c3dc2ef406e3af7ccf4e4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia7cdab2a88c99d9780bb267234b2cb87946009484d21f4419c50e7570438e645;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3245926b69b2db031c68574a86f56671d4dac371989b6670fd5cbf1106c85606;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iacdbe6e2ae2cd5fa475cde0217452a14f05bc8d499b9ddeca568f6cd96ad6a2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7e27c6552a8a17a2f1f9fa61cc6b4c478f1030f1ca44dcb98424d65cbf10f93;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5aaf6ccf4cefc2732732ddd816c3eb7aea7146c6e7abf913a5193f6906fe9497;
reg [MAX_SUM_WDTH_LONG-1:0]                  I37d8e18c384970e7a81bebcf85fe71c569fcc09b47de629e2258eee1c837ff31;
reg [MAX_SUM_WDTH_LONG-1:0]                  I96d8c1b67b028322f3d3e46d6306eac0333a8f3fe45073c08c5267157f73b71e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8d5e26d702af2d2b53b135bac7ec7097af7f878392c518c52571ead31ec485ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I600b1d1ff12460bfbaf32de67aff0e32087306628f0ba7db6736a81354309a41;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1d7ba7c6a56849ae78cfb42345e7510951e81fc92ea2aeb04addc6d3962e2873;
reg [MAX_SUM_WDTH_LONG-1:0]                  I225db641808b767d3f529e5ef2ac066e3abe953b8b434fd7bf4e02b57edc0f27;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8248e176e10a6ee79f77bbd56fb4f86d032c600522b20afc7fca399010fdfee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1b7380bca98b56ba1a2c2ad5d78fdadc1112b208e8d98b84c8d950f3f12f1658;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic35e7904ec654dd5f5e382f1df5d76cd1e4cd0af95a57ed979a5b369ed8ebdb1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I651492ce35fed9d77d5167dd211125ace0af8d55b8aff148e760d8919d53b6b8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I412c9dbea5975fe4fd5089a5d5b7e4270992142b7c2a5c4b59f2f6637215558d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id732b4b9de3f715537d32d6eb6eca4f6f9fa6d634bc283ceaef531bdef605537;
reg [MAX_SUM_WDTH_LONG-1:0]                  I480a5bbf4a2b6087f900087a2dc6c595ae36127a85d6551a9586443ca5c793c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I78c5859a565a68329d5f75effa2fbe77e16d86bbfcaf79d5480374f8bb87039c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2d42f8280d91ee6fed549f956ed81dcb31e70acdd0fb1fe4f63aa2bd3a7878f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I411faecc88c5a9fcbc433d784eccf7024675c9b009564295eeb765079b8069c8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia29c45f92e3672c1b0c186b711e5f0eba39186fccd95905a2bf9791609b8bccf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic429f74c6e97fa699700391c81e8a8ac449270476ebded49a8bcf8161a19260e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9572b18d2f9aa917168f389e7066eb543c9036fb55680d5dfda1e70b4d7a1193;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6efa3ca79fc64053e7e2744a4248a5c0df63ef15c66542967b53b2fcefe0d286;
reg [MAX_SUM_WDTH_LONG-1:0]                  I447026649273854452afc7335d4d52926fffb5950ed7a209f9f31e5aa95d6336;
reg [MAX_SUM_WDTH_LONG-1:0]                  I00827962c46c637f5d74d450ff4eae848b4cb15add5bf1f607708b76c8551c21;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb1f8fa764a70745aecd528189909af5082393c7f4d69462d6c069a011df5c6a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6cb1364420f9bdd072770a684de242f89990e3f144f160c2f5311bb00fe4daa0;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7730750ecb044040333f33232026110e55becb8df689868897b76fb093b5bc8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41bc9fc093e9f311e6376edb8aa0640709fb3bd420ff8a7cb2092844fbe0e121;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie2ed41aedb52e82863b3dfd580f2d2b7aff367f1613d274ddd5a5114316f858a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84519b5d45c05d737fb27ebd20ddbddfdaf7a22125df9eea17400856eed27992;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb92f51d1c0528dfafe1997ed4a9539f2f3d1b02900558ba6828e873a098789b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3af2de27ab7a899c5e55f150a53b7ef65e88309f4280269afb3eda2b1b408d05;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21742c373c52ea0c4872995841566c199318bf1f5849f05df796b79e171934b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I988d8e969e2a2ecac68a36a5f4eb0d6cb2c325e4be24c4716625070057ab9538;
reg [MAX_SUM_WDTH_LONG-1:0]                  I541077747787cf13e4c324b089049dcda6ff46c252b180e3d2c8f5b422217533;
reg [MAX_SUM_WDTH_LONG-1:0]                  I63ec7fce46bb02bd1662b19d58025abb479c4b57a0e4fd0642404ddf7f607077;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1fa1de74e664f3ed0ac923d6bf1a11fd74a6337f2c8f983d8b3dfe0f6737dc4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I086c1b2b7346139212d810647d98824eff245a9e24fa84006583fd56f1e76926;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3846e68c708bbe037e97544fc1cd70e7ed94539ddcad0d21984791ad35556d88;
reg [MAX_SUM_WDTH_LONG-1:0]                  I401154446147692cdd273c1d6dbe5a225e466799d41dd00f9477c586add460a4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b00e353fb14caee3c8e659e4c76b55ddaa6a17394c90f3fa53e52486059030c;
reg [MAX_SUM_WDTH_LONG-1:0]                  If832820141ab4f3c34efb429966b47ce584cf58fd34d38a7ecd976235613c541;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc3f186e24f214ba2d389536a913299116a402cb32c161f67fc854d73396e087;
reg [MAX_SUM_WDTH_LONG-1:0]                  If13409b9d8c65fe2127031b0e4f953f55c8a66c06811c6a5d261372aa2986511;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia86976aba4570aa0ae88d5ec887ea058cb4f7b49d7ec46b0ca215162564b1598;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2bc1d218fffb230a1505feb20cfb5229db9f3e2b0c7bb005bc8c59403fa35ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f93ff96a38e7ef38f5fe0f41333327e06adb0efc0ccc4c442058b75966ab5a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia1846f3088723131b0fc158b2d942749466887bf940e29340846070ac9d5090b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a2901c60b8a175d5462c32e4922a0bd931a186384b519b751929e551b477efb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5d5edfd68cef65681c36f4bcd770ec84a721eb515bc1d0fb7603ee0f5a63fabb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa5a98aa90cec881eabe5a6eee07f971778a40613c80891ff994d5a32d9ca6dc;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9efcedaa1cc036ad8613f9ba801ca4ff4afcd709f5e4aaadbcdcd130d1263fc8;
reg [MAX_SUM_WDTH_LONG-1:0]                  If367e1e075614957d2fd83c76b45a3ebe11f58723f4ce4f310646680622de4fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26dc2d992b646fe215751740a4406ce2a30e06fa2251f0382248aed7a08071be;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5001dd5906be258a2388828d2ea764df15f9efd4d2ed03ef3182e4ad7f3adba;
reg [MAX_SUM_WDTH_LONG-1:0]                  If25d531f7d1101b94167fde8f48549338e9b003202bc68bcb851f94fccb01007;
reg [MAX_SUM_WDTH_LONG-1:0]                  I499268c16db9bdcaf38ee694fa0269ae0c5ac8bc01e49cdc813244d8dd10c3aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e49103842dcd70cc7795bfb356ef7d178c1e87d94c08cbef0794b0956dff7b9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3f4ce0299be5d6b63eecc05da273fd2626ee66b8344d7cac0519c35643c8f487;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84b78cf1294735491099a4ece1a26f5a1bed53ffd09724d3383bc63756866721;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1894f875406842fcd82bee8824917bd78a61df725b719ed831ca04d6ee0845ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I964fe2ac03da8dd1965fd87a79f3fb2adf8e1607b64404233c3a09867227531e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8f3d1beef9bff167f3b3e18f1121ad15059b6030ace5b42de03ffd20167678d7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I58df6e4342bc054f0177b7c91a68a1afdac21b2d1d52434ef5d8272b92fef6d9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33e0fe9272640febb568aca8a4b79c740a030fbda58477f8c5314fe3dd6ffa97;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac61de7786d6ba1a40fc62f7d70b3cb366469c6674ebc4ecdaa21346903a58ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f8e0b3d76f589fcc9b17b95c68db92dbbe51ce063ef7ae57c527dae2bb92b50;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c94620659b19b26861b2f4dc674bd9b9ddd8a378f11b67d27bc0f7639e0842c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib3c97690b15aeae251f2ecc0b59366eede5e54cc23f96c5f55a04866d540dabb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4aeb03994ab1826b4bc249e1cdcbda394b864bcec0ca3bd6a0897fafa6d280f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia53a9dac8ef5ed6ca6e7d4a8e3ce09c23057963286442c6de8154990774e0c50;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d24219bb14476929c0d4b4bbef3ecee057061ad24af5601a8de67871680ee10;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8baa541fc5fd694b934bb04d8be6893f071225e454e095c6a69340d24c29abee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6729f7458757e512a921fff6abb9aa05fb498db59115c3b041bad959c15fad3f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47904cac869d3172932ccef3ee79eb5e70fa1dedbf4887d2f23fc54456756d7c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I543c9825f790b1e9264e3f6b5e66e64c773dd0866bda372b2eda0201910105e9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb2735bf9ba202c3ffb7d50c14e63bb88305bae465a10fd9df8e1a516569b257;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8097cf47b760092e87e117165f17e1f66afbaa3ee78160fd0e2a597f613883ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36abf86ea52d7dff510cd8b2223acc503829bf031477a5fb94f6cbeed88c1929;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4eb210e31e4ad434958f477b79dcf5b2694caf5c18f801a8d3b3b612eb0812af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb48731efd9ce27f84725ef47b1e6733a95b4753274e4dbaef808d4764a470e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40b6ad89db699e7f672e55f672bfc979d85a462330e526aefd63b9724ff7de89;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib45b2ba433dbdf77fdf6bf72c9e7a1b60d7bd8977c20cc9ae07e7320c058252e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I014e96c75acbbe2bf38e1c89b52e1a331eb3d31b984a67946eef2a5223b87855;
reg [MAX_SUM_WDTH_LONG-1:0]                  I30cb24b52e864de98a09fc41e8719f6009e8642027c70850c80dd90844b08093;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia3588e449670d7edbf99e52ccf0d7c8462b51e3d24ec5f0f7293290d47154f72;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62abc4525f5ddd159fd9af8e17f6b7a271d8aa70617eca684129eb9320ddefeb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6b3108db71d5eaffc5606fb88fe909a0462a77232258fd85cb6792954ad28c0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib5945692324b161750a7e5b6d9a2cba70565ddcb2f85ce9665da37e06c256ffb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55a1e3e076ea304ccd72b18524bfa076977a0f791806719d752ed020cb6c3e37;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3fc3cc1b4558877a3148d5567d5e5ef929459603af3c07214d2a05a5c9568e2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I318f0ddae7fd42b63d856ad6923268574eb4f8f71cbdddcaa420e917a1d7ea51;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie399b6c8ee179bfbefe764089dd280841d5e8bfa73941f40de3d7a293c4618fc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee19c6e30e6fb9258878db36251e2e15a071b41364b59473c9de2c0f0b8c9ce8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b0bec74dc25dc927944819c56c35d1df298227cb0fd804ca1b526db544b17f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4a9362c36b4a88ee5422688ee5550c97e8fe10b4cc23b6538ee81bfeef1472a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8007db0cf24afff18bc9922f5b33406c49079a0374944211f7ca69ed7dd8b4f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9dda3335af58c2daa92010ef90e217e0842b7740a65ce2a029ebde5b65e9fc86;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia79976d64cb4e1c9a542747c4a7ae62fe509cf1f8617cff283529b36e86464e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I996cd6ee71fdd8f4b109acfd52bf495951439b9e49b87a6db4565bebbc7d1e1d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5889799635ff332461bf6d25cf95f401edf86feb687d4013457a3298dd943c4a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I705cf789e535bcc9523034b7f4743daa8f66f1dfa3d15c77b87e9f1845563690;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3f8872c22051e28cc6cb6beed2ec233c7d8b79ed058acc23d862b30f0104715;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4345f323dbf4da279580851ea1d0b7a2e5109f518ca914c88b6ac91e9ce8625c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic620c07652badc1f7831a4e487498f6f875cc1d9c29604b1991dc89620485abf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8a484469fd2c86173f27a68b9ae6c15c3813761e5dc1035c2f9fe04b24a6d73d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I88787a9b8cae593784a9ffa45bb675bae477cadd18e0cbce021ecc9b4461dcea;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic6518d2e4de9b3feb98b24f5ff4fd43edb699fad33847f2e67ff731825f15177;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id093cb8cc2ca70696c70703a5a623de87427b286fe83fecbbe236110c68a8e8b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie147f013af77ffb57ecdf0bac185fd60648505960bec48f3f18094b1b7e319ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  I789fc42a39562699279fd510c6fe748b90314b0586a7e051058bad4b84370347;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a51859ca31f0b470011ae2b3bcbd11fd2c79f03c854103f016b54af79028ba1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae8a2a117b9f71a954b7368532a41c443d18950b56dcc9d12a7809dd4b6f9033;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1f5d36144836b1c2e41164adaa02934f77b47f317c3f6e7452ea483c756b4ba3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I386d1bd1bbf4aa7d9ccbe2cb4a9dbd9cf9bdc1fbccbac9039b32d0082f2442ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie1c46630d4cd6028c341687f4df0c2220054b63f8263fab4a11d3ad89f6518cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I588bd9ed21e23969799b7c1ec15350266ba52e0eeacb1bc20803f8aefcacab6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iedab2e8aa599a943abe7d0d1dabb0f7a5a7d4b97f36e982d5f548a4acccfe2c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7045e20c9bb1e7137b3c996fe61c7aad0323741b7b5dd70d8fe2ad840a816000;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7ecf5c9528425bf54c120398b0e5f75dcd4acd18b3088fd8a16fe8207a592bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id056954ad6043df8f15fdd039c5180035a585020638d2e39e1e1392e283942a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I355cc82d012dbfaa00529a9197d4fe0b654fc609360a0775d398ae0b3e95f2cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I213da828cb42a5d0f9025d51b36ddb92a677c7878c1f99496cf0c921bb8674c5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic0c2a03a257040df478653886a3a2400777322b4d4333c0da94211227433697f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I74a97e7cb539a14631bfc8532c9903e23e1889323443903126eefa3bc5e5be05;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic09079bc0fb0e140e7285e2e5af8caa802db98a774db8ce0bc5158e08becb4c1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie31f193f6b43563eb5a1cc4fac89514b8e972743354f7a28c0b6c8c8e70f1799;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia7d33f990e505c818a46c2a54c13bd6680e3a34847708d89ee6f38999242e0b4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a3a48d2c08ae2a07dc1e291c0d51c6e30be91af52aa6a439849005a958540d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0c87558b4bcfed105da91186dbea82b0f8d38c2473b578fb874ebd3e844edf51;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib93a5b2f4b149124dc2bdc6a90438a5bddd75a83c0717b52fdb47de0cbfdf8b7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a7f5ab868cc2f4e823808a238df41f5e29c98d896557abab5eb1b5ac4231eeb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76e90676f89b877e33f8c96e6fd6d2f1c2da1fa8602fb65bf8c1aa18d8b6269a;
reg [MAX_SUM_WDTH_LONG-1:0]                  If3574e7d834ff9a2b7247d3262dcd4265a5aa04a73495afc4e8098f7da4cd0ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d7cad2d595d0e7c85112d240714aa5ccb684bac4b8fb57f4e8118890ae82063;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5187aa2268c0345b27861b3f411a57adfe94104cd1a48c7573407a0f79e345d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia153e17a2ae12333c7982319dad7b3d57721e5e6075d2ee89f61dd6c8b06f73f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If54927516082a9fec583e3cdeaf09539203d2f351771381d6c29c7961dc6f98a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief4ea9c80ee182d2353b1a258190c80085fcd78a2379cd59968ade8f12695d20;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e63aa98e26c7163ac7e004f9b363177513859fd81ce1d6be355e187166ee55a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icacb23d3c6ca588b3fbe8371627f9c6de649dc63ec23db2a94d3b532660a8a8f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e3f1705d8ba2b2cbd6b7749bf249716ede50edeca032e277396a885c69399ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5902d24b66bb202f53e54816fccd38cf887dcd18bdf15dc6893dc55bcb6ad9d8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc29a95902384ae5ae3858cc3583cfc2fb39d4634b67c3c9858b9b6b9468fc87;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ife31d9500920174f7dda41fc67b6e54774505ed3c35a04eea45ca45b8be20457;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ee26418f368f28b1dbc386529fe4d0034170fceeaa1cf5f4edd2132db250ab6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I658eeaa8e533a4e2fff6e0c78b3d12aae697a38c0ae02a835e4c62eebe7d946a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I82393d9631be548b7d2f25eff102ffad6a2a1b7a683c82d8046dfd07b66e26a3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I77cfd243c2c2f87ba6a4f19612488bb84593524abb103ab9808275bb0a3f3c09;
reg [MAX_SUM_WDTH_LONG-1:0]                  I61291a36d4d546d1cb7c79a8a8c9ccbb4da2bf3fe853e05a56296804d5fde212;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2fc93ebc02fddfbbe5a6cf5bb7aca44f0a664be4a2c8273ac638ff7f94c3b896;
reg [MAX_SUM_WDTH_LONG-1:0]                  I454cdecfffd5c06b833e81e8990b07a9b326eec23f31a7b6589b969f610d8ed6;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8fd28316f1fd0fb493c897bdf978233c0a1bec3cf2136146e8471b86e0c0f67;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0d0472e7c0ef483f8cb46ed393b7bcd5ea93f12dc2885368d5bf587c24198980;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2452b31eb1cfee03ef6f6c00ed42126b741fbdbfd43b74377a675383e146ca22;
reg [MAX_SUM_WDTH_LONG-1:0]                  I33dc9b3b4f5aac0a30c5ab73b222441f5fbeedb26b7b8749a0ab253f239598d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2117d5fe8b672b3eaa3c257a2a7df3819e54d86ca29f980dac153f8a9da37607;
reg [MAX_SUM_WDTH_LONG-1:0]                  I70ea317892671f95b146604245efea2c83830d5e6b03a1dd19f2ecb28b47a9a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90c54ee94f70ae9ae84529f1c52175bf663de85a58c8ee420146322ee9faf1a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idf920a1de857f846c8ab2646a68ee3a6053d935968cdc3d6b46308a473be4099;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifdd6eaefa7e96076232a2d0f399e537f2eae4cf57a837693be785373eeb8f160;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifade018f22d237bddeb6fd8736ba424241846d20f2f32d2bb7fe779462ed7261;
reg [MAX_SUM_WDTH_LONG-1:0]                  I939c9cc4a14510cd9b1d69ec5f5649e80399a13c355e0f8bb8a5cda6df224e8d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9318e8402c23072dcc49ace45bb9814c535167574af63bc61463059dbcb0067e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8292477c74597003a879f491614abc033a2366dc024d96a5b38edc6517561f4c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic0071db5dbcb92ea14e4b31a24b9f9febc208bf86bb0634f07d9cd3763461055;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0e9f54539d4a95d17f80a316734c90dbf2799dd8311c6bdf7cb06d100d576254;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64cc4cfd27023e75e5cb557e7bac31506d466107aa2cfe7809e148d8977f8393;
reg [MAX_SUM_WDTH_LONG-1:0]                  If475d646e4baffa57990168021c33001ce2c5d28c7f22a83d42e35b6fcf1bd22;
reg [MAX_SUM_WDTH_LONG-1:0]                  I560502a76e2a6f15d91f55a12133213d8896b50299e0a7ed30c5c5958d5f5ec5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0122a25f242d23f81bd7c99bb094666594eb9c2ba1ebbfca379b384411257045;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7813b9f4f76a24bbf99a0f2d9cfe1d3a53eb0ec0fa5c72e06f1f86fdd1801c56;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id0e600a5ace87e9d404d63fcecff3d7a6b212ae81456381885943b78b98aa2aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia81295e4b9400e1737a8a8d335ed9765fbb59b817f0251f1f032ba3e48c6bdf3;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1febcbc92a43732fd85592bd9013cf0e14fd0e3926826badba0e53cbcdec1fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b7c06b48a33586be508f2334fc3eac5befd9ff87751db1859c5f01cc6d44b15;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id88407a8f20b0589f462959accb7d6737ae4c244083469d5207033ff09f7eb89;
reg [MAX_SUM_WDTH_LONG-1:0]                  I63860f7f2cc2e0814f98ead1e90694f745ef7a70e90f0af487d002ca46bf2c57;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0b7fce50c3bb3677721cd1cd0867a43bc7e7d172db559dd6e92617f65eb3184a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I48e0ff7c513e9892c552947f3bb0a96d7b00d0ccfa3d7fbcf067d996b3d58dc6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idba8e69c73d0fb1bd1aeff84e1c6d06234801f1b37b84ce20a98d29b69e98915;
reg [MAX_SUM_WDTH_LONG-1:0]                  I904078f4d964b6f66502423cb801a285f9cf21964df0a9fc1b8fdb9e35090265;
reg [MAX_SUM_WDTH_LONG-1:0]                  I204e9aa975645dee8af1ae12716c4c3a3a6f3884a24fcb113308d16a718f5f74;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaed17e55ab4220ad1c1485ce0b5e5518cfc682531407f36561bfff3ed5026ff6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I21423b347d172e9152d4a76123a9fb34cceae15bb211e99de5a3f25dd54b3d92;
reg [MAX_SUM_WDTH_LONG-1:0]                  I101c35283ea20516f74f90cdf4ea7f1ac3a008d80dcb4b80235a17483b1f5211;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c1ab87b7496ac411fe34c8295734d2eb6e3dce0c3770f06c2e61f1e9817f3e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1184b619aa3fb52506bcb002a57a421ae2f9d3a85502d2ae8132f38092c38fb5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia0a6c602c6591f708fc304b12d671520ec5327d8e45f7f066d24195464f454f0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I08fc2b9a844e2c482e2bf89714e92b5baa0ff2b9bc456c523d6360e5b5bbe2d0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia440e9ed203fb96d0b71bec0c8c3f8aa3ae0cceba15ab536fb4704dcb62e27e4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5617f2c448f426aa20d4dc124625b298648c40b73307feddaa9806bf571a71f4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f640efd56c0cd13cd6a2f7cebd9483076cc85b4668036f2739503dea91bea34;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic9219b1b4792455d5f1c104798cfb3ace66806e030172b83b652747280a3ea8f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If34c9fd9dd42116ff47c3db0a0a293a36fc2af3d8b66c4342c75e3c98bc969e9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia1e3983b6aaba9149d835f0e79d761b34c608f894259979b9e02f9891b0e04be;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5076cad6c2fedcd5c8e31e38043edbf8800ece300917426b42b72eb475bce88;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd87e183657088945b5a8789b001bbe566368ecbc0a773fb784a3d26cb6886e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c344f207e2150409498a524af2c7238e06c755329a5f2bdc5c298c2ad34d4cf;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic67c3bded52308b7875b1fe59eac4e253898565ad36a0f3cb39051d5a1a0289d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85328b4628dee41ae779fa1ca104a03dfdf089ad3ea8d7eede9a0869b1ddac71;
reg [MAX_SUM_WDTH_LONG-1:0]                  I496a0976329e8a4f6d29dbe1b1e9319f3f99afc9f4d3c645f264f4675b7ebf7b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d0a71f3a423efa567a3a55121fb24edaab598e2f36e51d7d2375c99e0554472;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93889e1f0f60b124844920662add026c1da1fa6650f347a6a616da18e8b96c02;
reg [MAX_SUM_WDTH_LONG-1:0]                  I830837e25b025c27a2e2957d7d0e12ac498d8eebb18bdea627b46c57ea61bf2d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9bea46de6ec248c77242ae2154d5c6e1dc17ff892dc903bd685badcbaf62291e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I802acbe8cfa680520493b84328e86b0cc0f5834df73ee11b2b35ed9997890e77;
reg [MAX_SUM_WDTH_LONG-1:0]                  I88a966d14bd155320f8f49d164cf93516a3822b9098c6417bcdb8a64f9eb1a38;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib29fb4c64cf1af8604b28c3cc158c13665bc570089df0e6ece0139f858aeada1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23c475c49d2504d72c81fcf2a1ca3122e6dfbc9f1e9faa0253d0d36c27881126;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5ee0d8bd36fdba065830db60c4511892d5e360e74ad676ce84ac82ba47d3e6f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib19a40aaae7bc965afa2506ee77fab296894319861766d0f6ede0e69e01ad17a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3e2780681adfda07b74c32d8a680f36823f2019a5f63c879113a2b258a339a24;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie10eac9c8e0f2526d443d3c8d9c007e29481ae4fd9bed2afac5a0861f80705c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I90657433c04f6300a3caf3c7aa1ea345ff62a9a5fd422d7326fe435a0236cb48;
reg [MAX_SUM_WDTH_LONG-1:0]                  I873fa9e73fcb148c0eab3dfc8d6163714e0a0dd5889d5d5dd73244c4f700f3bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e6b7e7d088f47fdb77cd0972877c65678f1d1e84f865a4f6a2dc3530ae75e8a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2d891a9027bcd15bb7deaddca0e282e872204770ad4e90ffcd4826beb3c492cf;
reg [MAX_SUM_WDTH_LONG-1:0]                  If50d96b50d6b829bdd534f141f7fd453812eab2373e6780f811dc8e43f61c9e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieae87e6a29536e19a2589665b2af980e34700c9a614fe1b7c4704a7a538a8f8c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I80f0dd7462a99f7863728dc9f513999e8df4d944672470fb4f614f0ab36b1bd7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia30f6d6396acef716d7383513ac1f4caface96330dcacfdc5302bbb0408697cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ad57caee3254be43c193b522b06af8f1b0603259b4c61f9db942f7d21afdb19;
reg [MAX_SUM_WDTH_LONG-1:0]                  I794ed9d1df776d692b623e89b6d6ade5d265c9869957ddd8e256061bb513d7ea;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97a181e9f8555a1bf3d9e9e1876e0ce599fa7c1fff5d905fdd14787e5b92956a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaaffc28ce6e25495dfad668af2f560c988f5a5abb76db94b71563231400c28b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie9fe82e8e7d32f0c47e6b0f9514a270018114d60c63841f864daed7f586a1732;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45324df36dd601c219634e39418995a9ab1bd58be03cb5dee89ac2d01bec1dde;
reg [MAX_SUM_WDTH_LONG-1:0]                  I28db4525c76b4ffd978720f47196c17b188839e095de0fce72cfaca9754cf2ca;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc26ae0a7d9ab347f3c75ed2ac7c48f6937f9cc035d46be065fb4b15699cc989;
reg [MAX_SUM_WDTH_LONG-1:0]                  I41ad0bce74c3d43c94ef9f055ff34fbcfadc63b49f45c24e3480735e706842be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8e22237e0bc0b24825cc53a9b88f0ad973a825d25aee1abcfddcbb6ddc14ea48;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied3eba558946ec39b989955200539b5593fddf4102f7811dbdc1fa0ee35d94d5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieff55ba27500b6d175abdc30224d7d4c703ff1ce6a3b5d86475b739903839b52;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0a0b709e36be096f2b7a9882b1de9c86a46b08e7693be36bd4e70082d5a7e1a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79948c8c3800c594e6e33eff537e1b38872775f3674ce78ad963f09de0091486;
reg [MAX_SUM_WDTH_LONG-1:0]                  I788b4acf11f5bbb2ad13fb9d931f593b149f2e9c252773e5044d8a9268cc818a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icf4362e74e763b339d2ba9634282b8441d0c293aacbc2879f95a53ef1a2122e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I674adba378ccde904a1bd264c3b6dc3f85faabaa01831cda8320aab4561fca87;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id6a3fad936fae13ba6503265a6a9a2bd1c54dc3fcb3d196623bf8aad32225687;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6039c5bf499421e601aa8290ecfe5a0e32552869e3222d6a881938886ee0e50b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic26999f764390a0c1461876b7687ee02acb7586ae1e24d171988084ca9d4aa82;
reg [MAX_SUM_WDTH_LONG-1:0]                  I823e547aea1e595b2a0345fc0866815d5195979bd55744098366f536832a36da;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic77bba83655ba517bc6313df02ee80ace5ba5e383e3794f971225d42bdf82690;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie728139df8a2d5d2cab83b4b4be5c462dd69107d1641666f7de5170c7e83d6dd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I01ac098466c350975d0ecff2227564446e39a21fd133aab22628a9cf3a866b90;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5e202ec46a29f008d78db131cfe4015f74fdf5a888f7dc1a700a94c5c18375c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97389ae6e03b0e2bee0e882909d2adf1aa34eecf73084ceab73088e850c24e87;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8df36cd42c3c76dd956f677770fc7b64fea6708efc711d8010a976ea719331d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I059c355ce17871c1a494b1a39b4ad3408ab5d28b886b143e04c71a29731f4651;
reg [MAX_SUM_WDTH_LONG-1:0]                  I020d4065b6ac016b70540fa3ec5d128c4c095e5b2f0bd807223b03aaeb730aac;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5a7256fb2ee0e45b0cc306c46856bd7cc606efccd221b75d515f608ad567603;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie79dee20ce2f12658f63bf8f47e8435a7993e0185c8c6a9aaf81a2f7951bc1fc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib419bb101d14a1958ca5b3a7c6a72d8fc15ca6e217fcac0f7eb84c776f3b0826;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8c5f6c0f6af8b9c18c00ab1116cb2cf9a93ec2f992be305dc553a7e858fca87;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie5a479b36bb003e0b2d92a68e955c1906c3969ee52a96b4aef5a84bc275f3f9f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7036a280bf3fb8f4d5ce054b2a19cc759ebf28fbfbeed38e6885b95899e1e4a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I380a702cee9dcf67af75101568b0a417c567c5ebc9e777dd1fd2d297c2455e90;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa80df411d8316c4d2acf8c1a094ba67ae97da2e64e440745984aff2f7a6061b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44aed07314ea5c6ed70e468558116a9b956c9a2d67e52229ac85b62c1b511d36;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d5d4c0a9031c2d7b9be5be76b42d25709e833098352ba533ad05dcb34571942;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f63700c8702ba858d076a1901ee015cd80dd29b33e109b7ce64aa14493461af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaeb27fc85e957ef3ea1cdd8db5ebfb513394c5f1680bd98e53b09552b554f80f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8bbc0d7554b094c7dbd8b4a06c4ef791cd6e66621e4c3b97464052276957603;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia109c552edbb715f4515acb56e6ce5edbc0bd73fe58165ed7cce5a35867f6332;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib65f0444b24cc43c4ebe5dc5fb7a2e0aad7c8d125bf92c527ba5dabd52d8f98a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie22b4331ce03a83f7b77b0ae01cf869497d506d764f6295831de5522518bfffb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I088890dd5f7391be17333396dc9b8cba40ddef39e657378c312707e1ea43bb56;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icd8816eeae15f7d5422c702821ce9d5fe0e272f5165cd7c6f100156f9cccca72;
reg [MAX_SUM_WDTH_LONG-1:0]                  I64fcddc23b1b1d72f4a5cd8707f8ec3dfb77bd105d279d01a99750b9ec4894d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2f34f393c20f24e86ee88f74da7085cae9c4df6d25b805f32adb16cb2bfc69b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I323a7ad384b7514bf52fc27d18b29da7effc88c35471be18c85d0b61ece11db3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I541091c82a0e29abaf2bb1c586f5c44501e90f7ac691f250690ff6fc4f186307;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iede33454e4e4f5856e3700d92d14d4b4ee573de70aa6715525cb1164348e6561;
reg [MAX_SUM_WDTH_LONG-1:0]                  If809f343f9007d972db4bafabd3a2c1f1a5d8a7a965cc6924aa965005763fcd5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6254bd01448c9d8e8b348c9cf6f62da72b3e66c76cfc692be2250a30039c48db;
reg [MAX_SUM_WDTH_LONG-1:0]                  I75b60c610ccc4ecb84b7616f74cf1cc68e4312dec53d71e99911cfc9f69ec69c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib50a67b0b1f097d85a05aefb1686e6d51cbbda0406226d20772af68de6e6d139;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifbb0c6db7e47972ee1ef163f0f3b0e8346b27ad9fe17801df9f1c4f9a79c6ed8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0809c22530a4fef601b75ff7573a7e9606b2da1938ed0918b43a958b9c2ddb9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied45ebda32de8ab6f352042b494f0350315f9a86a12bcd18991d3dc774876ce0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia0febef423616e7d4ab3957eea2ba1de8a8bba8b027652658ac2ab5aab11b9bf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I63bc47a8fa8e183d1451318367b43a76386d269e4ec267b71169127ad5c5a46e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8cdc972ad763857aa9a0cf1145ac106bedcf7897da19e06cdac06cbbc52e0141;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6a82ec3534f3eacf85d6fb59ea0a6d640df62089427d83d5a9f494661e44e942;
reg [MAX_SUM_WDTH_LONG-1:0]                  I10d197005aafecec4bf8c18547bda5a551dac520da311ee42db394ac67f413f1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I63f3c451c1d8566df035f6ebeccdf248343fabcea08423509f9caab46bb7a75c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb166c946a1916a593a1931a1651288e452553572b5b4e272aaa917a4afbc42e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I955d2b4663596b343e2ceab53a3bb73447741d4f3c8c935f35d72cf9b44249e9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3ca7faf1b6e8e04fdab54e1a4b313720f91992013d31b492f9aa49e54676aea4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf7b181b75b6f0fca207af49cfb93611fb71c31c28a5604de13112e8d521d008;
reg [MAX_SUM_WDTH_LONG-1:0]                  I77a2d0c0f26725cfe51712e4d1fd8663cdcd4668405e3fabd33e72bf7d008343;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6198ea973d8346b504b6da6f2fe193b989253fa47992f709c17ecf344f3572b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3c9445224e3dc806a499c5a5faae2cd5691cfb5497852d3aced39ec164d9a5ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2dda176f6e7f4c75b5cb93278b95ba9bd30bda61c0d44c103e5092e71d4db7ee;
reg [MAX_SUM_WDTH_LONG-1:0]                  If86de9d134174799b06582013809be1a492e36de3aeae4cab7bdd6a827223976;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8578eac4c908240f9cd21d004858326a5c6d88ba020a8b0f27955896bd227e30;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c7e61c506c8d841d4747e5963d49e0237b106ba6cb15a0fc9e4680ccab02c5e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ce58155e37948ec0a5842ed20258c382c0fd9889e697912d1ee1018a5e25d74;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c17caab5e5aed3ddf7a867cf514cdb5f65c3591789f1058a756265f97aabea9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I13016deb611dec6abdc3b14008afeb343ae5cafa44375dcbb1d09da08c80cdbe;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic818ff3260f1543c8d940d36c72d644a7a3a243220548792289117ca6a793c02;
reg [MAX_SUM_WDTH_LONG-1:0]                  I046da9b39f69a49ca827ae6c66c4164d2c64cb390dc8ccc238a70c68f00e29c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief965ff00c0da0a12a68cadf50622567e99dd688e9bb810dd46f69e3eacb7285;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic7d0c1eb012c5cf07f8df74a28a53ebfb026d43c9161bd7cb0de0fdf8bf6a9cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib4d1942b7949b0a4e79441e13e3b6b7b36bbb136c2bed6ad1adba30a840f4b55;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f53d47b7607b32c4f7401fd9fb07a28d9dee9a3119dbcd0b6f09292a910107b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc7991125ae81f1c0d5f221c7fccd90e5aaf92e72e0421aa687e6c1e0f8afa9d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I46c1d6509155e8a243b0d4fca0c08cc86e520b8142ff55887efd0b27fc9ec619;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic1e2fa322b42a15a886ec6ba9f67656a39c8bd6a13af883081336da43d9d0406;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8a41819311f3c31efd56be044479263c2afbb88f7c90ebb8ad570237506878b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibdbd014d7bbe12aa223eaa43939e3459f35b9970ed075d4733932cb66042d281;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6c2b8dce255f31b35ddec9776805ae6b3dd2d4d843a755375f49d28a7f7f6d8d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4dcdb2c22db70cdfa468f9249fea4262e91120e0d995981b34919e26c9b5bc5b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibe35c53955eeba706ea61cb7d516b391278b1e27ae1eb5f796d45dca20a11928;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2f6966ba5ca0aea5cb187d9d90bb6b743b80bbc7fc4547396dac13a22603e7d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4df41d0da488a9cf1999eb318b6654e68637641f78ce9be4636203d6dcab3285;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibec37c7599a7f7cad52a48cb44ea0ffe117ac5ea206590a3eb8a2c661913c9ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I79c3d77c250619b76005964a5d8b3dc5480c395f1b541d7234d846955213a0e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieea63392582d451f7570a458bd235afaec2d11a7427d4e706bc1d73128993792;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0997b7b9813944c111e41c7f375c0925dab34b604959dfdcc8dfcaeb701d6d62;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2fc14612ec75b59c28fa90d7a5bfd1bce6d5d1fe0c46ba45f77ee2f9aa9e481a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie6e358691e81a9c1ca0a585b69352779f083e4f3e26d03152194b1a9238f0f0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I876dccf88204e4113c5f80bdf348624dfbd5a1439638577670da4c6afe1d5f70;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3480800eed0a0bdd9a7131caf3ce773b28d952484926c279b3a5e6244925a6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  If0c1eced668b91b966c13a44ef09ca1209f96723c7e3d030a757d45d0b61141f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ddb5092da74c5ef9553f80099ceb2798e717d25b24053400181825ba303c5da;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5f3fc42a6dc35a49dba82814b80238d6a9f6e9c8cfddd4d72749a3197115b969;
reg [MAX_SUM_WDTH_LONG-1:0]                  I552b1b2def8af8685711597e1db1da516b0766591b757ea9f33c666f9e243ff8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I677e11f6dcc443a45cc24e28c955adce7dc006e6b26e0ade792740c59d91ed6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia5703a4566bd7f99d071749104ecbd4712bda3f156cec8a1c4d4d40303e37fc2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I703d9bd8f5b9435c814d93ae7e2327a45e0febce37b67b770c2b93f30ba39972;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id5f32d64dc52d3fa4da97ed5a432d520af0cbc1e4714d57788e668a7bf3fb310;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d518a62a0a46b493ab538e6ccaec00b9b2cd08aba9695482997b884ae7b006e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9977445235192d6416fdf5221fac29c4586af4f83efa91e128a0cc18cf648281;
reg [MAX_SUM_WDTH_LONG-1:0]                  I67fa42eadbdacb43b464b7246fbecac6c261d3cc37d501efdc1e83b9b1ff6055;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5fbd149fabfe16474e75301b3ec4e0ecf4c70537882f00d8c8fc630e7656b368;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb5ffff327b8edefda5ee44436f5f31deac21a01781b65e2429b1e1a025c997c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iceb61d5ca2b0e3fa972b66d7215d7e24047180d638846c80cba9b4e84e147d49;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0384038afb05788ee28f773a244ec49cd78da115f5d864f8497df2b36f37ae54;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac3ec84d526a71f93a304493831b4f9597b2ba176aea1b62dce09eebb9dd0e4f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibee29fffd6b844b0fc4666fbb35c295ccc5a7b99dbedce125b370508cf6b0b90;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib6afefc545bb77d065a44983762a6b83fafb326b323fec8946ac2f7b11865d26;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8f9f47f8cf0ac244089271b1cb952cac9d90aa94b91eef48733afbbcd992952;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9781f084a762fe71955603c76c6d57791f2a642ab73c8393d5ed79b42dca7b66;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie80058ecf96cf544095e34ccc9662fb679b8da3cf6f10797805cbcaddfd63804;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff4386a737586e5cd21336fe2f577e54c5c8bebdca0c7fb944923f8a9ef09d2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I680b7384eb5b44faf98980956603d7db164a819fe394beff4e94872edcbece0b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1ebcad455793356bccaa94bc33207b868ed70c398881b3ff78c8eab610605708;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7bdb6b57635075a7bb8408a878d4ef7f2ff136804287cfbacddb40bb20dd053a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I068c9d5ac9f999a475341bd2e8328de90021df28cbe517e182ad5de16d1a0f51;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27f0b66e246c474ca71e1ae20503843b31921b5552092c5ae6eb872e76808395;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1524d287bf11b9e8bd9c37a61011f3d9a6d18bc1dc48aa254cf288134bbef748;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id81f3fed6908e777951bdff6448776a9a80348c44058ba0f9450999a26f6155f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e88cba4b7ba164003b35e7b7266a2d22b85b731144db715c2675eb9011bf01e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4655a76ed253aad70f2340070cd7b6f2041e6782a87be16ea66ee0fa2e2ad74;
reg [MAX_SUM_WDTH_LONG-1:0]                  I18edf674979e3ba4398115ff3e5912b2a41737a1641df1ab7c7539e10cd53785;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8acc445f4b9f01af1a8f4f34ab10028472b79a2c1d1d3b8aed7d040f5ff4cff9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib8387757c67a87e7a37c530022a9539aab577c140512fc5481f00fc9ef52a140;
reg [MAX_SUM_WDTH_LONG-1:0]                  I11f1c07733856926d4d980234959cd48f8b0247270d6485cc57dc3456ba7adbf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d2bf12a647b50d4ab9b14ca939986eb9960c3019be93049f9086529acdfee39;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26f2f2938065d9336a83a2edcb5595f6976c5c434c76d4c44e771cb8a0c685c4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6648e8e7f5ebb09e748ceaf1dff7eb3cb073b8d035948f93b25c45bb10b2589f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I059b4a33ad6774feb79158ff05ecb4287420d94dc0c57650fb90f11fb7fb83ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  I248153dbc85025b19e54dbce1436968e1467457e71047a73fd6b1365aa362259;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a9e162c226e402630bd217ff502dc5aa823ee7c089801803c5ee091b5ea4026;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iebae6187f539cafedc0df54b1428bc9b57c6aeb3320a5bdc212d444a9a4fbcf9;
reg [MAX_SUM_WDTH_LONG-1:0]                  If30f29822c81c32a3f153165fbdd82ff6cd9527a6a065627852ca8d5d1a0b122;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9b9bf6eb31652e7b62bb383e61221c03099b628ce1f87617b7c90805088c161e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iec9d3d3ad44a5c22fbedf1fc73a01cf348f8c4b16c5f3f0cf55c85f8d92ca22b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8b61d2b7d04b31046b959b2e56f86603abcd13532e8c5d7496b769f872bd6fd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I94452304db6f03a077cc46cd087cc756c098f85885a9c8a60e1860ebb0b23a60;
reg [MAX_SUM_WDTH_LONG-1:0]                  I294ca2d54cee0e207eba2b6bc501af13d7576edac3409f1d345f26fe570947a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I59d79bf88b865cc38882adc0e8d69f2a1556f9cef906cd558730ea7a902de6ce;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee74dd10fa4b539456d95de7258116aa77db37667ec4ec2decfa968bf6f602aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I022500b8d9cd3b589fb75b90c1b633a96fdc76c0e3e2ec514cf7b4ff3ccce1b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I62b9c19449f50c6d47f459d20978c10e564edeec60593f2213ec4a45203a9b93;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9936f1014242296259237c4aa19452ea56509e2d970ce60c72e7c4d18a66752;
reg [MAX_SUM_WDTH_LONG-1:0]                  I85c9fd61717aec721a675c20933429f4e323f13065bcdbf79eee199d97d2e56b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idad105c150f27de4777164385ed4e2123966f63d2b2ff32add6d18a95be2624d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23746c5cc5a886c61f469589a55b57fd6e8b77852b50e814c672a2c52802f253;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice1023bfed1f964ccc66c7d914378cc899ac310a76f3d694302cc688bb560e45;
reg [MAX_SUM_WDTH_LONG-1:0]                  I806e92d3c392bf729c0f36bdc2b5d398ef947f073dcc733e4301aab45a73d08f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I372b0e45c0d1e8d30830bd3cac2c3082ec36f9af195380d0e1b7d62712123fa7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9fd1bb95c6a2213084ff79a560a6264130dbc55ea0ee6b2702539e00fbfc67e3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie98369c31ad7be164b6fc0f16fd6d1a5193f2b00a3eb10ee1cb478b4653b60fe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6644cc3a42774e6d8fa09e46158d631bf6b48b406b7981f8feed695d22959203;
reg [MAX_SUM_WDTH_LONG-1:0]                  I80f30106eccbcdd1f0aabed1521d2b09a4bb56a421079ec90f81527a903c6643;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iae221cbeaae99099c7066532f85d20ecf85ca760a449bb238696d7821a729c21;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81349ebf72720f77a8902dc12d9cf986ddec6f8fe30f7f76f9f4dc54881708b5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I304c658d3b58023c7c85b82e12d5e4eec7336cf6d04c3468e591bb77e4cce5ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic941f62ac4a004ce3dfdcdfc5312a3be16a5307024d1ad292754532cec3fc90b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57d74f096ffd259b46eb1b76f49ec20079d2b15d7453108f95f5f6aaf6a272f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I65c4ade7c4c23e62f5cd1846b0a739c70cd498087298f54c41f89bbd9677e705;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7e4b87e71ac1fd30a6139a3cf27f76002a1c67adf28eb8d4e382866afa224cb3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d548bf4a643564a906a42a32acc4fe6919c91f43890f1b921b9e42100b92e68;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3704a80d3cd58a300a6e4d721e00950f5166111d44d9827c6b492524d4c556c6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id89fd01703e5a1c53c89a64885698fdf565b791620408fb963b53208a33e7f47;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4e750ac2d9b11787d2cabe2f06aec65d630b6be5185d7ec5a3efa12565000e2d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8467f29aa6da06588468e21697c56464c67e4809c135d2d41e38d9881715aee7;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia2b84466a2783970d94e38c4a99be0bd22b7e574580adb621eb579e8f9bf81b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55ee374c21e5aee6b0ada78409b18bdefed20abbf3dc5716c62daa87b418dcfa;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied4d22813a35e4cb32ffd1cdfddcdcc877dbfc83dd6d6780296ec5c5c9960925;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4285be4ac50db4da7f720fe115c342ad8ecefdf6dbace4af4c9714009ae31e86;
reg [MAX_SUM_WDTH_LONG-1:0]                  I11bcf52f915e80d94647f8fa66ee0dbf0d31537d68a896fd62b4fdfd8e76aee6;
reg [MAX_SUM_WDTH_LONG-1:0]                  If37e3544f587a047696dc53e30f6031f848e27a13e2328b2c38a4f51421954db;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibc1d752fb7dc31452424184c390d0348180fae8b0901eadef67aac5bfb0bc449;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id9067d2f353cbef30dc828f16a97436418af2bf3e5fd19300471de394f710fff;
reg [MAX_SUM_WDTH_LONG-1:0]                  I26105c08050f06741f732eb11726ecee4899cca05c21e1aa75eefb07c60b695f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I93150066a1cfdd9e59edd1d42cd2611eac0df4fdfbea33d913804f52dbd895a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib75010a3db964882380071e188e4d75235be279058fa470c1a758a97a7ab518b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie296c1317a499d9d35191ae9de6c681e2b521a2966b8837ffa470e3de6c8530d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I32d23e06facbd4ea9378cd4d72ac744cfc0ddfc54bb1c22550b09176ea670372;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0aecd8795e3571b4b428903758f7dac78966a9a928f64c26a3e6f00fd61872ab;
reg [MAX_SUM_WDTH_LONG-1:0]                  I84baca35ef199aa658e78c93b7dd27049c57dc70d92194ae59ae657ac001470d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0bc6fa0d581c2d2fcce482d2821bf87f00bc84606afa8b56d7f4cd88bead4a3d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7cd8396ac94d8c37d3de99389d6b06115b7d36f1e31faf88cdf01c5662fcbbed;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idfee0ad9592b445c7afa92c1099d49c458d1eda5605ad06e6ec975e2d9103e11;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47f3b89a5acb9ee2c282930b7d311145f48b3aa49a1ebd406b76412db2042fa4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic700c1c29d2fbb8e2e85fd9871082303e3dada09845afca88fd7c35f9d41affe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I40748060a17eaeb7d8f1a828d0767e42c09c2c104161262b5adc72249d128df6;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie1342b74cd710b1a52ba3de5ca28ee42d03eaf53a42a6cedab9ecb6d987d7b55;
reg [MAX_SUM_WDTH_LONG-1:0]                  I580aa2ffd81e1289f84a7d86e68cabc547ca6c8bb698bb648f6cf57491c18289;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69f8afa3d9aea957a3c1a9f3dbfd8ef8dc6370b228a7f67f0a27113c094992ed;
reg [MAX_SUM_WDTH_LONG-1:0]                  I89baba2fe1581baa53e6774b196896f7a0c32f88c5dcb0f6ccc7cd4911992b15;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3b017b72afccffaac4ff923e52843d312e1cd5e1123575d6daf4692f81cfe748;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2e381e0df584249b04ed891c499ded7e2d180a403ece202bb96f3cf8041dbbd8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I100b4afda393740a5fcf563e8e5fe34d5d7bfc439f2eedd77966bc9b37b3d602;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id539ba7ee7b26dc8f610a6298e8fb42f50f810b490cd75ca72f0875a2271c8b3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieeaf4fb83c3c92f18b21f65ff2a951f74693fa6da2ec322ae6a4873d26729f51;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9826aba6d5de9618406c264016c229e048ccc60817b1edccef930d6e6bfc6a0d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I27ac039dc48350ce90d2a8a3953936d5f7c97ec1098fb20d853cd062f2d4a6f9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic211c903aae638bfcdd91aa6d092f085204dad95f7e45bc78c9269816684ce42;
reg [MAX_SUM_WDTH_LONG-1:0]                  I224433de24984b12aa905ae86eeaa53ec459acd68fefdba7aa1e8778abb89408;
reg [MAX_SUM_WDTH_LONG-1:0]                  I14d3a54a6919ec76c17e6d155fed5dd3848ea7e567f997f659d5a09a2100190b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice1b30668532ff63b6ead40f37366b805ea21a65f6fb7067bf9d3b5d08eced46;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idfa486a97bc44780268cdfe3738e6c0a3fa58e51f0c4bad523ce7ab24b3fc471;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b6551d9c8b14c787afa552e23234fdbb63c8fdb8fb285416ff1b72a38e7d898;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib486f88deb674197e70cfa4b28061cca75c06176b05673ded7af5c62ffe15d5d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24ade58e2190b73f141a858e6812d93a49203181d6d427a29415d014a9cceec6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I958b582efc12bab546e1da193b5687e5c19e401a03bc7d6fa5c7bb1108ad911c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I55affee832ae4e480ffb916ce8a5e3b12fb6429f1ccee3a8f9a668aeb8352f7e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1fd2d5d75d3b779da0e3e1c3c66053704eac857ecae818b79be59c72e04e0b92;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3f2f052f1d132cf1a83172a044968741665a7b85e421658976109057a3d00ba1;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5f8b823e2d28fc1b521af24083f2fa271ac7a29129e8cc1cf8c5eba46fa4583;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibbe3cd91dfae5930a6ae5799a27b045ce6e0c59fe00a38b5fb4b1691949847f2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id068fbdc476f28f1695939e90fef8a08e2cd9434b1368ddefb14cdc950a76a2e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icbbfd81a7f066da629076f9f7c26eb457be34298a6518cf45e67bb39e74f5f2a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia193fe333281870ef7d810f61721dd6c5557204828bec993bb47bf37c9ab46e8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I762a7e10d310500a1080b7b46a9a30bb003c7a7d48011e96501a647e1de0cb66;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifedd253513982e9c918cb3e4a65f4a6034759bb977b8dc42b00ce4a97cbdd5ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idc9ce24f8fd9ca7372ef25d9e2b8414a4c8051c796f9ce64b91a6f3e70faeec6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6ebc1aa84acf73083137d13ff8d907175d13ac8031ff97e186840f851182fa28;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iffe887b6857424a57f7b7bec156197556dd869c44a2eaa660fa66760cd88888a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d39228cd05d50c7151740b19887493bd52a4504ce3b2090dc14baba0b03affc;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie7328907da6b377ef494c54a5e6fc2f90992a99258967af4bc2205d0d42e9db1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3369e19a0c3d22229db15bfe65a56d3f45222928f405a8c28bb7dd5f5f6a96a1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I98616ac468624d04fcf2487684bc23bd20a87b719be4d4533f987ecb1bcc8d5c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6f621b228fdc4c92d7bd7bcdfe69acfae45c715d228e99fc566de1e72163faf2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieb0d5850e57aa2cd83ee69ba71c85e9e047a9cc5b195da367a9f042a39559f47;
reg [MAX_SUM_WDTH_LONG-1:0]                  I86236809a2da5af49885cd9a573af96295f9f16b79a784c7803681cf5494076f;
reg [MAX_SUM_WDTH_LONG-1:0]                  If6bf4d8f739928e726bca59f6307a2b78966853a5aeae6bb7dc4786660382ad9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0bda102a3a10c710d14ca95940f86071834d6ed6cad335022b18ff8f2cee8602;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3fc232b4e4ad45bd25aaed0b1306112944d63174fc4f473899349954e94895cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I00dc832ce34e281f748daed4bf56bc03e171d8124f2c72f7627ed6a5004de894;
reg [MAX_SUM_WDTH_LONG-1:0]                  I07c430087a2a880f756db41ba39cef794ad6d3b28723a7c22df5aa719bf585c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id5fb94774f7af4bb8c727a46f588f1266ec3fde633c58ef0844ea4f486782842;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff963f656b33e8c5d0b4155f3d4ce0be5ec1c056727223d45af4ae070b006272;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7fb0278bccf79ccd873d9a4bb72a48982ed0d6c1a8702c009bde652c84c90acb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I44d78165b52487e966d2063495d2b76b8086031f3d3f0bac7713717f1e56b721;
reg [MAX_SUM_WDTH_LONG-1:0]                  I345d4e8e18ce7ca6151e381d432ce605af1865671c5aa141b209d1818e2c06e0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6e5de0450866fddb6d15781d26a3df126ea57faea36d172ff9c08fbed711ea47;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b2c44feae2f93582dfa6ceaeff78800b79465d7cafdf52289855eba9ba3a236;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4db811b4d839e478783694d956589c702666e122689ec06c5fcd299c782b1a7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1d109f4a8531b0b430e5010ec4e2619c94fa8502f3979e8450c9b1d09206660c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I23072d2753b8750a9cd8da42f6ec9fdce24f0ccf4c201e983c3aa96963421ed3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6a87ff2f8cc2aef5244068df9185b2f8a6b899cf3e6ad460439150b1f2dee99c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I96d2ff73be5717714513ef2406648446833f53abe34481e91be763d63d3f2d09;
reg [MAX_SUM_WDTH_LONG-1:0]                  I645eb770871cffae4c361144a6b3e428d61327c7379b25e3de9ec083b7d9e299;
reg [MAX_SUM_WDTH_LONG-1:0]                  If7d7e9843a2eed7a0478c5991a13e140b1ab83460cc8ea6a3bf24a85b8d8ae49;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1fc6e041dc759bd5cb34a694328c83cce92d4169f00f674238fcd140226fb7f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I61ea75f5f583a43e3691ab2462210c213f53492dd6a4a0a41abc406a7a828bd8;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic803fc5440f03ab206425c2100f94823b03ff2a6d6c238ed7407fdf71237986d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2668038e4b55b5d2fbdfcb8fdc56d43beaf4546ba92b39940b8f055a51d7013f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice1dfd35c5faf0569fc1f6572561e2931d4616abed72917aa2f79010b9949786;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia29b333453d0a00fb718748060cc9eb198035cf24697fefdcc6b75b450e5fa6c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida74a7b5fe7355a18199b5b942096f1655f787e2b340aa6954243923045f59a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9c17b85d3c4d97f0a7093e8007d812455859adb691cd79d2e41e78f95c44d2d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibf7568c1b00603b724362101a10a23918bd964f364af6cc21399eca4c9a7f17b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idb9949cbe1d38f86e61e1cce9211aa264e0abfb2ea1afa05be251144a4a081b1;
reg [MAX_SUM_WDTH_LONG-1:0]                  I636a373b59d09734f347126322958163d4e21351a4fb1f1acccc9209429fd38d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I18216dc1eb7be60021a2be1d64303e6b9838aaaa2a9b1e6bdffd2a3789661432;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifb235b2a210906a94a1dd95f01a9adcaf8fd76e786707e99bbfa8f0b4bf36e18;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id8f0e532c3fc4af615d6cf0967f8a54e6971c1f3572b4383c25360f5f8204ac3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f513306dcc73f879dd824e41b5335820c03331e576edc90cf579cfeecfc74ff;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia59883b6b96f3bbe38c2326bfca00e25d3b596e7ddf9287bbf70107666855849;
reg [MAX_SUM_WDTH_LONG-1:0]                  I54e17ea4294cd67ff4fe7c421e38999b0b6c6eaac95124d86c6f19863061e935;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied4edbf18ed0371b7d1ffd53ca5d98f1344d1640b4ca9733d97af5ba5c1c2a5a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I122b25621999aa119574ea30fab73a0dfa43bb5da1e0e76082f0844cad371a4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  If9a4d7f44a518a3ab1ecc6bd5d4e05d8e8f78615ebada754f1ef1e7b13a0e956;
reg [MAX_SUM_WDTH_LONG-1:0]                  I32549ac0c631e47367790a831498738385979aada71ed9fa5d238c4128be632f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I53fa59c42044794f03f617ff512486e58e173121f75b8dc3eb292e9246f7740f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ba7035cb5eb95ebff5d5d7e549a4ade921979bb4fa7e27f5810134ac2890d2c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9ae27a7b654a36e4265449d861213978965e4cc3bc7f36b77c6a77cde5e24f77;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic14e91de88b33f4702b25a3e0b4485ba5165438366333847b3e2687934315ccd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9dd84c850b5e32710685c595cad935e3249afc0132b04ad8dec94cf13e16faf5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I119671afd256f916b0acec0f5212868cd2dab6bbbd5b158a5fd37320253cb913;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id59c354fd382f5bb1b276d565cfc2a0d55444ebe928c144c3d0b5513d53e3787;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3350bfb01272aafbeca7b9bffcab3434116b885a4ecc32cd92680d122656906a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idab4a7def7105c2e615a9138bf503482df9a2c434aa1ee7c4937acf6d0e6bac1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifce65e25bb01c5dd7349a1766ec452a1658f643d6bbe1f877493527cb46e568b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0d0ba52491ed5f98c69d74967cefc454cb2be9dc40bbc5bfe16c8ace0231dd70;
reg [MAX_SUM_WDTH_LONG-1:0]                  I000e12e2ac3967d4da10fb33efdbb5d6e58d70ec6be81408ba9b7a0995925edf;
reg [MAX_SUM_WDTH_LONG-1:0]                  I05291a3275d232592dd880dda626cf60a03a62c655a2cf4b811f5325a07eb5e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id202333f4219877a36045cd10102973d3a15c1dc91156e14961f1d09744c6a6d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I141f0199ad8f1dcd707f6b0553ebd7fd04217fb960f13cf25e98511ed91bc7aa;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9a92d30f7a49d8556b1c480dfa0ab3a0dfee73aef8b8e5caa76e25a3df6742c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I11a01802ccb6a01458a2cb2be3dea2f663acc531821edd809b95e10fb5a2def7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45ee0619e5d6be949b89b7356b7d5a6c42d33e44c5a8885fe69eaacfc56ba8ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id76b3104f5a076b0f43f85da8b35a62b36a68d76bf8f26ff0667e085b37ce0e1;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id94d619696cf4cb1820576796ffef7f4fbe3a8a300c5fec44516ec9797164636;
reg [MAX_SUM_WDTH_LONG-1:0]                  If5b73982b4248c4d2cc32bc28f0df8b37553ac0b034c0ebe3009bdfee069f642;
reg [MAX_SUM_WDTH_LONG-1:0]                  I82f65771b72b94319cef82f095d5719ff7dce631f5bc2769ca69634c978bb4ec;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9e3cbc961652bd76ec24ad12037b6384d8690af30372a8e0e5a93c57e4fb7b70;
reg [MAX_SUM_WDTH_LONG-1:0]                  I6566d75140a54ab2f2f601ec74a46508751ac02ee7bf86bee304dfa07d54c8e2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7107302bbea73f0e5ff5ea2791a6d536cb04a165b68ef03ebeab0c0bfffe92cd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3a570d5967f92b4061a618a46c8d71292ae290fc212c5e3356651a7a69c22da7;
reg [MAX_SUM_WDTH_LONG-1:0]                  I561f05c657c3171c43fdfbb59215727da59d919f424597533b1890f7afe7cf07;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id348d892485f4cc1abbc4a897aef1fb7fa4f27c61ff633c9582a1bf733f5d55c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I81789766f2008122a36b608dce3f08425ac203a154b4e43f915e0e3ef19fa022;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0697f4ec5a674060a0fe012ca040842a7e13ab1391df2b3d09398a7ca857ba3b;
reg [MAX_SUM_WDTH_LONG-1:0]                  I678953f2ad317e167eea663eef2246d68cc67776d905877573ebcc39188a9a4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifad69639fb069c42f4ba17d17a3313ac3414b948dec1f6ad011824925fc5a7a9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I048fdd325368b2b72c83a32e9ac2c0208f392416f178445db74ceeafe56c8408;
reg [MAX_SUM_WDTH_LONG-1:0]                  I604729a7799bbcf6bc10010a36ab4d0bd909a52c6ea58259e7c532c28c19b1d6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I16b1a9836d7b38707938eb48bf60f17f049403d2fd29d5245798fd1ade1c2531;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic42634514b28215593b2b52782e8b58dd3f1e9e4276619e8603c5de34b4acac5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I48c21b6fc24c93dae3a01b55b280508297e0ff5101c7fbc7d17e823d9a31fb07;
reg [MAX_SUM_WDTH_LONG-1:0]                  I78f9a0c586ec95915e1628e57d58d38942d01562658ce91c4409571459bbda96;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9d5c1ef1f35b4d40b4f20dcd2c33691152683bf308c95aa53adbf785defb75ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I18c23544d10425853b73e8bd64411a829f4bd9fd145e5352cacd6ecf0c764945;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iec1baa5364573d0a9866494a039a3409a32b4665d4a79e2a729b54d370ecad97;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c79c03f571f276bfc03a16709012424498a1d7d53208213e600cd300cfddaf6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I508c79d6f4d56ea0e8100825c438214e4b5087004f8a5041b4beb900509cfde8;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2ce3e228247a767e41b5c376457e5be0d11aaef621b0d63d7683741f275b3f4e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id55510ec558d15440325660ab2ac2cd9d4dd682c082479a742118c9ba1923cae;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie00142d305ce51cc78575481f10dda9c40010d6ae4a3fcb4435961983c8aa98c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I000c117a768755741005775b84eb6e4c406d2e29765ca9bbab991217963de8d2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibd10325e424f3c8f0a460f2a4fe7bbffbfa3bc23e74abe4dfd6ec5b278e2c4be;
reg [MAX_SUM_WDTH_LONG-1:0]                  I95d510e99cd368229106d7ef60f9438bc186adb5359c9483b645b255a769df90;
reg [MAX_SUM_WDTH_LONG-1:0]                  I47c4e3e3263c6533efa2dc2e7f1ec4150499e8360e38b1cfaa524071faadc4f5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4cb9b54295972404ff2984e0b2a225773e067803925fc434674a5ef2439df4c3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2b48e805b3470041470bf0544dba31d75214a8834e8c456aebb8dc5a12e8656;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ied36baf05b90f7d785653eb1e7f699cfa84cd0a1eb3a985047f57e2885dad2ef;
reg [MAX_SUM_WDTH_LONG-1:0]                  I945dbc06fbc44959482d5670747fc5c6044a790ffc0a73ca0f41f150e8d59056;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id3947617c14deada0b43f71b47e700dbd8a1ac15820eed783d58774c249d5f24;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7d3a0a0dd3aea84fb203c8b51f1e4424f287b9ef01410f3cc5ac7e7579f2d4c0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I846f9754b91cbdf37fc2662d5851bfffa4926c1ef01f4a23f20b02d9588ff3d4;
reg [MAX_SUM_WDTH_LONG-1:0]                  I297e0d55dd6607cd32af52aac3e610ccf0fdb5e52f2ba250dd2c929616a33a8d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7485137b6eb30fbd6f06453139f9cd1ebeec411e566936bc598f0aefde881251;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id4d7fc501da443ac562b3578778aaea5dca1938dfb4563d14632481d1f453eb3;
reg [MAX_SUM_WDTH_LONG-1:0]                  I152ada5197e26088aadb2058a128099d201dc6e91d564b80b8e3930567a1a929;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8aee3ea7ce652159455573562acaad5e41a877766e7fda11580be1d60194305d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic86eed327a12ce5bd475a6b82a5bdc31777526455fb541a8f4e842605bb34ddf;
reg [MAX_SUM_WDTH_LONG-1:0]                  If787f037863d4eb15f1371255724977e8b67d17ffc783cb726ebec744a0ed62c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic1a3e7a14eff1a6da9e96ddbd750086b011cdc44e8aa1189879b056fc48b3a27;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iee4c52c7ebe29b796d3815def71a1869f8acb0bcdc109ad21b59ab2aa610c807;
reg [MAX_SUM_WDTH_LONG-1:0]                  I215ee2b19d3ea96eedc62d8cb097051dad2d917dfb2eb2b0e1ed0ff697955765;
reg [MAX_SUM_WDTH_LONG-1:0]                  I580713ee6afab29f13f6dbda18d77ae815138af729f981a455d34aca294bc4d3;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibbfd537ee459654bacd89b68f7d66565efcbdaa3838dc0847f83ba17c49b404b;
reg [MAX_SUM_WDTH_LONG-1:0]                  If18d826ce7582d4bf76e5968c9c86b08281682d30b790679e01e9aafa86f195c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iccf845c102c65fc97a1244cb2c0182925c72e95fb4a9b0dc97379f5a32837612;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iff4ecb0f057c396e2e94c919920695cc67ad53f6b463c28baefee01ee00e4942;
reg [MAX_SUM_WDTH_LONG-1:0]                  I32562e9f1cb6c7224d2efbd29f393e04c0d655e4bef402c2689cb946013f5d1f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb8d3dd7bb86ab8f1237c04d9d07d1d6046f07c618a3bd3308c59483260b7365;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8ee1c7843334dc659003797fc7ec177037e184855e8e80063c6e490425de9446;
reg [MAX_SUM_WDTH_LONG-1:0]                  I63450ac287a1e882703f7362bc499e7c779a7e68a1fbffd944aaf0e770fe18cb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5c6a9cfeb6a0354276fa86b65ea21b018e71d37b366f907012b41156aa22bfcb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1288c340fbff871d0fb4e5aab171e965bdf5b3b6cde30bb17f6a8d04ef546109;
reg [MAX_SUM_WDTH_LONG-1:0]                  I76041755b112a333460289875673d3f2b054918770d3a2cc46ab7a9f92b50eb5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I559a54fedbda0d961279ffb3fc4d2eb644cf2b77f805acdfde54df03ba0c05f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I30843beae9ebf34c0f73f773e1af0422e40b3ced201574b6f87f400cb37a7175;
reg [MAX_SUM_WDTH_LONG-1:0]                  I628a71f11553d99c7d0f19a7932ab7250a9448868d3e118479c70d70e1481ecb;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7f99ba04346760d4ee2589662be79b19673e741f07d1b9c0c35b54d4bcd3cfc0;
reg [MAX_SUM_WDTH_LONG-1:0]                  If06e126d9560577dd7525491f2092e8e9c9ff9e64c0ef94b3d0ca2b61cb6392c;
reg [MAX_SUM_WDTH_LONG-1:0]                  I311c88c2854536dbb8f578bdf98823eaf5888a7c772bc2c6f0cb49c9c9c79500;
reg [MAX_SUM_WDTH_LONG-1:0]                  I42760d09b067c76aa603d685d09ef8a3fb0aeeeef30a19648ab2cc69233d8514;
reg [MAX_SUM_WDTH_LONG-1:0]                  I073f480ce57215d8a9930ab34bbed6bcf5e631613fced0e782749a390615672c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iba06a153040bdb18311bb9c6826eddd28863470c44a75683bff1dbb5d03e1d39;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iaef86ab80a38f09821c64eb7b93cf066c0ba40a4b315075fd4652eb82b687bff;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifa64872cb59e066ea755fd8d50aa1fbdf10fbe3920e9ccbbad20c899f377207b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id523ce79d9f7a6b24c5979c58855211eb2bde238c81e549064c23ec62a5c7a3d;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc225eef673a329e451a89e36893eee8b9d8d9b8cfc911d6bf84a2ecafea5e4e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id27c2a1647e08c46fba102b41eceb3513a697df9876d76b23fc4118f16b479a0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3bbfc044ed936cf51599cd8977c7bf894621c83e1e73c4cea372dc54a1d6c028;
reg [MAX_SUM_WDTH_LONG-1:0]                  I54a09dd4115c1f70cff7fd7921120216494997fbc08a7e9eb8e59152ef12a9e6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I809ac54f05fda9abf4917b1e555505f9eb41cf89a9a9fa098fd642e90bb635b0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5a2063e62c2c96b172ecad9fa950c0b42c413214e30d94796ca9c2b8c6bbe522;
reg [MAX_SUM_WDTH_LONG-1:0]                  I3435109d555534fce5a4cccb9709c25bb5ea401158c144add8e4c09a6a68c8f6;
reg [MAX_SUM_WDTH_LONG-1:0]                  If0c2c0785586996991da246fc01722deded4e3ca8550290626324c5908d770a5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0fc48ba2f5bdf67aabf15071712eabd08121ca31614dbbfb3ce3eb7cf6287364;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icb2218fe2214af22ea6fff2b9ff3c8d1772fd9318efa83c7655b0dfee2f6ab4d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36a6b8814b16f2a3e44bf1afffac6416088645e41a495b7dcf9053020718e983;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0c567cd54c6fded476f507a4a35d7d93fdbd2cd1c555e10edf313ddaf4b0d64f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibbfffde74fd960499ea7e7ce9dbd03e057746dd164bc9af0e585839225056f42;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic49fb172f5523a522e94efd83b5827b8f63c2d8fd7c76263249d96a00a0e25ad;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0cfea5b22889a1b983f14e6d1c3bd847f20dd9cd96b0cafe80e1705be750eb96;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibef81155a593cc991eb8f0da7ea8dbc27f3c935dc1fdf7b857110407ef449718;
reg [MAX_SUM_WDTH_LONG-1:0]                  If34a395225bfb809ae5327b364a127aec5b1e5ef9e4fc9bad4baaa13cf13f661;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id1c35604f896316440f1deadc55ea39d16307edf0e2ddea1d7d450c41dbbc705;
reg [MAX_SUM_WDTH_LONG-1:0]                  I31edc2dea3cdd499a9a2035d2460448786e5a44b1d828d6486d7c3ccb959892b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic00c95647ac3595e199e62c4d3e75956755ac952e4cea464b27066ad8f09415f;
reg [MAX_SUM_WDTH_LONG-1:0]                  I31d6cdf7439ddccefec7a19dfdc442d351d609dca8f14aa276c22741a45aecee;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4d89a637472e8c4d071c44792883afdac1fe1c6ffa9d08f7259525884000b34e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I2b2cba74c6c9eeade51d69171bf22d1de38947948b7af485a5e64aa9bd90d71a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I081fd1385ec974da04b64bc5764efd6db252fefa40f518ed0ed4b01ce630064a;
reg [MAX_SUM_WDTH_LONG-1:0]                  I45a1490302e61b9172caa0feb0aea621e97a5a95b9e8c525d3ad875898955f02;
reg [MAX_SUM_WDTH_LONG-1:0]                  I57c394b657ecd32691fcef200ba361abaffca7d8ddbc7bea22502a9f7bff9f5f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie22f10e98c9847ef82cfedf9cf3ca17fc0307139848522f58fe0ab8f92d253c2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia14c31a81641330844c0c48e155c6f7630695ccf3e7238ad6eca01c8a45a104e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia40a2c6be098446003dc0b6caccdf75cd1ecce9fac58135f83551b0029ef7032;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iffdff1b757352d5f1174deb338f337fd8841ce8d132c2e0a16f18fc1a97313a2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifcdbddb54d9293f008a7bf068e7733c4ce75f38ee2cbe8ab4247bc4200a604ac;
reg [MAX_SUM_WDTH_LONG-1:0]                  If8c3dafd18d6fabac3e4ec4dce257aba397ab0d341e25a1bb88f9e32909deb17;
reg [MAX_SUM_WDTH_LONG-1:0]                  Icc54d76cca75160c97db719151bb55f2d112201e3812c72f002b3dba5e61575e;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie4b741e2c3f5dbd43bba89fbaeb4cc6b309042b53629f8db67121eb22a656ee9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Id2df947b4126f71a866a204090780296b99e4ca990d0d27c7e3750ffb4d11451;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib1a3877a6c9f5b87fd3c2104782a0699748b68ef73a12291b34e914344db9d25;
reg [MAX_SUM_WDTH_LONG-1:0]                  I8601156c6a18f07b4580760c232a62262c2eb8d656282d9710517b6bdb886459;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ieab221c067f0649e88f307dd8c46981653088853874e2a256b99f7b7a8bf93d5;
reg [MAX_SUM_WDTH_LONG-1:0]                  I19e014466929e7ddd8d4a2a3f0fc6cb3d9eec8d39e8f7a81458043ccaaa90ee9;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic80161feee5be9576086dd9d1ed8adca369a841f0052af01b2fe93d46af669b2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia24a2450394a5e7953feb8631095648c20bd71240699f481a0c3b748e665aa64;
reg [MAX_SUM_WDTH_LONG-1:0]                  Iac4628a0a7bdc975990c2664a736112cdb2bf1b1b30f89ae1e6827a44bdb4474;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5434f08cd24b915586080bec92103df0eb2a3d6d14ee496326046918db03b549;
reg [MAX_SUM_WDTH_LONG-1:0]                  I7da6920e7bb85e837e61b04ba09453237164470bf2eb7607af94194e05407bfe;
reg [MAX_SUM_WDTH_LONG-1:0]                  I536c65ee87da658790b4273c04e7acefaa2baef5da84d48a9a53686c9ad20195;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie3ca82b8d601f023d408833c7b5445539ebf8f17bb678e486fb3f650b2e01d9d;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5ec53ebfd7533177d3d5a1d97e18c9e5f90e4caad316088f62d8bd0ec6bc983a;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ifc8ba6aad04e3418146443a14c520552e32ac2f43fabe430ef0d640b4262337e;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1090417ca7c539e5bb1077d4b96824cac49fc6bd3253fb6d0348ec13edb97d2d;
reg [MAX_SUM_WDTH_LONG-1:0]                  If1aa1bf1d7206ef9c00f8c1aafd738c03603858f9757a3f671242af1b139cc64;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ida31fcf4f48fdc3b391ca3e4d2c7b1c3ff6ce6ee53c2dfbbe1bc863514845a19;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97205d95f7ff115112b2b1a7eb32bf70ff7c1e2fb431785547ed7f98d5fea0af;
reg [MAX_SUM_WDTH_LONG-1:0]                  I5b4f25d6b0cdd33c4b4f5f200eb9ca9d2ad68b01b48f7697100305c1456f35af;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia6232cf34275276641c494e4f4cbd7a8796f1f946733ed0fe15d9e11cd8c740f;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic98f738736b6b689361d5a77495e45e51874de01c86f1e7c10fe07e2c0f3ae82;
reg [MAX_SUM_WDTH_LONG-1:0]                  I24883a74ba0e0eaf8efff93301dd4d714667c28020ff65d73e4056b2d014e287;
reg [MAX_SUM_WDTH_LONG-1:0]                  I347c2eca1405d163956cbc4ba007b08ae0a0a751bee7ecde367e2336fa308e26;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibdd97caada239a1152f2155c8cb9e25402600931810f6bafe34159894246d962;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ie0fdeb73844872fe9e7af165cda8d1c865df24e572180803760f4959f8e73ef0;
reg [MAX_SUM_WDTH_LONG-1:0]                  I4ba3a78d1129b6b95ec4421b8dc75b90921b67ed09cc636c1fe08c778c9a4c87;
reg [MAX_SUM_WDTH_LONG-1:0]                  I69baa1c18df6858ab86b75bb25b5f980db3508a861fc7da408a38ed95c910b16;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ia8fe4e59fc4b364c711cdef5a6718ae33543de2e35744d9cda4cf33f340d7add;
reg [MAX_SUM_WDTH_LONG-1:0]                  I877a8619724696e16819de80d99f77e7ec18579f9e3cd99092f4ac0d358ab35c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ib0319b3fbdfab7c4df3ba7c1d710d7ca176cf8cd4223ea11fe12102cb5ac7f12;
reg [MAX_SUM_WDTH_LONG-1:0]                  I97f8ce585d26cb40e221f7f8bff17e80cd5565540b9108ef64628053a3d547fa;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ice9d3685b31919d1cfe76a96ac6e1738ef6c66e069de55830f61665cb5bc0ca2;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ibef17646fe9cd45fe72647539df79962a2f02d56819071f9e7740a099175decd;
reg [MAX_SUM_WDTH_LONG-1:0]                  I36a3a77efd095e4c91274958f1ed4b9fc929f2b6794e4b879b8275f3a01ae48c;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ic2f933f79277b6967efca4d861031734f157410c96568f6370436fa3c94443d9;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0643791cd1c7ee5c205da45ee4720229c6f7b61e98a7f642afc47506f6e10210;
reg [MAX_SUM_WDTH_LONG-1:0]                  I34e2e324da2cf6bd7804e6c3d9a2e8af1ca0799f9a15e7c9597f812ee6679831;
reg [MAX_SUM_WDTH_LONG-1:0]                  I485c81ca3402c9b70ad8a10b749c0ee5e81569d1a64231a5fb25e3af8cc4abba;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0784dbf1fd934c864e5c23e58e5636d5e4e72af359af2dc3cc1c11653a96d26b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Ief695bef8a02a4f5e89c14ac6b89f84678cc7d7a9d71bf2a5e3c1abd44d1cbb2;
reg [MAX_SUM_WDTH_LONG-1:0]                  I1e024678e8d8668a4b3744b819e48699d59c21dd2856723a6af255d20bd83297;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0ce015383446aeba50b7677c9060a1e18dab91eb8040a718fcb7e104a700c29b;
reg [MAX_SUM_WDTH_LONG-1:0]                  Idadca14723005bf0db40379151927d667247f30071db43f735c3395db88dd110;
reg [MAX_SUM_WDTH_LONG-1:0]                  I9f790cf09f0d8b1c047cd0df401052898d374d930d5ccd784d142c544d8b54b6;
reg [MAX_SUM_WDTH_LONG-1:0]                  I0f94b265dac20d93ad623db13d43a951cd09643250c48e9d8f58e163ebb406c9;

reg     [22-1:0]          Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626;
reg [MAX_SUM_WDTH_LONG-1:0]                I96fb06aca6108479f7e21e1835a091a9060c2925cc6320c8ed71a0a0092bdeab;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie000dee1e3953811fe9424588b71a7dbc88f41ec69afd16e17e8fabf141c31ec;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie873b138e19cd7f7e8afa8bd8f8c4610b65d0fcd647e76d880d25f6fe36c54ef;
reg [MAX_SUM_WDTH_LONG-1:0]                I8ab1772a3bc752331b0bf62069643cadb48bc13bbb06ad3eddc68ac603d73654;
reg [MAX_SUM_WDTH_LONG-1:0]                I4bce49360270b653e45b914c493ca8e5b74beb0b6b85838bb3b54f1f39389fe3;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibb4ff9ffdb2771ff640bf958798f8447a0dbcf15ed0ef9f82068826ec621de77;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia4691d32d9e84827a250e0b3d6ea8142c24c9df4ade01c19583e6cfca06cd990;
reg [MAX_SUM_WDTH_LONG-1:0]                I3a1380b85cc7f797ff92d02b7081d1ec3ba069aac74162ca059c399daa10690d;
reg [MAX_SUM_WDTH_LONG-1:0]                I14919dedf2b4d4caae8efa1726435d1946f48e1e9b1052133bebe8affeb3556d;
reg [MAX_SUM_WDTH_LONG-1:0]                I852a201bdaecd968b6f9c9b6bd64dc8035a17fb92ffc806a690781666354b069;
reg [MAX_SUM_WDTH_LONG-1:0]                I345c0aef41ee2863a96a076a78d92c7498f50ef90e82e75565df1d1f38a08161;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifb94a220081758ce91634fef64be084898a662f7c0e8cc9f86859bf3852b3efe;
reg [MAX_SUM_WDTH_LONG-1:0]                I5f1b294a0702ab37f94304ae67fe91abc04c397dd682d371126a7ceacf7c43ec;
reg [MAX_SUM_WDTH_LONG-1:0]                I81aa911c9f6f4bd88314aa3c5310efef6c40219ca93521bbea3c1afcea7bb48f;
reg [MAX_SUM_WDTH_LONG-1:0]                I97f674eaee005fc7a54ccb648f5a0a67cec041e895d62eacbcc9a37068b912a7;
reg [MAX_SUM_WDTH_LONG-1:0]                I7628fd0a5ee3ec547c1b4798a4d76de651807424cd18f0b3b8a3bea849e6fe0d;
reg [MAX_SUM_WDTH_LONG-1:0]                I1d8a992801d3f6a457848578ce286b496d4e2a69937344bdcbab4e8b1af1fe4e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia28f68b737aaaaa6b98aa5e9696b937e564754edef217740c414c16fe2e485b6;
reg [MAX_SUM_WDTH_LONG-1:0]                I099e314496f03784e5504a35292defa79dc063aa81e6aa8764802f7fe3a47114;
reg [MAX_SUM_WDTH_LONG-1:0]                Id4bcb557769f043a7275ab01d6d9794d4cbbd9309be38f58acc307a1e693f347;
reg [MAX_SUM_WDTH_LONG-1:0]                Id1bb830ea0f92a1c0ed0addc915fc85198e4744c4bf7369b4ee1f7131f5f8542;
reg [MAX_SUM_WDTH_LONG-1:0]                I31009872a3e84f78bbf1f12a7da708c45e3b708bd943b6f4561ad436164b12d8;
reg     [22-1:0]          I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56;
reg [MAX_SUM_WDTH_LONG-1:0]                Idd9957e5b52c4d33e24910559d8203415afdf467bbe1c9de950145282c7eacf0;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a09910e62aa0cf665f69be80c9ad61f2d31115012314b8188cf79fae365626c;
reg [MAX_SUM_WDTH_LONG-1:0]                I3d6f6b104bd2ffb35ea6782748bb777ec7eceae47ef2e1d18d37d1677d56cb80;
reg [MAX_SUM_WDTH_LONG-1:0]                Id5055b759fe480d476c4bf08c420a5dafe9e65cb03c6d6991c1d225af0a51d7b;
reg [MAX_SUM_WDTH_LONG-1:0]                I93e543ef3d58bc8bd48a279299dadae1d7f4528c3d09d7106b969e15565d3a15;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib6ff050679c6366efde7b9809fcf42051f107c18863bcea79d41b5fee0603e9c;
reg [MAX_SUM_WDTH_LONG-1:0]                Iba81256fd46cc69f1367fc6ed7b712d2695e099c52b476f9b39f0a13404dceaa;
reg [MAX_SUM_WDTH_LONG-1:0]                I608b794037b45c46a29ea01e378b63a1f267c4b489b0866fe2f6090936fa9d44;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic48347f5264e8e479996a8dba0171a108b602be1e1d24b2fcb43cd2bdb82f61d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib62b5b3c80d193b97bd6b5c0d5678e424026381949c3f24546d367df930cbcae;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia7900b5a01cfc1c4db79ca653f072956c13e2040cbd94cf07de2f1d969222fa8;
reg [MAX_SUM_WDTH_LONG-1:0]                I1aa136009f34c39a8dbc39b4444642cd09c9cd2f01bd6310287d4ddc9bedad85;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic195e053a186bcb0e653c0ddec75c57d1b3210c583162dd90978858c98fa53f2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic859d34db6baa83e73a8627c251c877e93f15653973d0634c42a8ffc9f628bae;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibeb23788ce301c724494a2852312b38344c27416a5604c0145fa330ccd1f290d;
reg [MAX_SUM_WDTH_LONG-1:0]                I5ccf8e87b0b8e8ce9bdf4b3329e4458a628f2568184f82b998ac62ea28bc0307;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaea7277e745e05f803325e0f19dbc5a54234878a9a3cb2cedcc013e3942e9cc0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic94e7c887d7f24b573b470820c36fe8a0fef750e2c46675f8867d78f2100f1f9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifa0b8243f5ab6adb88a70fc1245e3480ea3fb3f3af846fdefd0613ca91d7b122;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia00cd24df6e6b22b466e1492500f1948b3ba3d70bdca407d1c22b4dfaf374eb7;
reg [MAX_SUM_WDTH_LONG-1:0]                I8b41f817a4008df0994e2efa6b33eb847e82b031082f90a767467ffc03cfdb93;
reg [MAX_SUM_WDTH_LONG-1:0]                I8d91c857f2c8154bb09d456ff73ebdf81e3b7d9bd1c57c2e6b8c2de74e55cf48;
reg     [22-1:0]          I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135;
reg [MAX_SUM_WDTH_LONG-1:0]                Id0f930aa222bd91b8a7d5f80a38d84993a63fa1c6aca3d37ed259294e08869d8;
reg [MAX_SUM_WDTH_LONG-1:0]                I58598429d44ad951f91139a213d3b0bdacac6d71f1b9753886dfe1d39d0024ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I3cca3cf08c967f80e7e255a590bb9c442abc535cd529f7ff304f25d5519dab04;
reg [MAX_SUM_WDTH_LONG-1:0]                I42d1b7202048c81ca3a8bba0dbbce65501cb7a519fde37085c68d01db7edd635;
reg [MAX_SUM_WDTH_LONG-1:0]                I07bdf8f629cfc9c094023be167a717880dc3a42099b01bffb431036521cd6019;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifaa925832248fd0e2f5841096d9618c2fdaa3c63a3130b57f493782f96473088;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c22aed0ed8abb0cb8906a35a4d44cfd7cc68b2924e474680a2eb6cf7caf5582;
reg [MAX_SUM_WDTH_LONG-1:0]                I31ca3705bdc7e063c61023d93193b3ced40cf440afd817d0d730f6c8d37f8b92;
reg [MAX_SUM_WDTH_LONG-1:0]                I789461a909fa4abaf3840dfca4f63bfa63fdab389e149fddb7d8ae2b876dc912;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ff3298d93471156b56cfbbea17c8dc0405bfe8654e9f830bb33bc6c9a649b3e;
reg [MAX_SUM_WDTH_LONG-1:0]                I9eb30c75f8d71ade925633d7c8bc6b948ae519cdff33ddb885761bf72a8b0869;
reg [MAX_SUM_WDTH_LONG-1:0]                I5456c559bdce4d65af540e4c71c19e44227c62e5c129b7de968ac7f311dd76f4;
reg [MAX_SUM_WDTH_LONG-1:0]                I98e4b84e98742d38b206ac059ad123966ee63903c616b9c31b4ba9615edb9f40;
reg [MAX_SUM_WDTH_LONG-1:0]                I40d7eae63827c6efe2ac480c8eb9f8a8f77bbfa845caae02d137397c9da822a9;
reg [MAX_SUM_WDTH_LONG-1:0]                I30a9d5330fac5c3ec7b63cfab0edcef0eda61dddb23d2aabf733b9982c12b4ad;
reg [MAX_SUM_WDTH_LONG-1:0]                Icbdf29918b91006ffdc8b68c707840ee6bb9c27779dabd372e2033888743409f;
reg [MAX_SUM_WDTH_LONG-1:0]                I7f6b89a61d6313029102fc48e92a54ffdece30e9eac1191d840c488be69d8223;
reg [MAX_SUM_WDTH_LONG-1:0]                I9471414594b824d60836981bf4b9931c135520ad1ae7dea177e0bc591c2572c2;
reg [MAX_SUM_WDTH_LONG-1:0]                I0e9135a0817e96971dc8c4fe6eec717a563c44738f7e38d5bfb2f4dda8c77876;
reg [MAX_SUM_WDTH_LONG-1:0]                I0847713503570d7ab3efee12577ba27aa81869a22b14ec8a244fbd4665d566f4;
reg [MAX_SUM_WDTH_LONG-1:0]                I7b529f16d1499766369f75cde5a356cb12c06d21f42a10932edc6d54146735a0;
reg [MAX_SUM_WDTH_LONG-1:0]                I1b93b1b2c5f55e2267a4deb4f75ca91039d6893af8e082ea85b7a5e9354117e6;
reg     [22-1:0]          Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678;
reg [MAX_SUM_WDTH_LONG-1:0]                I7200758287b0c7ed92552ced989756e1d49b5418181b9e36421da7e2694ed3a2;
reg [MAX_SUM_WDTH_LONG-1:0]                I96e7a523360a0cc0f3abfea09a566658e5e9f3316c3c412f99fd6340d1b64235;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic4839247bb24d460ee6d963d31fc390e8d9d679cd73f058d94ec34a18ceb39c0;
reg [MAX_SUM_WDTH_LONG-1:0]                I23ef4f4232fa0d8813a25ddca38a2745fb660c05dbe9ddc2cc33c47d45b3fecf;
reg [MAX_SUM_WDTH_LONG-1:0]                Id5e78e4ed6db0562ed51d1da1f34242f54def8255088c3a1ccf0221ee8fa153f;
reg [MAX_SUM_WDTH_LONG-1:0]                I17cdc222663e370d6ef2539ad03c45a7949d9606583c17568a24c528a3e8c12f;
reg [MAX_SUM_WDTH_LONG-1:0]                I65e452247faa2c9d6b01dcbbebd5e8c31884c88e70dc8ec76d55aac7e77e2d46;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib0641eb8fe554f69ebb57e8e900f995c07bddadffd25c01781ba234b87af4a94;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee9c2c6a9b8e84402eb1e0de611c1cb8ae1e802226f2c07833bafaba74f1ac15;
reg [MAX_SUM_WDTH_LONG-1:0]                I443435c78145236b927711299e8bedd0d29a743e3784ac22f70b2284b6be11c1;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a86387a3136768ab52d320fae7fe63c7c74bb5541d18889faa263c71b2bfce6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0c4bcb29e2939b889fb7a5a7b62b49a3eeb3ee6f4555518c9059cb34dfebc7a;
reg [MAX_SUM_WDTH_LONG-1:0]                I3de9fbe37d08009f5fa66bf7c59debe7da836dc078e212968afdc608b100e3bd;
reg [MAX_SUM_WDTH_LONG-1:0]                I7c6d90cd79e1b85ce9a5452570cfeec8faf9ce3e6bc886f66495ec2a66fc8c7e;
reg [MAX_SUM_WDTH_LONG-1:0]                I57d80f41498f8d7b91410dc02e646a45a3f05d45e9b5871ae95d6432ecd2af56;
reg [MAX_SUM_WDTH_LONG-1:0]                Ief90cf0b0997823c3071eb46b636e384077579beae3d85d29e639a7719763396;
reg [MAX_SUM_WDTH_LONG-1:0]                I295d7aef060ca978805bdf65138e5bf134551eda9c396a22165a77a3091dfd28;
reg [MAX_SUM_WDTH_LONG-1:0]                I73a855a590363c762c34008e77f73f961950c0dd71b795acab3adf40c4540453;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie38c638da580ca7d25fc0754497163d0369f31a6cdb4bd26663a759b74efd588;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c635a0b11af3be4774428af79ff5cbe6a32ede6ad03ac197ecbb3ca2ba78f8f;
reg [MAX_SUM_WDTH_LONG-1:0]                I34a89a8aa68b1657dc7137437574877b170659ebdbcc93a772989e2b8b5be31f;
reg [MAX_SUM_WDTH_LONG-1:0]                I9f9d895211b42c2c9d491349dbe7aafbad775942920197105c34837dba6563a0;
reg     [23-1:0]          I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777;
reg [MAX_SUM_WDTH_LONG-1:0]                I11c6d693bd6c019722571e1aa6eea0507f351a89cfc6d16f8fc51997981aea81;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib53bac100fd49f57a5185ff4ad973dfe8eaef6de1937bb32d9246dae9459442b;
reg [MAX_SUM_WDTH_LONG-1:0]                I7ce5fe43a760b5a43815388233952e1bfe5d8b5a7c002f26ae2d462129aad434;
reg [MAX_SUM_WDTH_LONG-1:0]                I3a2c9aabb8b064f82bd6f6571bdebdd704abb7526f4977a7b98613f883fdc62a;
reg [MAX_SUM_WDTH_LONG-1:0]                I52f4d169be660862052b60924958cc9a0eb99b1454608fc48d47192452f8b390;
reg [MAX_SUM_WDTH_LONG-1:0]                Iade009d6c5b9e00f5459c53b0c254dda356081e6965366db7b7ac42a992e3ae7;
reg [MAX_SUM_WDTH_LONG-1:0]                I52dd625c97050874c15b1980a389843c4a7a890d73f6efb003c4324c029772aa;
reg [MAX_SUM_WDTH_LONG-1:0]                I11bf8ca77f64484279bd3f36febe1c6869fb79b4585a800449a0e5c683c6aa18;
reg [MAX_SUM_WDTH_LONG-1:0]                I255a6c7b69c31d60711a86b1f0da51040ab60c48952002406e028a200a835049;
reg [MAX_SUM_WDTH_LONG-1:0]                I24bc395a7644f2a2d7702656737c32662f8c2e8a7e2b2d4c1bca200dcdf49219;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia84166c5479fb08b9d5bafbf3446230d231e77cb1a3034b53477e2f0632ca74a;
reg [MAX_SUM_WDTH_LONG-1:0]                I544bba815490c8592dda0fd85cb612828256c09ba1431bc2632b74cc9cd2aa29;
reg [MAX_SUM_WDTH_LONG-1:0]                I7b8225b7ff4972426858a8550dc67a231d85fe94426bf0812906f1aee0e2d097;
reg [MAX_SUM_WDTH_LONG-1:0]                I3358739f5e55263208e661a339d6b29f188f07ef07e2ee7a63a24011a4f8568f;
reg [MAX_SUM_WDTH_LONG-1:0]                I5eff39d324b6a8910fad41786d651086c622d331987e649ba4b3baae11ca40ce;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a5c4f290852b8c1baa90ae00400045825f13c24b546dc4a7848f91824185f7c;
reg [MAX_SUM_WDTH_LONG-1:0]                I9af65d3592633577409561b2069e30c73196d1a4798cb92f4d2f14db8771895c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie2261f6d4e2c2ce04997cd365593486e02a7d85106b9c3b568ccdfcda7a9c352;
reg [MAX_SUM_WDTH_LONG-1:0]                Icf0b2747a9e17f2d2672f7a17111c6bf54bed7d8fedcb5260f25fdc4280ae727;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifb6bf654293ed3bacd2a4ffc883b8ca5e4dedea39e338bd1a30b21e8f8df2f62;
reg [MAX_SUM_WDTH_LONG-1:0]                I0f4ede6017039c42f04051822cfc539cbcacd77427efe92d393ade1c10a46462;
reg [MAX_SUM_WDTH_LONG-1:0]                I23e0423ae4012d108a4e6a495814e0e6f920fa6dcab900bb35cba7b95f590c9b;
reg [MAX_SUM_WDTH_LONG-1:0]                I571233769cc63838bcc3d61e7a5e95805c3f4116c0053dfe86831eafff7c32fe;
reg     [23-1:0]          Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2;
reg [MAX_SUM_WDTH_LONG-1:0]                I7fbf7b7f7a1f0155cb188ee4219620cb35a2fcf98d2687cddfa2508273b70154;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f56f225d6fa40e0469f803c2f72ca27e9c45768ad2af9af9ad10e529e249aa0;
reg [MAX_SUM_WDTH_LONG-1:0]                I634dc6f7c843c6e4c63ce6a21b9cd7a386600d1155c0696988403fc1ab790217;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieedfb1902d1f76f95f5f971b578c2440fa5de47dd78e9dc70c35698f813048cb;
reg [MAX_SUM_WDTH_LONG-1:0]                I88272c473a90efa576a83d0c277090f5814599e5aa192b878cde74215909c46b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia3e877a9f66cb7582b125e56b7c3f79601eb8e700f54e14f967a4d9df9b5725d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie278ca9a470ffe4ac78bc335aec472b66707cf02bd91256aff2e7c73b5d2c6b6;
reg [MAX_SUM_WDTH_LONG-1:0]                I5ef535b2e573d96fd518cbd837132928a2a0c6a25d4eb3c360f1cc0aed89656c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic486b9953b158eae95a2d8914f8144e669e056675946d245c8239bfc249a16ac;
reg [MAX_SUM_WDTH_LONG-1:0]                Id89c8a47964d1e4aa4bb9e96a79092cf7fb55eee5808d6323ecbdecf8926adcd;
reg [MAX_SUM_WDTH_LONG-1:0]                Id1e80f29821e7ae727d759f44b21e84843025c938468caf7c8adfba52f1cae43;
reg [MAX_SUM_WDTH_LONG-1:0]                I7530c712ec14c8fe97d1699177ef642847c5c1ce6185d1eab39b8416b562b454;
reg [MAX_SUM_WDTH_LONG-1:0]                I41b365f8c613bf86dc5e2ed41719ec6823046127babf87a083503ebcfd38ae75;
reg [MAX_SUM_WDTH_LONG-1:0]                If9bd4d7f3740f15bdf597de00eecf1cbf2e3b4efdbacbbad889c0946a6b34a24;
reg [MAX_SUM_WDTH_LONG-1:0]                I31c470f2adda0a23b85c3245646a168f2478bfdff11a434c1455be20db703c64;
reg [MAX_SUM_WDTH_LONG-1:0]                I9fa9c98579041b6735eb78f7b3727824dd61991c6a6d91a158c6ac65cb20b05d;
reg [MAX_SUM_WDTH_LONG-1:0]                I9fc6fbd6f2f888b9750fa59a966971aa6ba6fe4eee8c8f3ed4c3ea60141a7d23;
reg [MAX_SUM_WDTH_LONG-1:0]                I8c133563a8b5e359a6a45a7f3b4e939fc84766f9fa09634d18e5d2101d0c0645;
reg [MAX_SUM_WDTH_LONG-1:0]                I84238bd7e53e0dd7ba07efd813661c8cd1648b76c44665dfe51fd07dfaa9b249;
reg [MAX_SUM_WDTH_LONG-1:0]                I6c3a9695a1c1d22809b1378e82cbdbebc1ca78428194df50cce0a69d6a159398;
reg [MAX_SUM_WDTH_LONG-1:0]                I4d032ff7482be75de7d2b816ddb2bebfa9e896e45fdade2b5f81b35c003a59ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I6b4d2a32c92c22b1cfe81ee6620c69af1850621deea406d75f098da0542843e8;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0964979ac559942d1da1c41ecb3d9e94c6c7c0da3d16177cf2379db8f37aa65;
reg     [23-1:0]          I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129;
reg [MAX_SUM_WDTH_LONG-1:0]                I236cce67d0aea9f9c8d5ea3c39cb598d55f734b44ad6e3972e7f6b91d56001fe;
reg [MAX_SUM_WDTH_LONG-1:0]                Iceb8741c9680982b02ba9fa2dd76d3b45155ca5f688b70c41d66f3b3690dce42;
reg [MAX_SUM_WDTH_LONG-1:0]                Iac9f4a2fa823ae63e73b655020376580991cd4b2b3123204a757afeefe35a10f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifb57457918458a6aa9c5df68dbb83243fbc49b3b7037575f43749dfe1bef373a;
reg [MAX_SUM_WDTH_LONG-1:0]                I91589fd8a2ab91f079bb41631c44926b2c6f83b82448d758d97578c314d0b76c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic20b5a20229313d70c01a5f53e13e96095c1d8695144668e66efdc81efdd8374;
reg [MAX_SUM_WDTH_LONG-1:0]                I53e90d4a2bbfaffcf92f2e9fd80c491e61990aa575337df13d24211a558315a0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie57b3acbbf1d1593e02ad38bc0e07bb84db2655f9282adb3ac5edc311e882641;
reg [MAX_SUM_WDTH_LONG-1:0]                I632095e999af63661b01bfe8bad0078cfc2e74217253d3971230968c235bc526;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a66a98136fb7fe52fd830d869dc53a3855a545aedc1d16927f76bc12e319060;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifea15bb5031583fe42f92f554866179105e46b1eac3c6b691958a998c26ac2da;
reg [MAX_SUM_WDTH_LONG-1:0]                I8b2c2b27add863ad56639a306f803b656ee8f91170e649d29aedc5321181f857;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie3290070e785df28e64ff4df124d14c370c9edb924d5f35b059a6c82e8373f91;
reg [MAX_SUM_WDTH_LONG-1:0]                I02ed3128371185efeae1e27046aa378006ec78d7c458dcba137f69c29c4363bc;
reg [MAX_SUM_WDTH_LONG-1:0]                I8dcb7a5498da4a9d3e4a76923e84c88a30ec174503cd435864a066ff0ff464ba;
reg [MAX_SUM_WDTH_LONG-1:0]                I94024b61447a332a2c36a75bbf305f3fd80606bfbfcc4ee8c5783e3910e9840b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibcddbd4e851466c5ff49f13244c2478ab6c089e6d8ad294cdfbdc8451ac6a895;
reg [MAX_SUM_WDTH_LONG-1:0]                I50ff347e89fb452beb071f112e4a51e074cb3d66bd903552db23c17670286e7b;
reg [MAX_SUM_WDTH_LONG-1:0]                I8b5ee5d271abdbdc518ce02f900da21e858d3e2530585fd859690a1a71502434;
reg [MAX_SUM_WDTH_LONG-1:0]                I54e64fd01d9aff7ddfc4babeff6703891da38578bb141d250c4ef5949d818cfb;
reg [MAX_SUM_WDTH_LONG-1:0]                I448065f71638c5abddd1eba1fcf567566281d5b4b23ec4ff2d2208d32a506fbf;
reg [MAX_SUM_WDTH_LONG-1:0]                I6ed6ee11f6983e96e7ccc4e4be6ed8c4ed166ca9075b9cd218f26f018ad2140f;
reg [MAX_SUM_WDTH_LONG-1:0]                I0678dba3dc1a3400ab26e223257bf71c03f0e8d284810653b5e507fe964427f4;
reg     [23-1:0]          I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856;
reg [MAX_SUM_WDTH_LONG-1:0]                If34d8ceb2732716c923a7f250495970948ae431d5f1e0a025618c1070940ec39;
reg [MAX_SUM_WDTH_LONG-1:0]                I60014273d45dd5019a1b82bdc0a65e44d9a16368d996c8c9ff312fe27e236171;
reg [MAX_SUM_WDTH_LONG-1:0]                If16869134ec7e59b567e29a1125f0d27eff7a3c612240e25462e2ee84a7e0104;
reg [MAX_SUM_WDTH_LONG-1:0]                I8d95c0be0c84d3ee590f8e77065a6ef224e0a75b50aeadea980f9ef4b8d25001;
reg [MAX_SUM_WDTH_LONG-1:0]                I28940d6e8fc5937055f8f50c0d65ac9fd892bdc9f0f2a571808f930c8ad21717;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifbf3cda7e0639ad343a64c5b3d2f45017f1d280bf72c96520cbf272104c90ad9;
reg [MAX_SUM_WDTH_LONG-1:0]                I4aabce2cc01e829bb9c3d6a984cf2b5bf9230cf3913db788c47a932ddf71b869;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic9dc8459f6cd65f223a6386c82f754469ef74fbab59ded4fd1370fb69136c847;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib22de4dadb6e63ea49c52cd8bc86dadfd7b73a002dd8e726a9cf1b7b299a8c46;
reg [MAX_SUM_WDTH_LONG-1:0]                Id6c8c2ebab66fb903f108466c8d15060ed1328fe9a979858569c39069bf050c7;
reg [MAX_SUM_WDTH_LONG-1:0]                I385f4177f3a22b6fa4a6352d164c7d54c94b980806080c51d00a65f030966110;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibcf016cc83d0fcc2c731aa53147c199b32b3dc7a9f1a255e1a0e31615077205f;
reg [MAX_SUM_WDTH_LONG-1:0]                I7e7be31550be1cacb2acdb27d5120769dd7a0a49efb833051ceb83c8cf691e21;
reg [MAX_SUM_WDTH_LONG-1:0]                I26d08096b43367ba37b8f6dcd919bf4ecb9c660a39f2c0ae29f655e42b88887a;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c200a5ade27683d4afd55e06371f9880a7bb99259e2ccda5c368fe46bb385bd;
reg [MAX_SUM_WDTH_LONG-1:0]                I92d28f6c97dab90de260df37f619e0a9000db48e278327a5c5d1528a34bb6dd2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib053c04dd4e330e6784846706317bb6c8b12f9b36a57ee12807bff7de8ba7f0c;
reg [MAX_SUM_WDTH_LONG-1:0]                I0f71479f871309f1717e7a1a2372ebfff4623c315cc31914588df3896740a074;
reg [MAX_SUM_WDTH_LONG-1:0]                If49d6a59c1d539e369406ee4e8a2ebb30199f46c335584e62921f98fd811001d;
reg [MAX_SUM_WDTH_LONG-1:0]                I051f072f564eefd657cb4d59c1c851b56df2e70861d875f3b4c9b95e8945db08;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifc8302f040679d23faab1ed8387a8a3aec85aba86ba9a78d3ca903126266af4e;
reg [MAX_SUM_WDTH_LONG-1:0]                I2747ce9b7349ed89e3265df62bb0d0e612706d8c1b61e30a2878094662da8ff1;
reg [MAX_SUM_WDTH_LONG-1:0]                I3619e836fee4be75d6700a0e72e84df3a5a61003227363b8c4d348b8353075e0;
reg     [10-1:0]          I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f;
reg [MAX_SUM_WDTH_LONG-1:0]                Id658b37d70ac8e3a324133f475a77c7948231571aa66ea0dd11b6460fca011a3;
reg [MAX_SUM_WDTH_LONG-1:0]                I737ae96fe290087c8ae686b90b2ac94df2185f7ad8b4252a6ec850278ba5ea9d;
reg [MAX_SUM_WDTH_LONG-1:0]                I18777be7a1745485d18289e0b4a6e43e8a2e6758be0967b8cea04a3b0faf973f;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c30d2957a73fc51bb7044b869e28e0a8f6e0378a6098ee5e244efb43ab6a690;
reg [MAX_SUM_WDTH_LONG-1:0]                I69f7964c2f630ef03f49c2a6cac12420e0998397470245e6afaed2546b33775c;
reg [MAX_SUM_WDTH_LONG-1:0]                I6f63c71eab6c2d7e3eb41fd78c9e18d6362d2dd4100c72b43d3e4b9d06663165;
reg [MAX_SUM_WDTH_LONG-1:0]                I23c91b29deaa2df1f4d96e343f6fb852a2b594937a4f62dc4be1fcbe0347c439;
reg [MAX_SUM_WDTH_LONG-1:0]                I8411087f9f6fa41d454a74dc89e5152e5e8edfa501c8753bd0735cec3789f14b;
reg [MAX_SUM_WDTH_LONG-1:0]                I119a98150511650722429eab31b5785e99128641bad59a3cb31e42158a648c48;
reg [MAX_SUM_WDTH_LONG-1:0]                I28a2b1ada19dc69ebe4949a75633b2f543159d2d1cc169f3bb6070c1419878e0;
reg     [10-1:0]          Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibbbf3f4aa7f74c37a0e8ac8a675ac9a9fec748ac720e6a78e9cf937dd089b8e3;
reg [MAX_SUM_WDTH_LONG-1:0]                I59a4b1b33d114a1b5bdd708e1f856f4bf729c6b86a4064967ca1faf779189164;
reg [MAX_SUM_WDTH_LONG-1:0]                I9b13cfb3566db96edc7c018b88f158faa57e4db029e3982290989c6fc08163b2;
reg [MAX_SUM_WDTH_LONG-1:0]                I8a1ba53134dcd1141a6f03dbed0f18ff7be9728dd9a6d6b138ff266c5307ba24;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifd2ca31ff3eec501f34892055a36979681d27574ed8007e4df5cc0109b71bd89;
reg [MAX_SUM_WDTH_LONG-1:0]                I6b2620e847ea73b8618ac7bdcd8236c4278de3bef0bf1511ee9779306438fa38;
reg [MAX_SUM_WDTH_LONG-1:0]                Id2cf59876d070e0f34ee834d2691f7fbdb039bc9273329e2ce8eddfe736f0a45;
reg [MAX_SUM_WDTH_LONG-1:0]                Iae213c2ac7729f8efe23deca256bf56f030403ef6ac00a3bc181414b6a3aa75e;
reg [MAX_SUM_WDTH_LONG-1:0]                I08e50de7e2aae48cc03a9959d08cab30d3c1c2ba8c4ef0799645787b0c09473c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibf22dd3f14f19c3fc769966f72e8ec980dc79c2991f69d03ca2defb7f720f880;
reg     [10-1:0]          I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibdd37577b403da9aa72ec3f4707379b1151c0b15edbfc4fd304c4e35c1672da6;
reg [MAX_SUM_WDTH_LONG-1:0]                I8e23f89e84e219d5351bdfd4aab58f61c1cb310cc731164c6e0dd2eac37b07af;
reg [MAX_SUM_WDTH_LONG-1:0]                I3baaba73f51f47e6a3f2310f692de9f7b9a871c65605e14d204d6965153ff4f0;
reg [MAX_SUM_WDTH_LONG-1:0]                I82d316ed1475017844ea73f32085b755d17c9fdafd8191df2e363496e1950869;
reg [MAX_SUM_WDTH_LONG-1:0]                Id9e3ea08b52843b4a9426b735967bd4ac3d49bd67ab8fc85688b0f55e6df186a;
reg [MAX_SUM_WDTH_LONG-1:0]                I77e34c24ea46e99b6bfc0f960d428d6ba3ea4f9261d5a183d83c386f259ab431;
reg [MAX_SUM_WDTH_LONG-1:0]                I930ad334ce972f0b5dbddf698f6101a196d8072e90d8144b31ce3f4b48a73e59;
reg [MAX_SUM_WDTH_LONG-1:0]                I4c0096e7bbf30db97520f824e05dbc28e6d1db344202349993fc68cbc95d6585;
reg [MAX_SUM_WDTH_LONG-1:0]                I75c796f56576dfba821e867b0de1a871ef35851371c3aa422532bd287f02ee11;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieee1d2436dbda6f58f19df70b691a4ff28d37db8ccc12e04413e45f80d7124e0;
reg     [10-1:0]          I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d;
reg [MAX_SUM_WDTH_LONG-1:0]                I65b0824920910c82c7d677c2dcf4216e86940b3edc0b3da85d8f65505f58ad48;
reg [MAX_SUM_WDTH_LONG-1:0]                I169d92aaa7eb4f8516e38745955b91d8f6e0ff43cb212186293bb78884282978;
reg [MAX_SUM_WDTH_LONG-1:0]                I492e47d35231729b266a9f31aba61a3ac2c93a9786a20f6a152d342cd1d0b911;
reg [MAX_SUM_WDTH_LONG-1:0]                I2624a2d841eeb09774127e5d709364f803826266b46f0fc3122fcdcf0aa129e6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6414b3aff6031e10856953f6b15ffdb0971aeb680d784a7199386be15624ff6;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf94ae58c1d9c9206d02651cd03cf2e02bba505f76b849158530a38382396ffa;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0a40c2a77389cda4a8333aeaecf37a2595fbda87854a43162ad1299544bd9e6;
reg [MAX_SUM_WDTH_LONG-1:0]                If692b993dc571ec401ce86f38a18ea4f96a797b00c04699ce83ce875b7c31730;
reg [MAX_SUM_WDTH_LONG-1:0]                Id5a74d0be90678a7b69691c10e4ab75b47914e213e67eae2f20d4b58e8a8d9ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I47b54f01ac82a9eb80a681633a06c4e1d432d358091e9d079f74484f40ab3e09;
reg     [5-1:0]          I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34;
reg [MAX_SUM_WDTH_LONG-1:0]                I6201d3c2d85bffa03f368b5862fba1b2e0ce3735fcc8711cb8107adf16ccdeb9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifcc25cd8dc442c6720ac0f764b432530aa63681953d8ba16b441892ff5966bfa;
reg [MAX_SUM_WDTH_LONG-1:0]                I256cb35fd6d4e6c6e1c1a9b42dcbc307f858e5f9525acee9fa7af42c820664f2;
reg [MAX_SUM_WDTH_LONG-1:0]                I67183da8c2763243a285b7cd41d838337f98eb6e59feaaa0a9150bcd6c29877b;
reg [MAX_SUM_WDTH_LONG-1:0]                I730fa6d01ade8f1439b29b955c5cff62700a90e523a4f4208ca2f9978e59afcd;
reg     [5-1:0]          Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d;
reg [MAX_SUM_WDTH_LONG-1:0]                I37084afdf6695d3b8fb0530643c8b03deb2499f4f68ead04e3b5b79aa4467f73;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee510842ece3717ba6eefc3ccd844e97a9718788683d4c7ceaefa6ca0030585b;
reg [MAX_SUM_WDTH_LONG-1:0]                I53d3de58d6308b770e4a8884447a5f0b92931c8d83c62c86714b6e539b498894;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e8142c7ece070c02ed90211fbeb423bc2a4ab19fae011793be99c68ff103705;
reg [MAX_SUM_WDTH_LONG-1:0]                I425913b12fc3c865d95f1caead00d8c49de08765b634aa444243f4a03a53d0df;
reg     [5-1:0]          Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibe0fac26b5e106fc1753aeb842e8a04067fc91c95e358b1caa58db8192381837;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibadfd4f0852067e83ba6f0d57699585ae20eb542d1ad8f2cce3bda0d043ff2e0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ife27bd449bf6acad3f06d6e337bfc29c612ba6b3f06927e6f9699ab24d1e836e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie130bec82505842b184f5dd86865ab095110bc65e59662767e152f427dd7462c;
reg [MAX_SUM_WDTH_LONG-1:0]                I2abc1178fa35959d8eb41342a7d7289e29054439c7bc06adc61f3a1d2e55bd6f;
reg     [5-1:0]          I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a;
reg [MAX_SUM_WDTH_LONG-1:0]                Id27dfca888552262f492b81fd23b881938f66eb15f7ab21afb210fc6056fa09f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia96c921ce4e0590c903d02dc69790c6af52898da90f4766121fa7b31e0ce6190;
reg [MAX_SUM_WDTH_LONG-1:0]                Idf239af48228dc01198fdd7240b8282cf247cbc6969403dd994aeac0e5f81898;
reg [MAX_SUM_WDTH_LONG-1:0]                I6687de5f8cb258492154a67fd3a3d5ee88d97a4db1c6c273ad158d5205ae3b48;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib924c4eaf872874debc3b6ee65921f0381331e1421cbfc3bd17e8caf273049cb;
reg     [5-1:0]          Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379;
reg [MAX_SUM_WDTH_LONG-1:0]                If53d34fa90e564a24f6e116baa8a7934ec4c51c5f0bce8160f0f389391792fe9;
reg [MAX_SUM_WDTH_LONG-1:0]                If0fe01f34db565bf669e2df82579abb4d3629e8bb001bbf874b9b76f8f780a37;
reg [MAX_SUM_WDTH_LONG-1:0]                I61f7e06790f5516eba113bb79388fb515faa1b3a3bf06598a07f534ce2845618;
reg [MAX_SUM_WDTH_LONG-1:0]                Id6b81456b5d3050b4e1fe80ccc8f992cf56eb0f08a1d29ec1e7cabe1baeb0872;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaa0b6d0f2fe24db548975f410ac5b79f687b7646169247f3891ce9e4644ee0fa;
reg     [5-1:0]          Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5;
reg [MAX_SUM_WDTH_LONG-1:0]                I45ade5cafdcd254cc640ea8725da6961717fd6c50f747242aab6976ace4e8f10;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie2e727d2073eda2be7642a6a2937cd3c4e553d8bb6ec56d914231b5bfb12405b;
reg [MAX_SUM_WDTH_LONG-1:0]                I1aadd9b378df1ab58a1b1af097539d1407636833d9c2d8b08c8f70be326fe199;
reg [MAX_SUM_WDTH_LONG-1:0]                If83264f9ff9f7b77429559aff8b14fce54040210c6ba3476b77824c28b95bea9;
reg [MAX_SUM_WDTH_LONG-1:0]                I1cf0e3016bbd2d8e5debffedb198273a2d019ce75f2f8352a285d17264d262f0;
reg     [5-1:0]          I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729;
reg [MAX_SUM_WDTH_LONG-1:0]                If9628510f239b2275efec7ce187b8eb7360beb042a425934ac81632815361368;
reg [MAX_SUM_WDTH_LONG-1:0]                I7d0cbdb63988e88f9f3f69b35029cb2078b97b6cc9008644b2721eda7fb6cfad;
reg [MAX_SUM_WDTH_LONG-1:0]                Iea2bd90043dd35ae24830a90ed10d12869de66637ab0237a1ad459fa916b57af;
reg [MAX_SUM_WDTH_LONG-1:0]                I0f54db0f4bdec3ff62a8f1b5f4974982e3600a906dcfc79789fb9fac058c353c;
reg [MAX_SUM_WDTH_LONG-1:0]                I9a4f77c8ba9a40c1b543070a42451ed37c0f22850a4734cdda393e69c7b54733;
reg     [5-1:0]          I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063;
reg [MAX_SUM_WDTH_LONG-1:0]                Icdea1f407aaefacb918babc28247d540a8a52d513d26d7fbb5e81a41797e7555;
reg [MAX_SUM_WDTH_LONG-1:0]                I83ec3e2a8ec621acd2afe475255e144f2158e1941ec685a346b75fc471b9cb76;
reg [MAX_SUM_WDTH_LONG-1:0]                I25600d0eb62c066eda0baba4269851387918088406d117377eb8bcc2e080e426;
reg [MAX_SUM_WDTH_LONG-1:0]                If45b8fca9a85788040c10a47569139b44384357512af96ee7bd8cd98d88f8f0f;
reg [MAX_SUM_WDTH_LONG-1:0]                I926233df0c5e8461173cedabbf49fead4b0ab577d82f2585af3a1fb6e3130e21;
reg     [14-1:0]          I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15;
reg [MAX_SUM_WDTH_LONG-1:0]                I979c6bc2b8486315e3db6888ef068b88396857d05a62470d4f3c33833cfde130;
reg [MAX_SUM_WDTH_LONG-1:0]                If2b1e365b8ee6d4afa8536f5c2f5c80d31e86ab6729b26795614d75a6a18ef42;
reg [MAX_SUM_WDTH_LONG-1:0]                I50e7a3df23a8147b9a87cb5e38d44bce7613b2a717d1e3a8bda1171f9522997f;
reg [MAX_SUM_WDTH_LONG-1:0]                I3d6bb14416567aa7b8883b3d1778b55c251a22ed42b09bb3cbae6a5210cf11f0;
reg [MAX_SUM_WDTH_LONG-1:0]                I54b0a17c9919d856bb3ed7cbbd8e42fd4ffa33ce8c32d45e4be1e28b71426ee5;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a6a17ada186c2bb60e521443c0a5a0248d03242c4ae01b751fcce4abe853065;
reg [MAX_SUM_WDTH_LONG-1:0]                I33d759e40b55a0d83119f5c19cf87e6e3181c7e3eed94eec60fb52f9c376addd;
reg [MAX_SUM_WDTH_LONG-1:0]                I84920b6036437109dbc48865b69f249d82da5c7288a7eb7744ea7ea567e03657;
reg [MAX_SUM_WDTH_LONG-1:0]                I78f0dcc6533ef218ce6959768639c983d2119dd518e988eb3dcd6f0b4de98c82;
reg [MAX_SUM_WDTH_LONG-1:0]                If64a23ad02d1da21fe63cb33f95d37c576739eb181b0fe50d7a5101817b4ede9;
reg [MAX_SUM_WDTH_LONG-1:0]                Id4cd4fdc9fdb1198c2894543e212f665c925298f1c92b4da9c432eca9442963d;
reg [MAX_SUM_WDTH_LONG-1:0]                I2e15c5739b990462c8a17b590fb7d60ac9c7e6648b79e75697139f55221fbcc5;
reg [MAX_SUM_WDTH_LONG-1:0]                I294ca1e2c287bbe18783f7043149078d4fcc1c59e24792d75655fb29a36e33d4;
reg [MAX_SUM_WDTH_LONG-1:0]                Ideae854591637828f033505e4fc9dee34d82369d02f7680ef6887c597ac1ac82;
reg     [14-1:0]          Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f;
reg [MAX_SUM_WDTH_LONG-1:0]                I597d0e1b64b5d47502804c7ba47fd0c17322bfdbd4d332b11f9742713f76855f;
reg [MAX_SUM_WDTH_LONG-1:0]                Icad68e9babee274d9a5b79cf432d9e2a1938e06f51aeb564af6936972b3f8e54;
reg [MAX_SUM_WDTH_LONG-1:0]                I15b5266ec781a5ae11540d23bf8b1a0b2eb45d94ab6f367a872885ff3207d5a9;
reg [MAX_SUM_WDTH_LONG-1:0]                I5c1a09aa19ef4bb254881dd92543acf840270aa36ad4e0f5f63a6182a4c93a1d;
reg [MAX_SUM_WDTH_LONG-1:0]                I9afcfde9391d485e865b08f9b8ff69cc2ecaace5f5e26e27b7e1775b625722c0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibe932d914d189b275138de8d6f3ffb914940d4b2bbecb574fba3c6aed885c44e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie2abebb2c2604e435cea102275e0726254ad91df1973aece477e1e5315f82d0b;
reg [MAX_SUM_WDTH_LONG-1:0]                I8befad7180232073f2f7db5a3f546a5a1af79b21cc9cb00a13e266db4eebba48;
reg [MAX_SUM_WDTH_LONG-1:0]                I3a9293b8f323c7e097a099fa6beb33ca299723796aec9396365d43334eb55e35;
reg [MAX_SUM_WDTH_LONG-1:0]                I52698fa0d5291f0dc20fb5f24c33e968ea63f47765bb7d231720330b624b2fae;
reg [MAX_SUM_WDTH_LONG-1:0]                Id8d0e36ce1faa76feb8cbe0331f2179ddfc066b70e93e990b5d5bce17f505440;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaef8ec1714d2faf3d3b947db31b7975161077ca31fee04842efc1f7159104d30;
reg [MAX_SUM_WDTH_LONG-1:0]                Id8da43222903044cc48243a7bcce7864e66d151673396879258ee4af7008a706;
reg [MAX_SUM_WDTH_LONG-1:0]                I8eb86c8d64d83d4ac46667af42b6383e4d165459475ec6be9d547a70ef0248af;
reg     [14-1:0]          Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaf205cfa67ea9b2c39d6705da465f081eb75c326c1d80e63e1331a098ca9a4ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I16ffb13aa3dfd9da5da39d9b2246d5ab46fd0fdb7c02781abf4d8bd754bbbdf3;
reg [MAX_SUM_WDTH_LONG-1:0]                I9a15ed1b2fa413056071c97b4f003717902f38d29805752222c45cbb2cf58109;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a10084ceb62d383dbc5871a208fc087b23de418b2c780813ae950bf4e594c96;
reg [MAX_SUM_WDTH_LONG-1:0]                I63f5ecb10fc3ed9bd8bf79403afed8ab1a70600ceb1e755de0d44af98495ea88;
reg [MAX_SUM_WDTH_LONG-1:0]                I377aa224e1817d2ab5cb02a5a290a723621782607fcd59b319d8cec1b092bc1b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib1310cd21337a1faa061ffd12a2670171f582e03471ab315b90de9f8fc30959a;
reg [MAX_SUM_WDTH_LONG-1:0]                Iabc9fc6e9581216af19559d8e709ea0842cba4f29f3fdfb05bd71d6d9f7594ae;
reg [MAX_SUM_WDTH_LONG-1:0]                Id165331f616d7e8f347cbe46daff955009fef6f8c0310c64c01dd35990231279;
reg [MAX_SUM_WDTH_LONG-1:0]                If17c7df712b5dd40132ac60628bd514bc70092122a0cb89ba7d4559439779fc9;
reg [MAX_SUM_WDTH_LONG-1:0]                I9d7506b5ed3de0e32e821ce6ddd1c28aed177910ccacc4d4aa2a8ee57212d162;
reg [MAX_SUM_WDTH_LONG-1:0]                I734136c95a40c62745d684fc7e8cd1114b883c6209df11cfe01b9174cffc720a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibae97ff31fce14dd0506fdfe7407fd6260f7cf8584a01da77312b1aa48594be0;
reg [MAX_SUM_WDTH_LONG-1:0]                Iea011619fa5b0fb7d22dc4bb4ce3fcc4856dfc7286ff393fb329ac0d7e348207;
reg     [14-1:0]          I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4;
reg [MAX_SUM_WDTH_LONG-1:0]                I954e0367a6f3af96a7e033da51e7256543d7eabd37191d4b03f3077567cb629f;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e6d7d9769dc32e1e014951538f1cd1014e9d07b675e6369e88ad5a6fd400787;
reg [MAX_SUM_WDTH_LONG-1:0]                Iac4172f940fcbc93db2047b26fece588f3fa63ef255ef404beb5e6ea016b2ba3;
reg [MAX_SUM_WDTH_LONG-1:0]                I0e9a7c6c53b89ca2685615c270e8ef3d3f51fad8619953972e1037edfe633834;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib99b447a19aa10415461faaa8d8026b0073582bd078930f2cdf0f531259d9c50;
reg [MAX_SUM_WDTH_LONG-1:0]                Icd30277c9d839d833f27f571231dd138497796d3e7818460d836a48b87e34d03;
reg [MAX_SUM_WDTH_LONG-1:0]                I2862bdd9be64c24d98e80e8b662a7c97c70943bab3d49cc8d39443abcd5c2c3c;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f73c51d25db7485bf4a0d63f95f14fc0661431870ce704f70cbb787eb336f09;
reg [MAX_SUM_WDTH_LONG-1:0]                I2647390c3800518f2251794a7ee4aa2d71ca9589534cf73eda0accbd2b3342da;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie05c1da46b594d3c94aac179f6c98334d0d667cea08108719b44541b7b0a2049;
reg [MAX_SUM_WDTH_LONG-1:0]                I1bfa3da571b0e3d943ec7b9a8c641283e080bcc6502fa8317ced3c0a6eb2c4cf;
reg [MAX_SUM_WDTH_LONG-1:0]                Idfa7c6c8248be1a2f8a95c6c74a71be3126e039a31f4e16e0b964476c6d47953;
reg [MAX_SUM_WDTH_LONG-1:0]                I5c43417b1bd96dfedeb36f6d3405fc7f6b73c11a55f21ebe6ffd675e991a13c3;
reg [MAX_SUM_WDTH_LONG-1:0]                I71f31c9a9943d9fd422d00aa01888aac32dd8b34236bdd9bdf3e660413a3512a;
reg     [7-1:0]          I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857;
reg [MAX_SUM_WDTH_LONG-1:0]                Icc43ea934f0c07465170977b52d2f402fe155ef77f3ca27119fa665a1d918694;
reg [MAX_SUM_WDTH_LONG-1:0]                I78abc91706fec0893eee10a69916f7247b718169155038bdc0bb6f8661ed1c3a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia428f915c49f84567006696ba3f5c783035325755b4fefcf74d65aaae1f3d3c9;
reg [MAX_SUM_WDTH_LONG-1:0]                If270910122bcee1c18cc592dba9b38c026f792d8d1472400a09edee9d7633e22;
reg [MAX_SUM_WDTH_LONG-1:0]                I1517acf28729695d689aced1c7eb358d9acfc4453fedf95a76fc22c972550c63;
reg [MAX_SUM_WDTH_LONG-1:0]                I8ca8dfb7a3a8ecb9eac34d1d1ef4768d31b86a757cb7b9ce61ef159816ceea7f;
reg [MAX_SUM_WDTH_LONG-1:0]                I2cb1ae23e53b89ca0fd3d1df98b32d5b9e478e9eb579b0875981a6b056e8ef4e;
reg     [7-1:0]          I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca;
reg [MAX_SUM_WDTH_LONG-1:0]                I1a2646b8251f83855c3fe8f6172f36500201ce43b9b5ba2cf0f25fd5d540e89c;
reg [MAX_SUM_WDTH_LONG-1:0]                I1d9a8ff2514f112838c7e4f568303dfcac3f86d94003ec4f1a40a35b79ee8ef6;
reg [MAX_SUM_WDTH_LONG-1:0]                I83c8ad082be8fe1a71adac4f41a3bd7019d2df299d19f8e5a293367e49b04fa5;
reg [MAX_SUM_WDTH_LONG-1:0]                Idc29625b375c44e890e371217aaa25d5fda337ba8177fcceca881adc72292a3b;
reg [MAX_SUM_WDTH_LONG-1:0]                I6e88f83ef5bc5f950a4bcb904ffede2603201e72e362aedb8db04412f7bc2bd5;
reg [MAX_SUM_WDTH_LONG-1:0]                I7ff25e517e328eda581e7637a2114a7cffe873df520114410c0487e503c01aa6;
reg [MAX_SUM_WDTH_LONG-1:0]                I463662fa980f8a5e4be086aa5f37db53b1d6ea8dfe11725b8c407f779a168998;
reg     [7-1:0]          I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c;
reg [MAX_SUM_WDTH_LONG-1:0]                I8db02445666e4aa12d7e495ba28ca0eae6ef411094d30330e91eb9eb03b38aa7;
reg [MAX_SUM_WDTH_LONG-1:0]                I8c971b4c1be575fe328c0a4a9ecc5dc75f08d36f65aa58642976d971a6c316d7;
reg [MAX_SUM_WDTH_LONG-1:0]                I09e6d011dacfba2800f9ade6a495076a67e4acc6a944fd649a7c382422e8fa6a;
reg [MAX_SUM_WDTH_LONG-1:0]                I76599c709cdbb3f3cfe4071b96fb7dcdf8e072fe85ad5c8e7bbabd4f6182303a;
reg [MAX_SUM_WDTH_LONG-1:0]                I0d9bc57dbbebd429ee5a5e5dabc1cd0bd9f4de95a920346b9e61cee83969ba0f;
reg [MAX_SUM_WDTH_LONG-1:0]                I91716015389a9d3b1d0cc77327f439e02e54be0d3524b2cdbeed886eea673b10;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibc3e77c4d6cb28599b7a21c7992802beffb168f54d8dfa650750ffdc6730df29;
reg     [7-1:0]          I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562;
reg [MAX_SUM_WDTH_LONG-1:0]                I34f861f0a748b0ad1550db8ce40149dc638194b0089cf22e2380a39a49f8c902;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibadbb4e272ab1105914763e2790898c8e37a553a1b6726e8818431bf5209b369;
reg [MAX_SUM_WDTH_LONG-1:0]                I308f551a8479d066b2a4b473206e8f407082cf83b37a376e6b0e1454f7ea2635;
reg [MAX_SUM_WDTH_LONG-1:0]                I58c6fbcd5f77398c3514e6a850bb69d9f57880a387f10132aa63079c0a1f4857;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia9d25b6cb880b9a00c9bb27bdb80c08988eee46afccbd578659eb98301fbb8a8;
reg [MAX_SUM_WDTH_LONG-1:0]                Ied710d5ba03554d4103468029a9d895c25c10765b6e3d73bbdebc54d7cc7d8db;
reg [MAX_SUM_WDTH_LONG-1:0]                Id7dcf87d2a40e82e7f01327d834d5207ae5873a7e5133c3dddead9d0cb9703f9;
reg     [13-1:0]          I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960;
reg [MAX_SUM_WDTH_LONG-1:0]                I982c94b61dff8249f2f3055f60da6e2c2b0b56c403f151168b28a5a211aa6428;
reg [MAX_SUM_WDTH_LONG-1:0]                I710a57e6c5c8e228325430ba2a5fc32ed9da101d76ccf1d8c9f3397859b39ef3;
reg [MAX_SUM_WDTH_LONG-1:0]                I2cb87b14b006ce6a36ee5439eb18a4287c5b9ae79748faee259c0435d0dac81c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ife00518e7b24a5de694b56a32211898b3c23d2dbd2df91a4197216c23fb5aa7b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ica9ef16b19711ccdfe32e34eed347b590635f1ba7983272eb02f980f80642254;
reg [MAX_SUM_WDTH_LONG-1:0]                I9331a9d6610ae5cb77aa3d477fce0c0ad7378a884c86c4872a1573f2d8a90d8c;
reg [MAX_SUM_WDTH_LONG-1:0]                I48d9ec419ebe83e2a5a8281e7beac36acc9e554b86b154736dc51ff940f5348d;
reg [MAX_SUM_WDTH_LONG-1:0]                Iab97067540ba8c9551711cdbff0c6aa3993534d3e8b352bda090a0997c681afa;
reg [MAX_SUM_WDTH_LONG-1:0]                I25c667a6616c9a94f6618166c99298b28d897f9ac8276bb85816e4b42582cdfe;
reg [MAX_SUM_WDTH_LONG-1:0]                I2d2137ac29a7c23160dedc43e9caf010f72f7d08b057e49fcac89984e616fa5a;
reg [MAX_SUM_WDTH_LONG-1:0]                I11775c069ab4acd951a3ca47bfa65c7632a6a8a369bb103d0bb719806dfe0c57;
reg [MAX_SUM_WDTH_LONG-1:0]                I6e418efd4b385b2a298c1c53d344e35f593e8380d1c27d7cb62cfe35223121c8;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifd66abca1532f04fc777617d91cd2d5f4d4fee35c3f075e91639a196780168d8;
reg     [13-1:0]          I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af;
reg [MAX_SUM_WDTH_LONG-1:0]                I6dcc482b16866339b78b922f9a7ec0f4a0ef311c353e6a4e107dfcc351abbb23;
reg [MAX_SUM_WDTH_LONG-1:0]                I8c8bc477ddc4000dde6459d7cbc4ba665fd4ecd97242d9f9fe97ca6825bb033b;
reg [MAX_SUM_WDTH_LONG-1:0]                I54da11ab334a3942047eb5953935aedd00ef1a24bb5361fba51504632ae61831;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide2ca364c5742f786e5408980fbe12322ebcc2920fd99ed322112d3623d9e372;
reg [MAX_SUM_WDTH_LONG-1:0]                I6024b75d70e3da7df4e532e712df56a8bed06352ba0a545ec355f59473929d41;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia79355adc994f77e150b93a3e38c8bd6f0a5848a212ac64559cf1210ee0d11d7;
reg [MAX_SUM_WDTH_LONG-1:0]                I1b68e82cfc8606d3a9325ff2da047f345e2f34b44eb428bf2a3bdcf42a6e869e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia1d4bd5d90332afbfaaac3cd0d8f5fcbc626ec4adbb0b0f16fc80923925f703f;
reg [MAX_SUM_WDTH_LONG-1:0]                I87af49f5f04df14686aef62aa27c16723af3ad05398f00e29788666b27784de5;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic1211f3a0703e281ce073a20afbabe9b2a698d1cf74f07f099d21fd89ffc8908;
reg [MAX_SUM_WDTH_LONG-1:0]                I2985f4f17b726f40ab6609b57a796727fe46605944c5e25c594caa8dfbea9f58;
reg [MAX_SUM_WDTH_LONG-1:0]                I6f7aa66db409365eac05a200d0a0f1d2b25e9c37ba4a7db3b58a7298af0fd6e6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib1e319af12dcd98c09841e8b06e7af86f2569bd7afeb1718bbbd26e30f65c464;
reg     [13-1:0]          Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e;
reg [MAX_SUM_WDTH_LONG-1:0]                I30e28a0e32497e3137bb689fdbde46389bc490300e15be88612f28eff07976e6;
reg [MAX_SUM_WDTH_LONG-1:0]                I0b525cae7fe005cf25a07cb0b1486152d726fc74aa55f03480f10af97379953b;
reg [MAX_SUM_WDTH_LONG-1:0]                I3df4fc0f2f099890a34d7b376328da6460d429e2516a5f8fd1aee5a8fee835df;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib1b15c9e15e963cc4f2e9caa1b6b132e338947224b705b51ebe710d7e0f661d7;
reg [MAX_SUM_WDTH_LONG-1:0]                Id364040d3b9f1ebf34ae3fdf7465d955b49d7a2f4709219f76229766d6df98a4;
reg [MAX_SUM_WDTH_LONG-1:0]                I7cd9dadb64725f4217f1330c893724a7537a616ef41d9dc49fd2794125e0dc3d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibdd77bf8b31352e365f7e6440a57247a8ba62e667b000c1347165bb39f3c7c2b;
reg [MAX_SUM_WDTH_LONG-1:0]                I35e7fd3f09acca79a1003b0a4b7ac62c4a2be93bcf333abbfb13a5eefd7d5eaf;
reg [MAX_SUM_WDTH_LONG-1:0]                I7e269b2e2d9ec70c47570bad75bce0ddf53e85e3cb4ba87f784ca520c5ff1084;
reg [MAX_SUM_WDTH_LONG-1:0]                I0c23517b9814053cd1f89a8b80a64fcff6ae65937dc97199c0b79ba8f7a34ff3;
reg [MAX_SUM_WDTH_LONG-1:0]                I73ecf8ab6430c6343bf7596e671ce01a3e3e7499813ed75c583a7103147b0bb7;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib7f659da098e577e33fc0f5da1c03f6d3e68b3883ad7888152d2e8684a6177f3;
reg [MAX_SUM_WDTH_LONG-1:0]                I3386ee46348e8c4359b1ea2153bc64afbe76f2b6bc9a312629b8c52762a22873;
reg     [13-1:0]          I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c;
reg [MAX_SUM_WDTH_LONG-1:0]                I8c2fe0c8cb55f09e4dcdbaa3960acfd815764161f53c6234273dffe4558644cf;
reg [MAX_SUM_WDTH_LONG-1:0]                Idc64cee034c1ee132335ae593844b2c46e3f1b1b2cda8699940df311735a32a0;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c7699448a10638886eaa021495d4c7cc378fe1e9b0aafccda001c15484b9419;
reg [MAX_SUM_WDTH_LONG-1:0]                I45b03b0185f9efbc11c707a64fda9203cc82ec2fbaee7ff34610c74d7cc1132b;
reg [MAX_SUM_WDTH_LONG-1:0]                I3097f16921e899a99f2a2b013a3f6d339ac9672fa5e17655ceba4de2d506e151;
reg [MAX_SUM_WDTH_LONG-1:0]                If0d62663c8a08719b83a27c76fa62525eb14d452d4ff0f33e94c67f58d7c86f9;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifedfb1db4b16b86149f5eb8b0adf06499331d423c368c0077c738a190a1814f0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ice24cd0bd76a7d12a0199df195b34f41f7f72f037177656693b3154d102ba729;
reg [MAX_SUM_WDTH_LONG-1:0]                I6148a04ce3733485aeb6c4d20b6117eea37a510aba76ac29e82d44980bec0934;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6391e6b0ad4d9fe4136b90a57d121f2b5f16ed4662429f1b85677591fee37a6;
reg [MAX_SUM_WDTH_LONG-1:0]                I5dfc39b913b8e0d00491e3f7f45b6b467a517b5e87baa065097e28e6d695500a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie538f6d2c778992e2324a9adbde215acaf7b8dc3a72a9230d4fba2332f3cab67;
reg [MAX_SUM_WDTH_LONG-1:0]                I03929e638a59a35fc0168772ca06f7a502352e03525042ce6d49cf9ecb671093;
reg     [6-1:0]          I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieb5e001b45961175497657da7a0340c2a15b6d8de1b72ad68ac3aa7f96a47af0;
reg [MAX_SUM_WDTH_LONG-1:0]                I6d58dbbb9b18e4b347b34e548c70a9bc0d819986fb3a6bcc3ff8a67c1fce9c9f;
reg [MAX_SUM_WDTH_LONG-1:0]                I82772b528a8c156f2932a23a720f8446f3062e9605839897b4652bb2936fca1d;
reg [MAX_SUM_WDTH_LONG-1:0]                Idb259e613b71ccde839570ff2e7f21a9cb7bf676ffd4aadfb08d6a963bea9640;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie9b1b4412060f1e9acccc1f3ff897bce33f24fea3bfc91266f9e42c1f38aaaad;
reg [MAX_SUM_WDTH_LONG-1:0]                I259a9b6041f341013e6ea0706c4e9ef9a77148bc003b3f0cf9593ebd915b30c1;
reg     [6-1:0]          I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a;
reg [MAX_SUM_WDTH_LONG-1:0]                I41a57b30ab1dd9c40a723f99315558a47412465aa3fe967250572e8373aa7180;
reg [MAX_SUM_WDTH_LONG-1:0]                I42968c25ee2870f891f69991ae3ad8bc1c3acde2f8f4d6c0cacc48f562399c37;
reg [MAX_SUM_WDTH_LONG-1:0]                I44103a07ffcd818c0d9280b96ba08c32f96edc83a981ec9748ed3d6e9c061d62;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c886223618a03ba9e18de68462ddcc522338cd26d24b5e126da9da1df1339f4;
reg [MAX_SUM_WDTH_LONG-1:0]                Iac242fc0dcf37a86cc334319d77aaae46dd223017f2a6489c4e33314eabc9874;
reg [MAX_SUM_WDTH_LONG-1:0]                I3225ba7b6d0e0c7a94dfbc8e074ade02b79a66f6aaf97580a451c2d1781a625c;
reg     [6-1:0]          I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546;
reg [MAX_SUM_WDTH_LONG-1:0]                I25779b63a47c05d4588d4b33fecaff61647609a62fcc90f0f541c6b30ea9342c;
reg [MAX_SUM_WDTH_LONG-1:0]                I05bd9a1d7818f4945ddc448149dee571e80dca8b6eba7ab79b17b6f84d3f35f4;
reg [MAX_SUM_WDTH_LONG-1:0]                I17eff5960d8d41f0832a48fe9a3ae0dfeef1bfc44b73eff506fe1d3813398d15;
reg [MAX_SUM_WDTH_LONG-1:0]                I1b02edd5d00090446500b1dbf66a7e674de978c068b81ff0b0fb7abb9ffb1654;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c865426b0f044469b391bbc13f977fdd19dc89c908574ba289388e382d55cbc;
reg [MAX_SUM_WDTH_LONG-1:0]                I2e557a901de23b8442e8002b3560bbf9cb8592b7bfb7a6e2f8aad12843a5a041;
reg     [6-1:0]          I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290;
reg [MAX_SUM_WDTH_LONG-1:0]                I469f4965961eacfe3dd0cb82fce4905e19e6695d71bec95956e8209d2ae39ba1;
reg [MAX_SUM_WDTH_LONG-1:0]                I6e148041c3612c795f1eb1513a9eba29e0509f02f94971fed189dd9f03d54a4c;
reg [MAX_SUM_WDTH_LONG-1:0]                I2f687e6270528a72aa2f9f9cc0a5a6368f8eef358270329cc40b56abc0e4a35e;
reg [MAX_SUM_WDTH_LONG-1:0]                I661bc8acd80497efe43e3d6fd92bc4107b1ca63eaf162cff5695b35f8d4a7e26;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic72f2f8a61b8ecf8960d476bcf8fbbfd4389e932377679286e7182cc12c418c8;
reg [MAX_SUM_WDTH_LONG-1:0]                I823e337e6437e5ba36ecaf0b1ac6b7a4e74cd2ed7019dd5447355626a8877d89;
reg     [8-1:0]          I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a;
reg [MAX_SUM_WDTH_LONG-1:0]                I1622b11941b00f6d2ecd90320158533a66501a6ddb78defb4464a937f132c232;
reg [MAX_SUM_WDTH_LONG-1:0]                I9ab473d34fac3327f03768e14c7bb20056aa8a3dd31520d385552eb6d214f890;
reg [MAX_SUM_WDTH_LONG-1:0]                Iedf1b21de2a0eb04c4a64f9eb34e2b0b3a152d90b1938b61ca45c880eab16ab6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibe3e6de02f0c30287dd89b07be5254ff70d9683389574d02f1423e792bd2d534;
reg [MAX_SUM_WDTH_LONG-1:0]                Iad8ee4f6cd13a9f415cd3519de0179a66cfc993a840b3101cee554b55c0e7e7a;
reg [MAX_SUM_WDTH_LONG-1:0]                I15123100f4377e14c62cf47fb1fb652badc3bd0e8f0ab4b970a0bece065a6380;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic0a892c18037ef674c8d94cdfc94cfca47d977ca2da9e678303255b96575f022;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c316e8b8cb6b499a7a8fbb513b3067829197cfacee877c35874a2ec686ada4a;
reg     [8-1:0]          I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib3a2af9bef5f5d8d7228a3b49a5e0d4a37a33117e057078a552588a24d46addc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia042bc20eb6866de0ab9ca9154f0db63f7d4ad84d553be858a0be88fbb8f7f33;
reg [MAX_SUM_WDTH_LONG-1:0]                I5b4ba308b0fc2946fb11b66aa5c24c7b5cb2a21955116b97f3790de65cd2a064;
reg [MAX_SUM_WDTH_LONG-1:0]                I005ecc3a38317079c7bc5008817e11017c33671f77364ad9a07d0eff1e0ebf0b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib63856036797d30e60f13453da509ace15e3324c25bdfdea5aa495d592e2006a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia9bf10fecfe62530ea6be4687ecf78a2ac08c6fc6e38328c2d64a80cb5a3d72b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie1447c9e1eb4ed110e6b0353bc5dd2cd14ec645355c3cf897df6f6c5808475ad;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic8f640e7a0c71ddb20a985259b5e48746d28d2898383765c3b78c577f281d27f;
reg     [8-1:0]          I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b;
reg [MAX_SUM_WDTH_LONG-1:0]                I3b1d695a626aefa8e5b146c7f7f26a8da119680783da7afb019209ac9fd719aa;
reg [MAX_SUM_WDTH_LONG-1:0]                I1d91c7e9c2f99df4e0523b7e01b6fa6ea3930382238ccfbc07201b7d3edcc969;
reg [MAX_SUM_WDTH_LONG-1:0]                I7c1e9623dc53c8aa8611b46c0375994510a97c4d49d0b091964cbe4671acf1d6;
reg [MAX_SUM_WDTH_LONG-1:0]                I1b5d096081c0190c0ce6a674de1afee9ccd766a9cfab0637a0aec33199061bbf;
reg [MAX_SUM_WDTH_LONG-1:0]                If145a331c8a8abde8c26d2571cc8b38e1eaf2768a4658d350cb602bf8614a521;
reg [MAX_SUM_WDTH_LONG-1:0]                I86e764dc3320206d9b52013c2d735ff4d27bf6e4a82227486e64b4ceb68dfe8a;
reg [MAX_SUM_WDTH_LONG-1:0]                I4a98524c02346f4b9468666ffaa9d996b9b868a5a8730264d798d7a66b7454bc;
reg [MAX_SUM_WDTH_LONG-1:0]                I1187dbcc72f33b4cc3442982af526be4cfca1b5ac65be943d4ec380421632117;
reg     [8-1:0]          I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f;
reg [MAX_SUM_WDTH_LONG-1:0]                I73ce2860dd9aa9ca2c0d541a6ae1e5069badd35988d922cffb6aef0038cde662;
reg [MAX_SUM_WDTH_LONG-1:0]                Iea2dd4d33966d53ae739a16876ac2cf04e1d95374a5af68e59a5703dfef2aa79;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic0a386f5301913434a3d6aaea1d56d6acb3484fababb7b8831d09563bd8842cb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia8a4fca33add1c3c58b04eafe9d023751882f409c5d2905f77aae3fef8c2b008;
reg [MAX_SUM_WDTH_LONG-1:0]                I9cd4ac82c1e6f2dab27efa85314df34a40d8747959eba18330bd424a38debece;
reg [MAX_SUM_WDTH_LONG-1:0]                I9bcd5f3f4630ce7a24ea4479c9ddfce59ed809dfaad9d767e80295c41b332f4a;
reg [MAX_SUM_WDTH_LONG-1:0]                Iac7a05e270cb898af4ba32c16445d0dbdffdafdcc5fae209f09367abcff9d6b7;
reg [MAX_SUM_WDTH_LONG-1:0]                Iad7f008b5f08f3ba94a0832261fb4add17f0897e3c7d54a250377b813e284331;
reg     [9-1:0]          Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic072a2fb2ce65ca734c05e747f12ad094cc5aaf9267dd94dba345b5c7b11dcdc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic20328b806ccf89387180fe6d88ba762051c6bc2c7f82494129e8c3600108804;
reg [MAX_SUM_WDTH_LONG-1:0]                I11855780f53e8711f8eca9370af31f472dffd126c02cfce8154a959f33c68af6;
reg [MAX_SUM_WDTH_LONG-1:0]                I39b8420e976cbdf011232d83446a5cb92c2ba58577792c9c61dd71358205e936;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibca01267ba9d7e2fe9f8df34a548836390ba12b9b782f16ba40965c00735213a;
reg [MAX_SUM_WDTH_LONG-1:0]                I105a7d84244a0d9143b9b2a3c64ea6964f7e1f43b7f8f5cb15d579885bbf746f;
reg [MAX_SUM_WDTH_LONG-1:0]                I1b0f11f3bca53713a53e2ed18fb81f5a25c7151c874be612677f5204bca28093;
reg [MAX_SUM_WDTH_LONG-1:0]                I434991f7c09dac3a7bd42fce3073dcbcf8b1c6579822074548ea94fdf1ef4eaa;
reg [MAX_SUM_WDTH_LONG-1:0]                I7fec897140c79264b7b7b7f3ae228ed090ff69351985c07d317ff9c0cab1e58c;
reg     [9-1:0]          Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf;
reg [MAX_SUM_WDTH_LONG-1:0]                I82bc7aad8e3adf5b7bd03d9fdac6eea60cb800e4502e3af7bdc9d49139563fd0;
reg [MAX_SUM_WDTH_LONG-1:0]                I218ab164221d559f1e8bc2a13f06a7593eb4133134762698eec270be5d4c3906;
reg [MAX_SUM_WDTH_LONG-1:0]                I4135dbaf658fb73b41800cd275824d1c9f410ab1b6e555b6c4c8df12f96c5861;
reg [MAX_SUM_WDTH_LONG-1:0]                Ief38674752576e92e90fbe2a7abcfc952274123875a95657dd42c910133cccde;
reg [MAX_SUM_WDTH_LONG-1:0]                I783b89f0c1e5463646e0fceb976f2b27aac523a677eff6e597e434672b0daac1;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib0ee967a174d7c841ebe71e144d6303bfc80a6083ff6ad745c76d488dea66d9e;
reg [MAX_SUM_WDTH_LONG-1:0]                Iea7b69c43ca4b3707d3bfddf19b27616b8686df915734ba86d3685127bfbf39a;
reg [MAX_SUM_WDTH_LONG-1:0]                Id36acaa2c9161668c95e2cc3e6e852e9243ca7f486ca6c2ae4d124b1a8ddb522;
reg [MAX_SUM_WDTH_LONG-1:0]                I325ec6d7bab5ccd6e9c4a7e9b02a3b8c30072df123bf6318bd97f1e8766457c8;
reg     [9-1:0]          I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4;
reg [MAX_SUM_WDTH_LONG-1:0]                I07c37e958136be68b3d658649964c73ca78160582248da1d45eb9ee82c1f679b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie17e17c22c7215d0482ba310638db13a96c0943216f9ebaf53c0c29c69971b23;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie44aa17133d02266160c8fd6f75716f8bc4a3775356cd1ef0f495b13145ba864;
reg [MAX_SUM_WDTH_LONG-1:0]                Idaf1699bc7916d99a2a5ce0174383c189dca6d7537734b19dc379bd634d0d209;
reg [MAX_SUM_WDTH_LONG-1:0]                I64aaf806ebf0ead2a4836251dccd62a394b984823592340be94f4ea02e12d766;
reg [MAX_SUM_WDTH_LONG-1:0]                I152b3a1e710e5a39bac6338591c6597ee2a38fc25555f563beb7a1a967bf4e94;
reg [MAX_SUM_WDTH_LONG-1:0]                I9ede22dbb56f48c045a1b5a05945124fb97b6ca7e355dd8d9dcfdef6e623b953;
reg [MAX_SUM_WDTH_LONG-1:0]                I30e30c2bee3bac86dd68fe8364f818ab63e91d65c4fa1ef45fcfd03c9df87cc5;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic0bef9008769fe36d726cf80506004d66e7c843a046653201c9bc2c816115c28;
reg     [9-1:0]          I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e;
reg [MAX_SUM_WDTH_LONG-1:0]                I252a77c3eaec2d6accaee6de3ba5d0b354636e2a2aef4992eca0e2a74eb4d25f;
reg [MAX_SUM_WDTH_LONG-1:0]                I5fa628cdc28fdeb96014a4d2c2d06b092136cf2a14a0420bd5d3861b83687413;
reg [MAX_SUM_WDTH_LONG-1:0]                If258ff7e66143201e30b3fd451e1b8e2ec9e46596c2653ec836617c093f28018;
reg [MAX_SUM_WDTH_LONG-1:0]                Id160a3b60a3c7a3ad93044461ade9ccf0b7a627efa4b1bba84a2ea0d4fbdb551;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia42e25bf722566321268c83de181d196619f062381c7fdb381ab5f6aeba6589b;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f96b4022f127e7d965786f2cac8ee6afdbee96980608c876c6b699495f80b0f;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a2505f0de03f3e2d303fd207ee819f5a1777b650930b87a235ab3cca5de6e87;
reg [MAX_SUM_WDTH_LONG-1:0]                I8600d4c5861319be0efba19d9b66ad483aa7bf648f2132c1a339157c43920c18;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic551d228c593c4304b4ef79a965ac1d9081774282af09d79cd587ef9abcd6003;
reg     [16-1:0]          Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe;
reg [MAX_SUM_WDTH_LONG-1:0]                I01d7d3d20ba0eab63d519ae054b6c22c5be4000c846a6a4883ffbbddee37663e;
reg [MAX_SUM_WDTH_LONG-1:0]                I4177cb2b0a83442a271f59bf4f758851d5146ee00d76a1177c9a34d4208b7c09;
reg [MAX_SUM_WDTH_LONG-1:0]                I5df828301af902c72794032c0e55d8e7548c9b2277b2edc77f53796ff8e04804;
reg [MAX_SUM_WDTH_LONG-1:0]                Id595e96924941a80a6ade8778fcbcef39b07a62fa1d7350fe50182fdae302556;
reg [MAX_SUM_WDTH_LONG-1:0]                Iefbb3d08b0b2fc51d2f6b60b25b8143f3f88a705e770396e2f6d050632ded97e;
reg [MAX_SUM_WDTH_LONG-1:0]                I71c3a88492c33461f93d43680f11eae8ef3e9402a4b931c5d31f959a2f8c147e;
reg [MAX_SUM_WDTH_LONG-1:0]                I7a7bbb1d7d9b77199c0b29fda08f8a63112052ffb0a502a05586ced336e13c62;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie1657c5216d7c6e743a23819c08b7c7f2fc8a56793e1bc67fa5c5f3b37976641;
reg [MAX_SUM_WDTH_LONG-1:0]                Icac36c9706c9e063b771faf556f6699e280687be228aebf6ce71f5ae775a9754;
reg [MAX_SUM_WDTH_LONG-1:0]                I8b3bb7a4701d3ef22c71a9631482e13afc2ff80f40e2f0ae75cb2211af5ce6d9;
reg [MAX_SUM_WDTH_LONG-1:0]                I6a24b9c3ea194d09d619dff007c4c6f53a3cbbbae5c9d3ba718bc3546eaad989;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic7af968d25c444d210ebbc7ae563688f4f8a48f38035ce5bccee100e10555047;
reg [MAX_SUM_WDTH_LONG-1:0]                Icb61d0767612534695d9de0380a1febbda612604f373afa55f0339c7a679e99e;
reg [MAX_SUM_WDTH_LONG-1:0]                I58d2fcb7085fddc9250ca075b010afdc2d019c4091f5d115d9520586224a1ae8;
reg [MAX_SUM_WDTH_LONG-1:0]                I4e5dfe1c7112e24769a5e6aa86584c09ed659fa5d05af38d18183db31189a3a7;
reg [MAX_SUM_WDTH_LONG-1:0]                Iff97998b0778cb649d03228ed3acc81c1b3a97f6bc47041c423120b1311112d0;
reg     [16-1:0]          I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35;
reg [MAX_SUM_WDTH_LONG-1:0]                I422fb05bbac12ca5df13eb7c0c3fd96a4e819de9669ccd64d40060b5db3f3421;
reg [MAX_SUM_WDTH_LONG-1:0]                I782d29ca9e53ffe86cec8809d7d413c9c5ebd9edb6a0d76db2d0c321312d224a;
reg [MAX_SUM_WDTH_LONG-1:0]                I0705e6f1954b14f35dd7fa8a64370c2f9e6e39b6e265857e72946815d1f994fe;
reg [MAX_SUM_WDTH_LONG-1:0]                I3f9e2f1be98a5d14a8b79b252e9b5a2b3a09304f27a3526a4a66b365b682787c;
reg [MAX_SUM_WDTH_LONG-1:0]                I134dfd9d579ba8b2d72bf1c47119a086fcfb6b7d591cc2c5558e451f57636d0c;
reg [MAX_SUM_WDTH_LONG-1:0]                I5f4870fc880aac0f84130a26e3cd493954ea49eb3804dd17a91b2ba1cea599f3;
reg [MAX_SUM_WDTH_LONG-1:0]                I918037e81d2f9c05c6a8b94c64724b1d0ec8afafe5666df433fee3e296171f54;
reg [MAX_SUM_WDTH_LONG-1:0]                I136f70cfdde5473f8944efa2b1093ed76f82dd06a341413ee2a56054ebef5fd2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic02dae50f30bea04d63949eadbcf892ce936efc5373a6185668a20311dd59f4f;
reg [MAX_SUM_WDTH_LONG-1:0]                I54296c97ecd9a699f171f4d7271c761aeea50255010a0a90d2dabc16a0cbef79;
reg [MAX_SUM_WDTH_LONG-1:0]                I50a310ea41e0637bf28b5f56cf11560bc936e15c73acee063c60668bfa905fed;
reg [MAX_SUM_WDTH_LONG-1:0]                I25d2b0d3ff7f684e508a62271f3d29c729dc46478248627013dd91075f8d2146;
reg [MAX_SUM_WDTH_LONG-1:0]                I7f9f83601cb61fece60f94c3120b43ca0c737ee36b8c67ccc917d3a428d8750a;
reg [MAX_SUM_WDTH_LONG-1:0]                If4fa37977e1db59d1bd7a30b2b0919c997b6e25e0438e01b62dc273d10497867;
reg [MAX_SUM_WDTH_LONG-1:0]                I66291192ca8d81c8e3f667651d5201cb41b6872f73283d13c6718159b008d8cf;
reg [MAX_SUM_WDTH_LONG-1:0]                I4bfef3f43cb1a77ce8b2bf4b26160a161e7f28308b8d2817e6e2840f09463e37;
reg     [16-1:0]          If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad;
reg [MAX_SUM_WDTH_LONG-1:0]                I0aafab9f9205eb4a8c16e213e116d949a5c625f7cb2b0f3d124deb80aad2c6c7;
reg [MAX_SUM_WDTH_LONG-1:0]                I9095fb177f965807ae5a73a45c76b1c0b6300c6800b17259e5836adea5a78ec8;
reg [MAX_SUM_WDTH_LONG-1:0]                I3780e5266741d9a9435818f002588f4c44ae518b77a30ede57a3823e1e1e5867;
reg [MAX_SUM_WDTH_LONG-1:0]                I360ab21cba3dfd419f0ca83f85d9633b918c3d24a00214399b0465d7106466ad;
reg [MAX_SUM_WDTH_LONG-1:0]                I2c061ca6ba4299d676b5c6f1e1cc920bc1104e7ac730d207949b952d1a98300f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ief44fc6df0864dd0766877e0d673847250f53ab137cd9029916ab7149446f9c2;
reg [MAX_SUM_WDTH_LONG-1:0]                I353e1673347daf260e61fbba813cd14f83c52ce3f6e5168c0fa6308d41e93590;
reg [MAX_SUM_WDTH_LONG-1:0]                Idf77a6217d51b2439f71afbf5956a52a241f2bf8722f54cb166d83c3b45f6721;
reg [MAX_SUM_WDTH_LONG-1:0]                I8ea9b55580c15fa584fb934e010debd92e2e893630de456e85036d583921011b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic36cf3da50983e4168cc0a31ec0a86c171714355c0fab18398b8daf57bee1a45;
reg [MAX_SUM_WDTH_LONG-1:0]                I7469c1791d81d0924eb0faa6303565dc78fe9eb371fa13039ff89b92b7f51a6b;
reg [MAX_SUM_WDTH_LONG-1:0]                I9b8a4dcee9668bb71803c25e0ece0eebbf704eb29cfa7b91c47cf48d61076803;
reg [MAX_SUM_WDTH_LONG-1:0]                Icf4d3544466d430d71abf2513cfbc16b575af540d369d405ed831753f304673c;
reg [MAX_SUM_WDTH_LONG-1:0]                I0568efb50e0bb85c39c9ac6d2ab3474ab38799257dac5693085eeb0d74859ade;
reg [MAX_SUM_WDTH_LONG-1:0]                If072f43c0b06c41c30d9bc40dae674ad9052e5533b1308adb97cff2e03821bab;
reg [MAX_SUM_WDTH_LONG-1:0]                I2f05dd0209278c1e661998552da73728c1521c024a7d26f4652d4f151c6e5f80;
reg     [16-1:0]          Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c;
reg [MAX_SUM_WDTH_LONG-1:0]                I17dbb17fb2770beac552dafeb238c5e8e7a948c35c7c543508e652cbcda01dee;
reg [MAX_SUM_WDTH_LONG-1:0]                I68ed84b705e3c00d0fb66182d6eeb93f43999532d713f81fab39a36259e0e7da;
reg [MAX_SUM_WDTH_LONG-1:0]                I9d1a378e4d5703b65f197cb76a1982cc10e0c17654eabcf10d9df091086d8acd;
reg [MAX_SUM_WDTH_LONG-1:0]                Iba503643311c9dc3366b9bb843dcc1ee2f0243c4cf78004a660fca224b36c5f2;
reg [MAX_SUM_WDTH_LONG-1:0]                I05806fb5d45e4d6f569c12116644b625b7ba071eb052ab97525f06fca03dd88b;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib2630bec8f9f78489ca6cfe0bf25746b720aa422b9d529d67d6dde2d045d9c3c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic57569daaae5eb0e66117615c8c6043b5f76b114b5c34b0df50445f66a22849e;
reg [MAX_SUM_WDTH_LONG-1:0]                I5cbbcfd1cfc35b3e78d01b29831195106ebd9ba5907f44dee6761c2b047c4a60;
reg [MAX_SUM_WDTH_LONG-1:0]                I6dc5ebe003a649f0e4106dc27f25387651d43259f0ddafad10411795ee48b40c;
reg [MAX_SUM_WDTH_LONG-1:0]                I238a5c9cd1dcce0d745817081a4b240f74de3de6f18a3abcc42cafbb19a0ad69;
reg [MAX_SUM_WDTH_LONG-1:0]                I53c29303c76ac3c1c02fc9a74eaff9595153ba06d67c08e07790c58e53b674f1;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia92993e9a66294adf7a4dbe1ea88a9e8be6367da1c05b8df343b3c7a38bfd8b6;
reg [MAX_SUM_WDTH_LONG-1:0]                I329448311438699d3d590bba6ab4bfc9cead805f96015b77617f42d957bde7d5;
reg [MAX_SUM_WDTH_LONG-1:0]                I717aab2686adb8a0688009c23d92aa4475e240ec0747735e6fee5e196a50c444;
reg [MAX_SUM_WDTH_LONG-1:0]                I13a54b612481fe0fdfe8b52909179bb82298c2bff4f10adc4f41215fa4396311;
reg [MAX_SUM_WDTH_LONG-1:0]                I26a27b64a7aafdbcf4a6d058181fb84e0e16767f4bd7a9c45211c4c1246d3b9e;
reg     [9-1:0]          I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie46448d24890ed6ffa2736abb97331dc3ed219b9324bc0e8453eed6aa2a4806c;
reg [MAX_SUM_WDTH_LONG-1:0]                I8ab86da421b01a03999daa91e41ae95ff58c6bc38566a3deff72633a5ad1cc18;
reg [MAX_SUM_WDTH_LONG-1:0]                I20ddfee724da47731a2062b2732598b429c42f7d22bcfb300dc084de362a2bdb;
reg [MAX_SUM_WDTH_LONG-1:0]                I8d8dbd62189397b5e9189ead2126a615d5b6cea393901e21cd89c255d6672615;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie79db7f22cab9cd57482ce0141d83d5c1ff720a7c3dca2c3664feb4a1e2f4850;
reg [MAX_SUM_WDTH_LONG-1:0]                Idcdcb2dd5e2f2aff0d7b362ddb4ae1ee4db08edc2c3df3589a7143bafeec0bcf;
reg [MAX_SUM_WDTH_LONG-1:0]                I525b9b85b14df7a6533a7e54bdc9bf40a303c890a4a410251c8d556d38b33125;
reg [MAX_SUM_WDTH_LONG-1:0]                I65afc937c55081dabf16dbfd02eb03c97204efbdcfbb523609571bb32d537d5e;
reg [MAX_SUM_WDTH_LONG-1:0]                I45a11cd2f581121ac03fe112ec78bd07c070673712fe6112a3e4fb4eba298e27;
reg     [9-1:0]          I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3;
reg [MAX_SUM_WDTH_LONG-1:0]                I9342de9fe82f2273da138f99da619acf144edf1f9c33682fe3b1a09d0121c4d1;
reg [MAX_SUM_WDTH_LONG-1:0]                If6cd81d168d83d5f6a7ca18051bbbcea5c7a9e017cfffcf72f31f73275c3a4d4;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie2c7966ff2c1e84a7ae016f31b0f8b9ca7aa42eec03467c7e3dda37dc34f070c;
reg [MAX_SUM_WDTH_LONG-1:0]                I468b28bee4fe1c0d20fe7abd9338bf844ce0a2e322ed6b6de11e2ac621572c48;
reg [MAX_SUM_WDTH_LONG-1:0]                I08c55e08731cbdc9703e607b481a65177e7e1e242fdab9bfb014964bb0d1d22c;
reg [MAX_SUM_WDTH_LONG-1:0]                I6c252caff8f1ab047efc25a950ce3e3ffb47a5b779e37a667c48bc1487528218;
reg [MAX_SUM_WDTH_LONG-1:0]                I2ade6ee1b52da04fce9491cad314947a07eb9aaa8b0a430db2f96e2d290384dc;
reg [MAX_SUM_WDTH_LONG-1:0]                If6e953221a61b86b1fc339b69af853f6ad538b60770f2f7b880d7aa15bd625b3;
reg [MAX_SUM_WDTH_LONG-1:0]                I6c6885b180013a16955ddefa0dc75c25ac85fb76059df9bf8b63af72c8c1fb4d;
reg     [9-1:0]          I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42;
reg [MAX_SUM_WDTH_LONG-1:0]                I907aa3f6584035b934017a601019d35f353b3f99c7573bef60fad167f9d9ffe0;
reg [MAX_SUM_WDTH_LONG-1:0]                I7ae7cc2f052d37b650c0abeccd841b1b18abb4049c976fbdbab72ea579a5d206;
reg [MAX_SUM_WDTH_LONG-1:0]                I5c0776e9826af1a98810296a7cb86adde5b1b41c434e6040bc6a5a30172d1bf7;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia244be7d571a1e41348c37534a23f7cc942b689cbcd5dff8c10043325b80e322;
reg [MAX_SUM_WDTH_LONG-1:0]                I14730b2825dc07428388347472491ef3abe06da3bcea9b7dc9c919079c22325c;
reg [MAX_SUM_WDTH_LONG-1:0]                I22670670d7018cb361ca0ffd92516837302d5528c26915b62d22505471ab7384;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibc34c6979b8f5adc5421ca8603b6dca91161055286758ac10d0c612263077758;
reg [MAX_SUM_WDTH_LONG-1:0]                Id39c55c4f0df8a0d8ee4f8b47f3de8cebf5343bf75521edfe38a695565eea926;
reg [MAX_SUM_WDTH_LONG-1:0]                I06a5cdf2e430e40b5c08ab617356f6b4b0389236041b77e2a57d9d314bfe77f3;
reg     [9-1:0]          I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d;
reg [MAX_SUM_WDTH_LONG-1:0]                I22c3d90c4ad5f41054f9b3dc7ddae143f567182c7fc695c5cd087f126ccdbcf8;
reg [MAX_SUM_WDTH_LONG-1:0]                I533d6897ed500a803f6f6468e36a2a922495b3effbeb405b47ffb7a5f4d82c89;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib8d3655f6360b2b189b79353d38c9c9989af811109144d45af0f8b68a3276149;
reg [MAX_SUM_WDTH_LONG-1:0]                I6b264ac5221269381b155a30c051523f4488ecdc6eb2cf60da80a8b84c49bd96;
reg [MAX_SUM_WDTH_LONG-1:0]                I5c3a945e8bd4c55e9cb38d19100b13668bd652bc1162d16b30f1562a6595a032;
reg [MAX_SUM_WDTH_LONG-1:0]                Ief691d56b56a000651b0a4c6cc9f26bc44da82f4a6382550d96ea4101b81ecb9;
reg [MAX_SUM_WDTH_LONG-1:0]                Icf55933dce8b9f95a57d7d019c9b29f72e08454428013009cf0e4d2c5b6edf0b;
reg [MAX_SUM_WDTH_LONG-1:0]                I5b0da0701e7399ca2e668c1602f494f41127e4c90e6fa91632da0016e7b395e9;
reg [MAX_SUM_WDTH_LONG-1:0]                I6106f96669a63f337b78a6bad5894881230f0ab6467c23ec877cf27a5bc76cb6;
reg     [12-1:0]          Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1;
reg [MAX_SUM_WDTH_LONG-1:0]                I566a76fd27d46125a614f5e0c72dff06a0c1d836c7fe4a2c4086129386b34dde;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic754ed4f2d29b948b422876f371df4f89b86976e25183ce1b9f664e1a9b19f56;
reg [MAX_SUM_WDTH_LONG-1:0]                Id7310932ca8964fd49adc052220c04855b028e29fb7a48521a36e2dbe1d6d5f4;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibae8222f76059e8f61dff938a64e23080eb668880ac50ecbb50de852472a22ad;
reg [MAX_SUM_WDTH_LONG-1:0]                I09673e64aaf6f35dbf4aae16ffba969d08a800d32ab25413bfcdbd540d7b01f3;
reg [MAX_SUM_WDTH_LONG-1:0]                I3ae1a42457a669272eeff1bc293c80c67239ef6b725a09eacb82b06ec84edd65;
reg [MAX_SUM_WDTH_LONG-1:0]                I5b4c4554a78c551dd34a93ceb225237a2d2540a0e05311c4595bdaa5a4cb14ea;
reg [MAX_SUM_WDTH_LONG-1:0]                If27288056468d3ef3052303952f2e4be67796c40d6224383047d71d996f98cf3;
reg [MAX_SUM_WDTH_LONG-1:0]                I12dfae8d4c1a0612c6d65c6f5493247af5e06ca1d8c72dc28f9ca41b0bbc6ea3;
reg [MAX_SUM_WDTH_LONG-1:0]                I295da244d8dab1563a5947230e49171eb905c3758c289526ff6d3e0c3efcebbb;
reg [MAX_SUM_WDTH_LONG-1:0]                I89cf2ce418b6d96c0e2b9c8e82167a47d40ade45a8f08255a1b849a9df9e6d06;
reg [MAX_SUM_WDTH_LONG-1:0]                I47ba4d6ad7b1889cb52ff7a1d42176e166270e39a1d2875f3a0cd260a1fc92ab;
reg     [12-1:0]          I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4;
reg [MAX_SUM_WDTH_LONG-1:0]                I08240dfbc0f698324c1ffdb8e769016bb8b947fb0b8dbb72839375cdb4cc47e1;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia9ea47bb0829c979af002fb7aa0e22072671c2876bcdf79365ff2b3691172149;
reg [MAX_SUM_WDTH_LONG-1:0]                I58df4f7ee4282cdb7bb80c9f1d907ff37590b1db22994f3a07b521132ab80087;
reg [MAX_SUM_WDTH_LONG-1:0]                Iadfdcb3c0764107a2b0deaaf039babe6a08f1018f3718f5539718ed6a5aa962d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia2417744c8f15898d5d951e15cdf8c03d932cdac6acd27e32045e0fbfbfe4f30;
reg [MAX_SUM_WDTH_LONG-1:0]                I6d70d8c6d44eb58daff53226cbb59eb647b6dec6bed37021a64e16ac5318d484;
reg [MAX_SUM_WDTH_LONG-1:0]                Ice3b06f04279add8283c8173340c2bfd4b4801d85610179943f070aef508a893;
reg [MAX_SUM_WDTH_LONG-1:0]                I4fa5ada2d589c7a90e700745aba8e09edcfb0252f532e4c74eb0809c712a36f0;
reg [MAX_SUM_WDTH_LONG-1:0]                I71c6f88cbabd48d41f42f2b16170c8955b79d20b8a8b211e174d1c1473567ad4;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e7e130607ec849c80f9e687f0215ceb767a2650626f20ee44a6fe677fde2299;
reg [MAX_SUM_WDTH_LONG-1:0]                I4c02563233638e273f05bac3e277c702b38c204fda200dc5ac163662c77a429b;
reg [MAX_SUM_WDTH_LONG-1:0]                I85d8f259f770b22a380d6eb5ace0281c57f0952506152be05f38482c47334988;
reg     [12-1:0]          I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b;
reg [MAX_SUM_WDTH_LONG-1:0]                I989259874d3f12b373358db47fed6245f192edac9e7df00531ea7ba75c360d4c;
reg [MAX_SUM_WDTH_LONG-1:0]                I2ef69d9eec4f925b598115d569d2d85a4545871f2ac62635f9b072ba718b595f;
reg [MAX_SUM_WDTH_LONG-1:0]                If8cefdab8d831c3db83e1ef615ca534f34c58b9903520c7741cafbc84e28d207;
reg [MAX_SUM_WDTH_LONG-1:0]                I00e5abb30adb527f6b32257212dc21f9797e9793ebbcc10feae9e524188539d2;
reg [MAX_SUM_WDTH_LONG-1:0]                I9349cba960e03e6068aa27e997993b0c466e040a1ee9e6053536d3346c84214f;
reg [MAX_SUM_WDTH_LONG-1:0]                I19797110801d39a7970e6d8665215c967071ad9a1bad12c33401b44f595772b7;
reg [MAX_SUM_WDTH_LONG-1:0]                I0d25b3618b50ff21e3f301fe44087368e38fd6b37b6f6fab004824aa9df51f0b;
reg [MAX_SUM_WDTH_LONG-1:0]                Iba62c53d136b455b7d575b868f2ebd2dadc6003981aa2aae72863a0eb812bd1a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6f2e4979fa9229a647a81a4fa3f8b2af809199049d2554ea15fa9a6ba2f90a9;
reg [MAX_SUM_WDTH_LONG-1:0]                I83d70d4886f48dce0888e203c2c333c76d35f0c73767dd9443ec8fa4790ecb09;
reg [MAX_SUM_WDTH_LONG-1:0]                I3f92074e96f2c2711248b1d770b4ad718a565a323e6fe4ebb379e6494039af47;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia478acf4034b69d392277c3d5c6683346547ff26d418b3a6c36a3f9a56e3cfe0;
reg     [12-1:0]          Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021;
reg [MAX_SUM_WDTH_LONG-1:0]                I06186aec49594899011a9d7bce163a3a43ec094d7c92033df033594ed5eb43ac;
reg [MAX_SUM_WDTH_LONG-1:0]                Icd8ef17fc44642a3c86a1cb62727eb607e3a4e6d0b021406b9b710ea5c96c06f;
reg [MAX_SUM_WDTH_LONG-1:0]                I2a3d1a32b282fd624497621815c6ff85c904f5f3fb50f18cf345c5a5d7a557ef;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibb57ab5a5468d08c8b299ee67b535b83995e94d6223d0c6d93dba8580906e319;
reg [MAX_SUM_WDTH_LONG-1:0]                I6fdc128e94d85f0f7f884ee1ff44fdb6de2ad5b93d83c3e36ae235afcd3d23c0;
reg [MAX_SUM_WDTH_LONG-1:0]                I2790277776fa84c3edba2332cf538f8ea3a40c1b06cece7463a3b4757b1fe213;
reg [MAX_SUM_WDTH_LONG-1:0]                I068f00aade8307d2a2e2ddb37d7429a04c2f6786232134a041e62733cadb03ac;
reg [MAX_SUM_WDTH_LONG-1:0]                I07087056bd31363bfb1f76f8fbeb18d1deafd5e4816ca1200d362c0797a77bb4;
reg [MAX_SUM_WDTH_LONG-1:0]                I01c264f9a89aec9dc11fa16206ffee1c8fb03bcb279e9e9f53fea1e94e9d8b23;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie42f89c20abd223240a9f93a89ce650ed2f581e1ceab0587a4fea2ddf9f4f98f;
reg [MAX_SUM_WDTH_LONG-1:0]                I44ba42cf2460fce5fde6d8a9fba799517336268d29b5817597d819a9eb83df0e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie4fafd34aeca2efbfd3bfd3bf45f73ceea27b613ed242a43666d85f3680ada44;
reg     [1-1:0]          Iea53e5522afe762dd4185f0262512abbb94b905893974c13e954df5553942b1d;
reg [MAX_SUM_WDTH_LONG-1:0]                I65cb4f1288affe61a7cd9981878d8519db25d724cecbb80eb3932ccedafcd5bb;
reg     [1-1:0]          If481e9fd41cf8181d432f397381b8376d9da7ddfba17b52e65e301e74c3b9b0d;
reg [MAX_SUM_WDTH_LONG-1:0]                I577e642ba232b9a606abfddc4d84ce4354744e2f953da3b285e417dbfc5aef16;
reg     [1-1:0]          If2e4ac195be838db9dd7b062319aba299887896862f1a340013226fa025b18fc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic68515eee7d422be9cf8950e48b81d743d5491851d5a117d1f9b70d1d9b55060;
reg     [1-1:0]          I40914301545dfe0b6673f76e0dc0d1ab3968ca3b18fe8f4ff63d5623c31bafa7;
reg [MAX_SUM_WDTH_LONG-1:0]                I0ca47358f982879bb85bd78f6bc19192a5ed8c62214073342b37b040aea331b2;
reg     [1-1:0]          Idf30e1a70a723113d32f621f0375dd85270da2f7386cff5ef4ff88cfca78b848;
reg [MAX_SUM_WDTH_LONG-1:0]                I1606027ef88387f2150285b55cef89212359f49ab1a49fb71e457a3dba0c438a;
reg     [1-1:0]          Ic246bc24fb918b7c4a32727a332df57bfb205adc05150ae8d944a77cbdc62822;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic09f51154140ef91861243d7b35f05961565b368264d44c8fd5d0f85bd0fa213;
reg     [1-1:0]          I6cac9957a16e7cfa8a125b40d8ce42cb7f502078a791b177d9bbe9589b612426;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie28425115106f4b2405fad6fb2994a76e64dfa60e7bc165f46ae67411932a1cf;
reg     [1-1:0]          Iee4ad1e7709a56d53cd8b97f587f1f791fb88bf278fcfef32a29fa05247ca13d;
reg [MAX_SUM_WDTH_LONG-1:0]                I64862889bfd7d2a15503bc07af594be59cbaa8758863f78311d6f15ecadcc99f;
reg     [1-1:0]          I16a4499c48e5c24fd8a6d49ec3bf63c20c85f440c0c897cdb840e9f28fa2e68a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ied4424f3e85f3fb92f4e40bc63909f4e77698a18a1d0ee651e54e4de06ee330f;
reg     [1-1:0]          Ibed209db0bc502e3fceb4ab86ac20a2ebf87c43391a546d592e5aa32709aa8bd;
reg [MAX_SUM_WDTH_LONG-1:0]                I6c850d46af2f31f4e3d31c3fd2b2d9c7471ccf817b452a4fa2602485f5e7f164;
reg     [1-1:0]          I05dc9e8db597a2123632b2934d864ae64cab5192401d8f66ebebd95618590ba2;
reg [MAX_SUM_WDTH_LONG-1:0]                I1a1a9f7ee74e17c4a0d7064ca9fae938002b1b685f3cb6309569081b0d971aed;
reg     [1-1:0]          Ib309786164a7d646c17533008b3aaf0fd86eda3c5ee167efc2080ef5b26a9ddf;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib5929b32be13a8436b74dadded1f26d3742e1424b6025d1eacda112bf4749a15;
reg     [1-1:0]          Id9bbd0f5c16ba0ffae6a0e5304e1726b97df06f06feaccbb1bbcaf0e01be3823;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibcb7809e1db6cb82ba62be017c5b8685cb6f988f85a0d29ce2459f6ac80498dd;
reg     [1-1:0]          I4294b001f220e009c2a65fbf8b36ce1d8961c317ae8ded31cbe5aa288191e009;
reg [MAX_SUM_WDTH_LONG-1:0]                Idb971d0017094cf8b28e639623f85e6e5fc2c03a1da1e19a1ef87b959fe8e1cf;
reg     [1-1:0]          Id1fe66d1340965020f513e73a4f77d18f4703c194c3954d40a7f1bc37fc1342b;
reg [MAX_SUM_WDTH_LONG-1:0]                I89373d12365deb440d5337a2586fcdab81347ca28ff6f261a12e35a235bd23c6;
reg     [1-1:0]          Ie95c9af987f352eca30c8546d306af7cdada8d2a8037200d303e6afbd5a4f448;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib8f9b76d6cf7a74f0d437f634ce888096a0d6d81d66dc6c60b62a60006b661e9;
reg     [1-1:0]          Id34d005cdd89bf304f95101c6fbfdd40d6c0b1742b5f3bee3bf043bf88c3d063;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie55394a5e3d49de60fbc4f33b3f9813b885da2049376036c935e8cd7c85010d7;
reg     [1-1:0]          I79d61ad4114817a49b1dc8e9314d9e3be9758d861974ead362ff0ac862d1d77f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6240db37d8e82731a264e5e3eeabb88e632dc6445647a26b4abdb142ff44c03;
reg     [1-1:0]          Icfe1fffea36cf64044389903be9550fe283d4dbb7f1b47aff2005e70765a6045;
reg [MAX_SUM_WDTH_LONG-1:0]                I4dfaddc409bf6d3698f255e55590182c2c8c067e0766311322460720dbd0967d;
reg     [1-1:0]          Ib08cf17b2065d04f587d1a8231ec1e4bbb6b2b15819de8a7efe18b477515ccf8;
reg [MAX_SUM_WDTH_LONG-1:0]                I1dd3e1e1e78d9e24a54fc937e7a25fc0e2514eabd1c1cc662d81ba73aa44680b;
reg     [1-1:0]          I21832b7270210e1bb6a23930ad9ced36d3da201d80310263e26eb96bebd23612;
reg [MAX_SUM_WDTH_LONG-1:0]                I80d4a0cc8b63f2ce0dcb344da5a47c95cc28b5f93d5bc6b77e9b875cdd58db99;
reg     [1-1:0]          I5dcc76c47f3c9129431152fa6f7047be203fc556198b45db15a9991647bb8c85;
reg [MAX_SUM_WDTH_LONG-1:0]                Iec19b0b63d20ea69dbcb23411a298bb6e833ee523fdf082f9343a695891a990f;
reg     [1-1:0]          I450f5b0f5d2b96636ae010048040ebd744fc4ca164cd764bb33615741ecaa62f;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib612f39370c6527c5f6eedb0eb5e7676212642673e940402586e823ddcbfb4c6;
reg     [1-1:0]          I35d64df6881fde0d4836aa408258db7cc1bfb2f066abf8c9345670b78c466b9e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifa501efa24e47050960fb3c383458a20f54abcbc5ca45bbe2d15a037670cd5cd;
reg     [1-1:0]          I11944fb91fa1b1d5f076cc36db77f0f8434f0edbb1236c7a9bcb45f79432ea9f;
reg [MAX_SUM_WDTH_LONG-1:0]                I8f088dd043a22011add21694f90df62fe1d2f6670cc72cfee805c9fb49756c77;
reg     [1-1:0]          I49642204473312df5a3bcab2692aa7558f44f21416226675a4ec10b0543cc5e9;
reg [MAX_SUM_WDTH_LONG-1:0]                Id86d515c6d081de87b9ed3c3521ab079e93ee082d8a0b396d44b3b70cac06b9b;
reg     [1-1:0]          I24e0d361a2679430549932a968d7cc25f980275fea5554e3453ed0a652d31caa;
reg [MAX_SUM_WDTH_LONG-1:0]                I4f94812066080b656de1a2807f5f669b2a81085bfc0470f9868bf5945856b451;
reg     [1-1:0]          I386015f8daacd2ac9cfed376d3418b56ac13f075a43dde939e4056c29565a926;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia92baf4463c96e210b460ea02d7775353edc6d475d7a315b594b9798cfd17900;
reg     [1-1:0]          I32832b039ae7e6f4b1e38cfdf680e5044e383b921a76189054511ebe5b8c0d7c;
reg [MAX_SUM_WDTH_LONG-1:0]                I9d4c230c86454c5c5f9ec98917ffc8d23fd19105ef93ba860ac2650bcf43ba4d;
reg     [1-1:0]          I09fff9b84a38f3d19685f9627d01a7183cf65d72110802f11e8da0e01194bf88;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia4a28d520896fadbeabee4130dcf862a9542852d87be480b1df2b67817f0ce65;
reg     [1-1:0]          Ib82c65f09934744abbba984b6e375bd69ce7231a5085bb00ba4e673cfd3aba38;
reg [MAX_SUM_WDTH_LONG-1:0]                Ide9498000905141bb106efc7e2184bd460d0e59a2270b10d42f981cf3bd514cb;
reg     [1-1:0]          I8ec5727130bf67c04580aa1b5b46cdf964db65750f2fc9ce55025b1c117b2bef;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie9a6b0e499ede3f80403e8f9c795ef4e93108ee8db755e12fb931259f1699712;
reg     [1-1:0]          I862dddc300df692e8bbf4ca45a24d840e51ac1e975631cf4ebb8337ceefc2eb1;
reg [MAX_SUM_WDTH_LONG-1:0]                I362132341c8e8a464a2bc93e7cc5b1d9d7804dd93965614dc340b48fad5c92da;
reg     [1-1:0]          Id08a37df0c5095196e2d760938c4d0b7e8716c25b55d9a9656d86c2c473f9c2f;
reg [MAX_SUM_WDTH_LONG-1:0]                I4b3c222863418745872c878545e419ee8f9c531f2cba89d28f0787992b0be8ed;
reg     [1-1:0]          I40204cd18eb803f82fc3ef933553c6ec41331f6d4a15538c287b8f57adebb89e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie39e570f1b5dd9f1ae893af78d81e458d077fcde2aeaba432209269b79785582;
reg     [1-1:0]          I677f733f4e801d99dc2fd1987683a7ac6c8609d84da6c95b8a7056ce07845665;
reg [MAX_SUM_WDTH_LONG-1:0]                I50ebc7f8f7cf324814b5885b2b18c90bf5007d8030744263d6e66880d836eea0;
reg     [1-1:0]          Ifeb10787a88bae5943b616e3bf751faff5e7eea80e45e24d60a760f4d6b0154c;
reg [MAX_SUM_WDTH_LONG-1:0]                I326b57b49d3fcfe654c4cb9ebcd6edc0ad7969e3b531f498e3c31270a5c4aa70;
reg     [1-1:0]          Iecc97eedc286cd1c3d301e35036e81a10d164d59da9252a92ca5f355a828367b;
reg [MAX_SUM_WDTH_LONG-1:0]                Id3898be2185f86831f58bd16651edee3d1bb21fa07b33a1928740ab496404178;
reg     [1-1:0]          Ia9a21e6f22a6cc828e041980ab142b418938a92bf8e868216402a46b8c614a19;
reg [MAX_SUM_WDTH_LONG-1:0]                I2aa77512781cba636ab96a5d09527e1ac34623ea2bb6c6a8d742bbcf6eff499a;
reg     [1-1:0]          I355f4f82732333ae56692d1c7ee89b368d938d9ce1d5f806be7e46482c10e19c;
reg [MAX_SUM_WDTH_LONG-1:0]                I225543794992ac9aa68ac3eeea38d41077ab5512b9f3b95fbd65a839294088e9;
reg     [1-1:0]          I9b2ce64b97ca55921bacb9b6aa4cdc8da5c1e33db4215a2470b7cfab3693576c;
reg [MAX_SUM_WDTH_LONG-1:0]                Idd1dac44a6f35d558d400160a087fe7628ef80ad72c3962df2b3a3809b89bcdd;
reg     [1-1:0]          I2d78ac4a4125ec25a02df6484c0ae640a37f915383b72f33b91e87cdf376fdf7;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic039114ea8ac4120b09973c79fdc044251fc66bdeb18a498dd6ed7265cdfba2a;
reg     [1-1:0]          Id727bdc545af53e8f89be0ac5627d0c0c0f0bd7d75030bcb41f198a4fe9c7d64;
reg [MAX_SUM_WDTH_LONG-1:0]                I21b3fa431ddc4bc8eacfb17a90fdac2bb32e4d0f4d0118715642c37601a1f883;
reg     [1-1:0]          I7661c17a1c73dbca82a6d3bfba2ab85ebb0131c1e513f093e1b0aec54907595d;
reg [MAX_SUM_WDTH_LONG-1:0]                I1c6d953c9a0e96d328cc4b515867b2ac21d2947a85e96be19f38e67a8b15001c;
reg     [1-1:0]          I553a83634252c50164bdde3576d7e1552a147490d02eac6dfd1140a46b813d08;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib823a58e9d4db87e4d73a81a772a02435af32a11d3c2265fb8a16021cfe4503d;
reg     [1-1:0]          Ib450c1ee41d04516060a410bbdfb605f0ce13cd8781596ce5218928ed207de8a;
reg [MAX_SUM_WDTH_LONG-1:0]                I3427390162b0952481e5f0728a20075c9cfb814431ecbb1a4014d407ab3b3afd;
reg     [1-1:0]          Ica745abd4de790f1cd3e2a5a32a9d0b5edf1b64e85759c49f3b4e51779443709;
reg [MAX_SUM_WDTH_LONG-1:0]                I35a9ae1cf23d8697091de65a1d0678632bd6889ae32408d7658e542a756e95ca;
reg     [1-1:0]          I6399b29558311ea40cda1388848ce13bb7593bfed01ca2a10fa5d8ed6700df56;
reg [MAX_SUM_WDTH_LONG-1:0]                I37e54e8ae28cf1a36cb9101d5afd4d523ca9a6ae244efe641c547a4114726bea;
reg     [1-1:0]          I6f529a4dd77f75d9af4350baf53ba61c1e9c5ea6227c26690987d244dfe71528;
reg [MAX_SUM_WDTH_LONG-1:0]                I9544a194d3d75c6c414169ea2536e111c09711ee602eb3462c4022350906a21e;
reg     [1-1:0]          I7a94e46f1351801c2edf76bf3b70e3b5100b8e6108d60d9341591aa59f4e95d1;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e4bc72a55efb8462410905dcb2c9a8412e2533ded854d23ca648e0e36802960;
reg     [1-1:0]          I0b761d71a88d70e6228dcf7325206f840d9da85892ba151c317e06079291fc2e;
reg [MAX_SUM_WDTH_LONG-1:0]                If2cec64e868d25d7fbad45ce4889c6a4cac0084aae00d2aa8963678edbb88875;
reg     [1-1:0]          Ic2ae521a3a6fef956f28a89da365b0838d535c9f7801a405cf60cc776ba0af2a;
reg [MAX_SUM_WDTH_LONG-1:0]                I73ad61911b0822e313aab2c484d1699cf2655a42a2bb0a1c9ab36228e41d0f7f;
reg     [1-1:0]          I01d9f8a8900be1981c601c0ccb45c1f39a0fdc16179245d80fbb2ad6d7060899;
reg [MAX_SUM_WDTH_LONG-1:0]                I218255d96e659dc8f60cddd40cac94a56d93556ed609b60157d88b298ec95f0c;
reg     [1-1:0]          Icdfc2f0ce24f01af7df8a99b58de3a74e1dda0eea5b41ff2c342106cb226abdc;
reg [MAX_SUM_WDTH_LONG-1:0]                I11284a18d6115421b4c76054c1a580c41987dec66caa7d5bd9107bbd4ac8bc2c;
reg     [1-1:0]          I929ef5474f10c76c4686fb044b2833b6ba1571f2e1c82b6d92cfaadfa44946e6;
reg [MAX_SUM_WDTH_LONG-1:0]                I8516ef195e4ba8f6e29a02ab5ea349a26bb68f6ebb4da847d56c03c942e9c20c;
reg     [1-1:0]          I55312932ff9d69c8ffa1e42efdb5e775ccb21a8f9e8791b080b67654462e537a;
reg [MAX_SUM_WDTH_LONG-1:0]                I2411dfbbf605c7590bc678373dd20b7241356a433756332f9a3445ba8dad57fb;
reg     [1-1:0]          Icbdbaf4eb2f30bb78db34a582e06dc91689b9eab2f8fdfe4fbfb41a8cce93ca5;
reg [MAX_SUM_WDTH_LONG-1:0]                I69d896cdb2303b99b73c4d6886f2686381230feca86c62fc064a85e4d11266f4;
reg     [1-1:0]          Ifa4cbbd5c3ab5e47a7d5135e4dbaf365e79c4c6a806bfae88c9c0e1c9ffe2fa5;
reg [MAX_SUM_WDTH_LONG-1:0]                If6ca882e537cdf5f458a2e11b7a11f057a3d2a00923825fe236afa0b0e1442c0;
reg     [1-1:0]          I2341907334935e19ef0e392216e39bb35c215730c464a85c0e1b804b364b492c;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie35443efbbf821e07284652a4b37347c4cfb959495dafa4fd2f81ffa2edc56db;
reg     [1-1:0]          Ic0bbaf8314688690b5a15a5613ab149f604a8bfb92a2b9ed014e7ce2757d0743;
reg [MAX_SUM_WDTH_LONG-1:0]                Id6d0b1fe00e5324e0ed7c37d41ee3e848f9c7dcfb4a85f5da2b82ed4d8942b21;
reg     [1-1:0]          I19ff0bebf62a994a2b5814ea41289f72cd62a38d2f37dc0027beb0f488926d4f;
reg [MAX_SUM_WDTH_LONG-1:0]                I0a309e8aa7f7e07abd837c99be6d8bb8c29dc1679b449111a02f49442d5cb432;
reg     [1-1:0]          I4f9435bbcce379d6d591547481382ab188003b97877c0f32462ef9e33aa8bc1a;
reg [MAX_SUM_WDTH_LONG-1:0]                I416c7ff28cd1d182ba2e08c3882c04d5073a014f7b9b41e56a3850cdc289ffb4;
reg     [1-1:0]          I9e497e3ee797c274b82ecca58218c47f9b663bcac21b1431b45c17d5e54e5a4a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie44d1a587dcdbb709546c6c567988fb0a19c276a1df7aced4c09a029196dfd4b;
reg     [1-1:0]          Ib929181cef39d751d2726a054cd0478d309e58350ecd11d3363ecba8bd4cb7fa;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic2b8d811fd01f5cd88dd60bb1b89b33163b3cbeae48d04e2316f15500c6a1a40;
reg     [1-1:0]          I64fa7f4fa09b7909840d8edb83f29f6a2379419e65b80f592b37d8ea00e59475;
reg [MAX_SUM_WDTH_LONG-1:0]                I85ff9ab4f9a4a3301bb8fcdc7107202263af0c37f091445efb5fa163a6b47a51;
reg     [1-1:0]          I35beac843abd6268c39acb691d3105a5c386f05461bca8c63b951ce1c2ed07bc;
reg [MAX_SUM_WDTH_LONG-1:0]                I39ab1bf4bdde9805c5bc7695c4700975d5a6094c40e107b82477192005d9ce21;
reg     [1-1:0]          I9d8fbde44d35c50f5f24ceae6f2e16ca2f280573caeb8a3021b6f69dec3d04b4;
reg [MAX_SUM_WDTH_LONG-1:0]                I602591ae56f1a42c64e50378841e065e79aee138622a0a571effe20cb48645a3;
reg     [1-1:0]          I507d851a78a765c18af6d529292384fb4cbb06cfec0e22d516adc79b8ea13c7f;
reg [MAX_SUM_WDTH_LONG-1:0]                If37e9ed3af8a31c989dc6ad554207cd464c591b630ca1e5cf56b2eca57a18d8c;
reg     [1-1:0]          I80fb8d450dd144ffade989cc2cec363cf6bbcdc267f5372163fde38313387499;
reg [MAX_SUM_WDTH_LONG-1:0]                I80099c7b01770cc5f7edb3a3551d8edfe9dccbcd2a12daf8ebbafdfccd141bd4;
reg     [1-1:0]          I7844074cddcce1b95a010729a9e4ce2bfc4f7e1962b84af0e0a3cbb2c2c08206;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie479ccbabaa8a00009152557e4de08bd240fd28f1b131c674dafbcc2505711f7;
reg     [1-1:0]          I88be0c0499713ce396832a79853e9918ecdfed2519fba6fd7c0bae51450478e7;
reg [MAX_SUM_WDTH_LONG-1:0]                I6364406b04427fe3a4cecbed48e12a67cb08dc632b2914b0fe52fab0ca541c0d;
reg     [1-1:0]          Ib585733bf4c3eb59a772866965420fc7397b01272410cdb701f289daf9549fc9;
reg [MAX_SUM_WDTH_LONG-1:0]                I610dd39f1d44d84764b0acd6b3fb1219fb6b6d6ca92e1b226ca76a389bf6c937;
reg     [1-1:0]          Ida673298c761bab46fb26d4e73caa99f5b3ade7f924d99fcedae4e47c70b5b67;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib9f9384ac4ec4bad29fbb4ce683ffda7dcab311135f02b6336e6209f5742fddd;
reg     [1-1:0]          I60bb81cc7cd9a6212f7b4261a21655accd6cd09e7aaf5f78f7f1f4dec0e8489b;
reg [MAX_SUM_WDTH_LONG-1:0]                I60980f76d468775bcc8a7052681fbb6ef4b2243e5e30e5365cda6cf598bd0bde;
reg     [1-1:0]          I85d3c885ce504524ab43daed7bbcb599cd7e5d6d3635cf46e278345134e97e22;
reg [MAX_SUM_WDTH_LONG-1:0]                I892a754f0322d92126d4731e8066760a24897f93e2afb858ee1393604d2cbb26;
reg     [1-1:0]          Iaa08a49e0ca4f92f38c7f4d115ae1b275e45c42dfa6fd4b6a2ff40536b7f5f15;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib0f8816eafd3b950f67cfbdb6a44c59ab7c0918979817a4a998d8305da847e72;
reg     [1-1:0]          I197b3231cb1da107c5001075809e9fa75e4089871d473490981a8b44d3ff5e4c;
reg [MAX_SUM_WDTH_LONG-1:0]                I04b55f2c45002f1f1f7a6176773a22730dcfea14662f0badb102ddb60b84cf9d;
reg     [1-1:0]          I384c04b75344f97c691f70965d7e08266ab9cd8862e04ba73b502a0f36ac5ea7;
reg [MAX_SUM_WDTH_LONG-1:0]                I5edc072d158ac583bd1cdb2449086d4f0b17e36d724f4cfde79820788ce57f31;
reg     [1-1:0]          Ibf95afb3941a2272d76cd7256d0789f11fb35a3020c3ccca5b099d335d4a2330;
reg [MAX_SUM_WDTH_LONG-1:0]                Ieb128919ed64e331affb6adba798c267e8c3ec924a7ef58f50b1bc0b29702c23;
reg     [1-1:0]          I885622bb1c7371f4afa3e9966f870d2bf7750c2d2280a2a993a5bd9854187994;
reg [MAX_SUM_WDTH_LONG-1:0]                I90cc372cc2f3b23eaaf2cb32da95ee715af64ca2eaee77195d9813647d2a0d08;
reg     [1-1:0]          I719a3e78d6a298f7db920bf7e355f6fca2c46135abb8ccd1cc3ea470912d05c1;
reg [MAX_SUM_WDTH_LONG-1:0]                Idaf65411d995039ea730b6ee4b5ae727325da17dc79c8664270d60f063828453;
reg     [1-1:0]          I1729b841d155c32b617727459f01aa9a9a6af56de5f464e20e900e3a4da30dba;
reg [MAX_SUM_WDTH_LONG-1:0]                I977557441002c273f9b9b8748ffa9edceadb342e028ceb581c3bbce9af103a74;
reg     [1-1:0]          I96affe6d042e09b07278ae45744977fd3719a31fa5d578adaa2b3a66b2c3ebd0;
reg [MAX_SUM_WDTH_LONG-1:0]                Icc10ac19a64065f5923ecef4f1353f13c7796c23f2555f8ae6566eb538d77677;
reg     [1-1:0]          I12e1e01b28d2d443785fac1d0314b477b221b17b715f1153c5379a85b4b5e3aa;
reg [MAX_SUM_WDTH_LONG-1:0]                I725c369a5013eeb6b581209bc8a921fccfcf1754137191e26757abdb72ced94b;
reg     [1-1:0]          Ie244ea5cb57e0b4c14c0c8c22592347d1389a6b0f53b821335b821ca5130ad6e;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaa02b7ddfffcecb763aa916a2bc4c3aea58027c89b515c40b72214d9dd44ba21;
reg     [1-1:0]          I5a07f349b1fd7d668d35583c50dfa3ceda070e5dc241bff1ecdddace6624bd57;
reg [MAX_SUM_WDTH_LONG-1:0]                If8737fa82b71d9b0e7223baabca7405e148621600bdaef02e65cd7bd175b2d88;
reg     [1-1:0]          I6e5f194e3acb27a7fdd060e05aff00bb9fcd0904b3f920d7db0fee84c1534558;
reg [MAX_SUM_WDTH_LONG-1:0]                Id85c2b905d61bcdc87d500d6ede3ca02d52bc3eaf278f087f27fe6f277c91262;
reg     [1-1:0]          I09780397509ca78f4b4aed5b08cf22d8eae797d1d1864cdba4a951ac8d583c91;
reg [MAX_SUM_WDTH_LONG-1:0]                I5923f41aa444bebfc18d13202747ff84e20a4753bc9cedf697b9ae8ec3418afa;
reg     [1-1:0]          Iefcb9b5b2f238005d0f37bc519349bbbc130e3e072814ec48b4edf9c853a6913;
reg [MAX_SUM_WDTH_LONG-1:0]                I4ac498dc826a9dbeaddf2f013ae7116e92dc772ea55987a4661f18e56a4123a8;
reg     [1-1:0]          I9835f6f38580d8765566723f5a9adbfb4935af8bf719b3e4918e1b746cf12241;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaadbb1b235a85c555a6f37d003e87a987b7d9b07148207555eb717b7332f67ec;
reg     [1-1:0]          I2266ca44e019a30bb553f955a158a5b075035c4b20a0b3fca6a3675ec79b9997;
reg [MAX_SUM_WDTH_LONG-1:0]                I6afb533ec993de4f9b04007b355a9cadf08488ee6ca02aec2d7916a4c98a7fad;
reg     [1-1:0]          I684ec077e37638f022f10b5eb31403e6f9117a83a606f2a5013c2c33b8d1a8ab;
reg [MAX_SUM_WDTH_LONG-1:0]                I01313177417c899543a67763ede925dea3ee58ef4a31714ad15a7a3746bb5be5;
reg     [1-1:0]          I9331428911b817ea45d1b5ae75eb3ee6e05c189785c995e5d2625f12ce4e0846;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibd0ba147d1a08acea707b8c60da14ebcc4ad62e67ef26634777b5dae38af6d61;
reg     [1-1:0]          I7769e8ceb72790c37b351c32983860280aef172974d19a2e99348607863a97d4;
reg [MAX_SUM_WDTH_LONG-1:0]                I1e92e18a915678cc96aa493a00627dffecbd341dc8e022615610061e52c1ac3f;
reg     [1-1:0]          If09c36408407b246848b29df63e789fd1041815243beb4f27db0e774e853f1cd;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia7b91fa4a1ef16f859ee162b91daedc97927244dc19aaedede898049daf85a19;
reg     [1-1:0]          I533b63eedc528cb36abc0a469b66b144a6ae5122c038eef85d8d0557c3dff3ea;
reg [MAX_SUM_WDTH_LONG-1:0]                I9918d91748722a47f8526008bc3fd4c498bc80205211d5c92acbc511fdb667bf;
reg     [1-1:0]          I051e3b709db2e7861d31165ec1e5ee679f1e6dffa5a951072831ce479c16f27f;
reg [MAX_SUM_WDTH_LONG-1:0]                I95d109e37a87827de1455b5ec479dda78a0218cb9db245b80710cdb1e8ead67a;
reg     [1-1:0]          I2fa018ce903921d0a174a63dbbb29eea8d5700b376335b2ba9bd448e8782018a;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia0c7162290e415f24699688e45850c243397b5cccf07daf0398dda04810b0690;
reg     [1-1:0]          I36e06c1d77080ff75778f3dfa4ed60e66f9a3bedc39b214e3fdb5b6c21f1cd3e;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib9dc17b2b9fc7c228eba40cf625a49a27ec16f8c8a91957de14fb6849ea49212;
reg     [1-1:0]          Id647e3bd88fdc7a3642092d071f66f74657c8364937caf63c723f1e027c157bc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ied32ced79448b3f92faf0dca1673559e07372ec338e8c51a750be1c6975a298e;
reg     [1-1:0]          I015b73e7e4bc4c2a3073a304e58d24f5c8c32e90299f004bc0f75eb9e18e6d41;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaddb000276bde734c13ec1395f06c1b3bf5606ad5cb138579d711cecf26ac88a;
reg     [1-1:0]          I7c211cef6a581c5a6871d4c9a2b7ba29a9d05d36b0a758106e006caebfc592e5;
reg [MAX_SUM_WDTH_LONG-1:0]                I211ada7f9095ced6b3d20f8f7f67b56cd2e73595481ed5d4c08175ca874d16ae;
reg     [1-1:0]          I3f2014435aac47a3c807e9ad3f0829179f9285582b7ff2e3bae250a25e800aee;
reg [MAX_SUM_WDTH_LONG-1:0]                I0d49182fe7486bcf54c8f68904b4b90436de6f3bc42fab67a4e47f61154e22c4;
reg     [1-1:0]          Ib27fb4891a6edd486a99f23a750057de12a5a3e3fc6a5fad7976aa7e961e0c54;
reg [MAX_SUM_WDTH_LONG-1:0]                If79b91295d25c503f6bf5ca7c6eebd2ebf6807dd9990ce31e844cee0d8f89dac;
reg     [1-1:0]          Ib58cd067e009a5f4b72af8cfb1e5c49c18f51a2ad8880f65aee683bf8ecd40ad;
reg [MAX_SUM_WDTH_LONG-1:0]                Iec1d04d20ec09595743b7a35860b5cb2ec862c20da87c6f899284069c60bdd71;
reg     [1-1:0]          I7e40bd6625b1d7deff82f67d46817c7af70f1da57561ab528b553b3d244b3f1d;
reg [MAX_SUM_WDTH_LONG-1:0]                I2126b1597a95d7aeb7d20d4e0f4270e1fc5cb0fe6eb5003b05abbb7e5e9a2819;
reg     [1-1:0]          I01949f24f74578cb63dd095e8ce639ce0d273c14da81e75d00097535e391aa4c;
reg [MAX_SUM_WDTH_LONG-1:0]                I72a115d9b3659f31366e1d73d6d9a0793e20be233c3ccab2b513fd79786224bb;
reg     [1-1:0]          Id8f2a0d3524b27621ca5a576bf16e15789e6257060225da04da2a5fcc8cf751e;
reg [MAX_SUM_WDTH_LONG-1:0]                I469b0bcfe9cfc27a8596782bab479f30aedaa132a5cd404feb1fec4b52a17d3a;
reg     [1-1:0]          I6020dcffd9e047c03740cffcdfe790eaf614ea1036a50fefcec9e13e5b5ac4bc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib4c52550766a2cbe0de236d6783edfb1a6a7cb4c2bb9333a9379e1b75680dad1;
reg     [1-1:0]          I815f772d86db329f78fa75c3326c129ccf0f6c5f383b42ef18033e48d11525d2;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaa72101e8c3e7fa248ac4d4336b3847c4f602b6db009e9cd74cdd25251d5178e;
reg     [1-1:0]          I2c8a33831a21c4c21dd58a300467abcc82d52e7636a73a12a003a4144d43e0dc;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic1381219782d18c1cb880970c062eb260d9d3be0b597e1465fc604c0c0c32c68;
reg     [1-1:0]          I8c7b9ead4ab28ae2c2aa5185a0746c9cfe9fd90bdd68f2ba05291045a296d566;
reg [MAX_SUM_WDTH_LONG-1:0]                Icf0c3c82c9e458a347212415d3029f192c40152e8525a20b5c9bfed88ccdb32e;
reg     [1-1:0]          I32ed4ecd4363760151c1accda085c9afa3efe63daf7a312feefc00b804401c27;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic5a87abf4c6018e9555de321c141d9754a7de91f1743d980e339ff9cebd63b7a;
reg     [1-1:0]          I6aa6d6c6213348ea0cc3e8b207bca2c1db81499441e4ed721ca0ee01ae831291;
reg [MAX_SUM_WDTH_LONG-1:0]                I3a27e4e3322c28e7fe85d7e76b7d5477f4d4f6acb8cdb876b9a54cba98b189b9;
reg     [1-1:0]          Ib4f23d2e5f8c73110ae24212c4ec0e7ef29c09c8178ec3850f061a5b0386feca;
reg [MAX_SUM_WDTH_LONG-1:0]                I11edfeb948852dab396975b53b12d09da7a5fbedc2dae9fe7c687768cfef05b4;
reg     [1-1:0]          If2be986b27ce8aa2117f87e9a144015a10acf0a07847f83acec2804b9e987e8b;
reg [MAX_SUM_WDTH_LONG-1:0]                I578437932d2d1156445b41a1238e0fd96ab5702bc3158ea337a9e37d14d6731e;
reg     [1-1:0]          I9f17331c6a9858b60705d889b5b77078042cffe9e956de20eb067ad7e70626b7;
reg [MAX_SUM_WDTH_LONG-1:0]                I3c2c5b5cd798851c7fcb0d0e66ddf81a516ef9bdf4aa4ebd4901532bfb2a651b;
reg     [1-1:0]          I2b70416e96231188e62b7bcf0300c4a5b2d2139449150d31414b92ae075aa0e7;
reg [MAX_SUM_WDTH_LONG-1:0]                I8153d6f17d832da24daaba2909a88f1609e523ad3b6eac7ad42521979aae96da;
reg     [1-1:0]          I29599a1dac362c87f4780a94478787a718f63401d2051ccbfe543b44e49b35bb;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic10ea001dcd0b864b987bc3080e95b338c1e91247bb90e884e161c926183fd2b;
reg     [1-1:0]          I5ff7defb023005e77164f9f3b852fa60ce897922c6b814015d3436fe1d1b4a44;
reg [MAX_SUM_WDTH_LONG-1:0]                I61efe7187a1aaa28235dacf68eb1e1dd97e7cb5900862790bb4d5872d7adbd67;
reg     [1-1:0]          Ie132a24e667376de85b8fff9a639698df164043422122a8058c968bb7996d3a7;
reg [MAX_SUM_WDTH_LONG-1:0]                I3c710fbd5e4dce0c97eb9da2d8e526f9d44d87fa75088c0421353614e6ef5da9;
reg     [1-1:0]          Ie8d5dfc9a77dc01055a551c5f37416d0b13ef83428bf751fb9f95c7d10442697;
reg [MAX_SUM_WDTH_LONG-1:0]                Ie02f677979058dda2291ddb93acd64f4461f6d75f3a33c21dac97129344f7055;
reg     [1-1:0]          Ic94f2b10208cb23bb5f5b1a46c11c3bbae038308b385373cfaad9a18e09ccb90;
reg [MAX_SUM_WDTH_LONG-1:0]                I2b78100b50f7334d563daa27cab8078fa374dca0c438157d1ad44ed3fd9e3456;
reg     [1-1:0]          I3b79a6c69be124aeea9d1444f9f985201b55ad0d7a4767a01f612eee12a6ad73;
reg [MAX_SUM_WDTH_LONG-1:0]                Icdfa68bdad11213dbaa576cbf43ca9deeb1f9f24225264eaeeede7d1aba5fd8a;
reg     [1-1:0]          Id3ac4bf805d3981ac1eb1b396b3da5c0dbc68754d89668f0a4cf7c6f2a44ddfa;
reg [MAX_SUM_WDTH_LONG-1:0]                Idb39db95234cbfdbbc89fdee230784c703e170b9e932643a5e1b811b24ae021a;
reg     [1-1:0]          Id77fd99c6146776bfc20804c67ae41b88cb0441eecba4f40b87828956b7158b6;
reg [MAX_SUM_WDTH_LONG-1:0]                I7141b42fce475b5502fd33035bf37addde06271b2259e158ba03a66843b66075;
reg     [1-1:0]          I650a7220fd4eb743f652c6c1f9431191621f9fb1a5b5d64bb9649b43bad5b8bf;
reg [MAX_SUM_WDTH_LONG-1:0]                I245e922da0aa5470370db389d5bc9db33327c905528a1740aa015b7ccdfcc29e;
reg     [1-1:0]          Ib7417e90e9dc35367f110c364878657dbbf66b1a714d5807e6347095b833c62d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia2ff4d61c4f4fdf29be87b50e206c308cf970cbad2638e86ba8c2be8d025b534;
reg     [1-1:0]          Ie59a4afbd0d65de2149e8c60229bce12b77f8f1b2b232a11fb9714371eced2b9;
reg [MAX_SUM_WDTH_LONG-1:0]                Idd383630385363471e1b17ea946a61194a3cb287d833af386876c3b4ee66e406;
reg     [1-1:0]          Iad3f7ae48f752d3ee71320875a2d1d170e879dd5ff51cdfd662241e6a30fca6d;
reg [MAX_SUM_WDTH_LONG-1:0]                I3daa8702e9dbd047a05e5ea044d14b670c2ae3849526cc514be6a511c5c45c35;
reg     [1-1:0]          I4e9c85ad6975994daf65df213a2d2fa5a6a2abd91e66d9c9a6f540caf4c2afe2;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia695c63ae87e9a6742c6fecea648a214f5b24ea2b652bb5d83f35d9a59b94f72;
reg     [1-1:0]          Ic8f9966a2711f4810086d09b86e16ccf0d31339d146ad5c38d34c973c757947d;
reg [MAX_SUM_WDTH_LONG-1:0]                Ifc31b600cbbf26e78cee82cd354c17b872586c1a53ddd132edbd25ce87d8aa9a;
reg     [1-1:0]          Ic1385b7aee4e3b643e13733b56157e3e92e638da28cd1234e275fc9263709f04;
reg [MAX_SUM_WDTH_LONG-1:0]                I261e70e693cdbc572e40e81c594f3dac624febb03465bfd0fb864d337e753499;
reg     [1-1:0]          I3a173e6b224a6415ad442ae28a0af62756975427859bbcfc0af6c8e5effd62a6;
reg [MAX_SUM_WDTH_LONG-1:0]                Ia6f7ae0adde8136c7a25f4fed69bbcaa376b5f28cbb4990afabb57a87ec03019;
reg     [1-1:0]          Ia5580120af4590da8aed890f81ca17929e4c998617df957686c095e891649c83;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic40e94217a2d2c13f4b1ad2766ab1ae4e8ded0b5e0a3522dd51ec806c3e9feef;
reg     [1-1:0]          I58a3910d475757bccbde2da0e6b5dd5723cbe44e1f4d3e71ac2973fd2a03b3a8;
reg [MAX_SUM_WDTH_LONG-1:0]                I78602c68a4a00f530bda7ba1dfa4820b7faeb0edabc636d6a2d8bf97005755d1;
reg     [1-1:0]          I1b76b0f61e714e21a844e429806d641f6a24f0eb19c23a3c2fcfb76baaf3e72a;
reg [MAX_SUM_WDTH_LONG-1:0]                Id8e684d92e6d0b6e10b5e7f7ff9656e6fc67c99edaa59b49e453844ae33d23f6;
reg     [1-1:0]          If0211848e6cda136970069df5b6156d4ac213717491c68ed49ab39d2cffe9999;
reg [MAX_SUM_WDTH_LONG-1:0]                Ic9d9001a209401fca8a3f28e39c4b89adc8f4e9d225aeffbb5d30893bea1a7b2;
reg     [1-1:0]          Id23ae21f713f4f452abcb1c1839b5524c452bb8bb0b6c35683f9bde212bc5f96;
reg [MAX_SUM_WDTH_LONG-1:0]                I97f666707f6afacfc6156ef498941fe5feeb7424834b4a283139aefb5f50a68f;
reg     [1-1:0]          Id5bdb0f5a920710b1af7cc3abade245196df9d1ab4b7f26277fd93e1bbee5556;
reg [MAX_SUM_WDTH_LONG-1:0]                Ibdaeb96b71f9ccccfe79b1b3bab77122aa32217b58037d80a3183bf888b60c72;
reg     [1-1:0]          Ic72616171e7fb8489fa12cc29be1f74602ff8e4bd28ea085e938da615238a0fa;
reg [MAX_SUM_WDTH_LONG-1:0]                I574e4843ab81be7ad95cb7027fc3284a8780b07fb8a194a9c991997988d7ff8f;
reg     [1-1:0]          Ia09db6bd7cba6c6e15cac4c6ad0d4c98235a7437beeabca1388fb1b4dece5d67;
reg [MAX_SUM_WDTH_LONG-1:0]                Iaa4463f258ed92a2c85fef0790c47e725c555f37c80dbe366d973c9599a5484d;
reg     [1-1:0]          I15ab76f6e4824af9b3b4f5062e8dd3c426e1ff0c5f68e4733828c710eb7bca54;
reg [MAX_SUM_WDTH_LONG-1:0]                I7102386e760e34e2d0fc4563b497acec7222bd171333a2169fac800df94ea27c;
reg     [1-1:0]          I12b276cd6b0aa86ca2e28dbb1f4008ab140668e16e4ef96604a6d1741c7f2f95;
reg [MAX_SUM_WDTH_LONG-1:0]                Iee34d958bf4feec1e5bde8a866a9919f29edd54f1bc51cc9c8216b71101d640b;
reg     [1-1:0]          I01577c8c0e65ca47449450a8b2455ee84cf5c48bb26a0799b5523258a039ae40;
reg [MAX_SUM_WDTH_LONG-1:0]                I64b0ef6642050de0690c95be2af9606797be36c1656f1306b87ce3e8131c4629;
reg     [1-1:0]          I63ba87cd2daa7c3c625d3ff5bdaca7f2115fc2d65e13972a22b2c2ae5b746d4a;
reg [MAX_SUM_WDTH_LONG-1:0]                I23f31ebee34c7f4f9c46fba41d41df176a7465c074ad8527205a5782edab6524;
reg     [1-1:0]          I576afeb6020cc0a8e35837b4b96968ed04cd444999558626adac849848fe7c6c;
reg [MAX_SUM_WDTH_LONG-1:0]                I628b9674d7d6caaa70c54539241df2e7a4be0441dde1739b442513c6e4ded8a4;
reg     [1-1:0]          I3b8769ce28405c0bb978c458bd6272f10cea5338af4170ce4e93a8932ae8dcaf;
reg [MAX_SUM_WDTH_LONG-1:0]                Ib066c9d790586949b27c4cf09dc957e7d28161ab00e8dc6920e4e0cc5ac665d9;
reg     [1-1:0]          Ib4638612fcabc0a2c2f2bba5a2b9eb71cdea23575641b3f81fb6220fcaf284f4;
reg [MAX_SUM_WDTH_LONG-1:0]                I57419941b1979cd06c4fa0e6be943f004dd80da502425ee5b6dabd2239139cd7;
reg     [1-1:0]          I16ea389c88e4591f7686eae3f1988dd5361bf893895697c0ade8627986a9fc5e;
reg [MAX_SUM_WDTH_LONG-1:0]                Iabb5703a54942b1bdcfe2213d2011c659ec812f751dc75943b2ce511c81ffaf9;
reg     [1-1:0]          Ia17edf214ab782c25bbab97f6bb4e04b2fc46d41f9a97fcf617418d54ab76a7e;
reg [MAX_SUM_WDTH_LONG-1:0]                I798a6a6074b50fc61bd4e1b4696560abd2e515c86d47f85e9a3077cf6672acc8;
reg     [1-1:0]          Ibcfba9f1fb81d976955a1fa7101f0b0db16c344c82cc5ce81f50dd3aa2928d37;
reg [MAX_SUM_WDTH_LONG-1:0]                I3f4a8ec7c554b1f0b9d3d2963b0e3dec4654bf07c5b836f8fd07c639cd19d588;

/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [22-1:0] [MAX_SUM_WDTH_LONG:0]      I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe;
reg  [22-1:0] [MAX_SUM_WDTH_LONG:0]      I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [22-1:0] [MAX_SUM_WDTH_LONG:0]      I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd;
reg  [22-1:0] [MAX_SUM_WDTH_LONG:0]      Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [22-1:0] [MAX_SUM_WDTH_LONG:0]      I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86;
reg  [22-1:0] [MAX_SUM_WDTH_LONG:0]      I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [22-1:0] [MAX_SUM_WDTH_LONG:0]      Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b;
reg  [22-1:0] [MAX_SUM_WDTH_LONG:0]      I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [23-1:0] [MAX_SUM_WDTH_LONG:0]      Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d;
reg  [23-1:0] [MAX_SUM_WDTH_LONG:0]      I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [23-1:0] [MAX_SUM_WDTH_LONG:0]      I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5;
reg  [23-1:0] [MAX_SUM_WDTH_LONG:0]      I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [23-1:0] [MAX_SUM_WDTH_LONG:0]      I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308;
reg  [23-1:0] [MAX_SUM_WDTH_LONG:0]      I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [23-1:0] [MAX_SUM_WDTH_LONG:0]      I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e;
reg  [23-1:0] [MAX_SUM_WDTH_LONG:0]      Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [10-1:0] [MAX_SUM_WDTH_LONG:0]      Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba;
reg  [10-1:0] [MAX_SUM_WDTH_LONG:0]      I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [10-1:0] [MAX_SUM_WDTH_LONG:0]      I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24;
reg  [10-1:0] [MAX_SUM_WDTH_LONG:0]      I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [10-1:0] [MAX_SUM_WDTH_LONG:0]      Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43;
reg  [10-1:0] [MAX_SUM_WDTH_LONG:0]      I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [10-1:0] [MAX_SUM_WDTH_LONG:0]      Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78;
reg  [10-1:0] [MAX_SUM_WDTH_LONG:0]      I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [5-1:0] [MAX_SUM_WDTH_LONG:0]      Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e;
reg  [5-1:0] [MAX_SUM_WDTH_LONG:0]      I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [14-1:0] [MAX_SUM_WDTH_LONG:0]      I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248;
reg  [14-1:0] [MAX_SUM_WDTH_LONG:0]      I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [14-1:0] [MAX_SUM_WDTH_LONG:0]      Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091;
reg  [14-1:0] [MAX_SUM_WDTH_LONG:0]      I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [14-1:0] [MAX_SUM_WDTH_LONG:0]      I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129;
reg  [14-1:0] [MAX_SUM_WDTH_LONG:0]      I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [14-1:0] [MAX_SUM_WDTH_LONG:0]      I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b;
reg  [14-1:0] [MAX_SUM_WDTH_LONG:0]      I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [7-1:0] [MAX_SUM_WDTH_LONG:0]      I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64;
reg  [7-1:0] [MAX_SUM_WDTH_LONG:0]      I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [7-1:0] [MAX_SUM_WDTH_LONG:0]      I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4;
reg  [7-1:0] [MAX_SUM_WDTH_LONG:0]      I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [7-1:0] [MAX_SUM_WDTH_LONG:0]      Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed;
reg  [7-1:0] [MAX_SUM_WDTH_LONG:0]      Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [7-1:0] [MAX_SUM_WDTH_LONG:0]      Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25;
reg  [7-1:0] [MAX_SUM_WDTH_LONG:0]      I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [13-1:0] [MAX_SUM_WDTH_LONG:0]      Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41;
reg  [13-1:0] [MAX_SUM_WDTH_LONG:0]      Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [13-1:0] [MAX_SUM_WDTH_LONG:0]      Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88;
reg  [13-1:0] [MAX_SUM_WDTH_LONG:0]      Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [13-1:0] [MAX_SUM_WDTH_LONG:0]      Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41;
reg  [13-1:0] [MAX_SUM_WDTH_LONG:0]      Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [13-1:0] [MAX_SUM_WDTH_LONG:0]      I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b;
reg  [13-1:0] [MAX_SUM_WDTH_LONG:0]      I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [6-1:0] [MAX_SUM_WDTH_LONG:0]      Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b;
reg  [6-1:0] [MAX_SUM_WDTH_LONG:0]      I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [6-1:0] [MAX_SUM_WDTH_LONG:0]      I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2;
reg  [6-1:0] [MAX_SUM_WDTH_LONG:0]      Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [6-1:0] [MAX_SUM_WDTH_LONG:0]      Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52;
reg  [6-1:0] [MAX_SUM_WDTH_LONG:0]      I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [6-1:0] [MAX_SUM_WDTH_LONG:0]      I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726;
reg  [6-1:0] [MAX_SUM_WDTH_LONG:0]      I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [8-1:0] [MAX_SUM_WDTH_LONG:0]      I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e;
reg  [8-1:0] [MAX_SUM_WDTH_LONG:0]      I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [8-1:0] [MAX_SUM_WDTH_LONG:0]      If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e;
reg  [8-1:0] [MAX_SUM_WDTH_LONG:0]      I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [8-1:0] [MAX_SUM_WDTH_LONG:0]      I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340;
reg  [8-1:0] [MAX_SUM_WDTH_LONG:0]      I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [8-1:0] [MAX_SUM_WDTH_LONG:0]      I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc;
reg  [8-1:0] [MAX_SUM_WDTH_LONG:0]      I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [16-1:0] [MAX_SUM_WDTH_LONG:0]      I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5;
reg  [16-1:0] [MAX_SUM_WDTH_LONG:0]      Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [16-1:0] [MAX_SUM_WDTH_LONG:0]      I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6;
reg  [16-1:0] [MAX_SUM_WDTH_LONG:0]      Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [16-1:0] [MAX_SUM_WDTH_LONG:0]      Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0;
reg  [16-1:0] [MAX_SUM_WDTH_LONG:0]      Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [16-1:0] [MAX_SUM_WDTH_LONG:0]      Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a;
reg  [16-1:0] [MAX_SUM_WDTH_LONG:0]      I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [9-1:0] [MAX_SUM_WDTH_LONG:0]      Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8;
reg  [9-1:0] [MAX_SUM_WDTH_LONG:0]      Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [12-1:0] [MAX_SUM_WDTH_LONG:0]      I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8;
reg  [12-1:0] [MAX_SUM_WDTH_LONG:0]      I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [12-1:0] [MAX_SUM_WDTH_LONG:0]      Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f;
reg  [12-1:0] [MAX_SUM_WDTH_LONG:0]      I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [12-1:0] [MAX_SUM_WDTH_LONG:0]      Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7;
reg  [12-1:0] [MAX_SUM_WDTH_LONG:0]      I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [12-1:0] [MAX_SUM_WDTH_LONG:0]      I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69;
reg  [12-1:0] [MAX_SUM_WDTH_LONG:0]      I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ida88a2dbb8109dff5f061f3ecaf9586a219f6355e92312ffd580a09126c72376;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9aea0703810e5cd52352d3b0ede17aa0ccb943f1e0507585e4cccd0d0c427e98;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I73f2fe34b7ee9a375ae43b6d3cbd515175de303a77f64ad277094e9bb8e45177;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I42c6c1d7cfb81335f01807b1d1c6b77c109482d338e81eda1ed174f739a6bf1b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9f9254e3af43fc1c116a2d33bee39fb18594b7696e59d5aa4c3884363616a5d6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I839de42c6f3369ef5c6200c12baee8c9e698b3108fd6dcd58a71351d9bedae54;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Idbd45e6a4aa2cf66d740fb7d3c41c5d4af78bdfe13d321e6ee7eceb153e03de4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0a1e88a592eeec68c060dd84ca2d75809b8fd80dd97a01a8d12cd9869bf94532;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie3a6f677abff075b84cd72fb72f4b4ad16dc2a915b2d3e06d8136c5073549499;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9114e17d37b4346674c23a6ef3a2aee35426292fbf73d7f30c895090bb749034;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6444b0cde8c0fcb1cc0b51c11d3937bd156b26f21a0eca3cabe0c6b0e696f7c0;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ife5225eb20e50e3cc959d9080f6faa318b4977bc9d04a67414a6cdf16c98e295;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1d41ad001c01e3dc84cd02ab5ba24e8239e273f81dad37de1fdf873305e073c3;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I28dfde2c443cd84194231fc87b8a1c6382ff3c2ff9b6d43e31e3a7116be41169;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I75cef0e0547fa056ba6e20b68cadef6bea875e9b12fe99c286e8d79a40c9043f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I55da00c15261d3abb33c69ecc3f2090fb2bb3c29a3653fd999f6232982cf31ac;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie4bd6fa32fac971db980d5dae63887ea1f4b75f375f1953975e4ead5b727d37a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I05ca033870ef7adc8ce911a962bbd120591a1fe3b3044782b7e569e2b94ac629;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I40f5e53051d38a2da1e0c992989c7740e6a7be23273e1412d01e853851b97a0b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4ef4ed6e15f48f289815b7e00b2454a26e076b8dc9b8903e118507c9688e905d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0e9c027df8259f9e499658f9ee700b50ea04b829312da04e92f13edd2af302ad;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I25e57b538f9a08a355a5ff8d26d94f81bbf2ebd0039881e74aec76ffb1dd48aa;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If5d8bf4cfab249bae208cb278b5fc90873cebd7a677b1d1e22df49b576863146;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I070ee6bd21603d58d3243ac556db2ca3c0476c64fde6d32aff54e0577b0472f0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I03501709a4343537388784e4e39cb9c1b52beb3749d09e2daaf1910dc5b1e2b2;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id2ede5f3d3ce0652bc9ceeadf1de91fb99234718893eea8cc1779cf900284e88;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I46aa1767826fecc6fede490a807238d69235f3cdf96dc753215e008a12454119;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie251294e2cb883a913e91485cecfa90bbd107955ceb6d60d4a9b1808aaadb2d4;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id749da645d127d8ff383558a6e7ab4a5c2a59f513cb7808fa4dc4e9f6f14f2b9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I983e8c64c323025590663edf53b0666d93d838f15879b5e3df245a8e9ac6fb80;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib15e62b641f64f20a1d3baff39f2dc6a403616e09955f5d7f47ba4fc093badc9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I46e5ca785f6f4304dbc4fbbf3816d83106047f0eceea77717a1ad5c41a9ca441;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I603d7bbab10dd31f19047e4a73046c804506ba70d1504351984be41bae1d180e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ibefeb67be2754ad6b9a6cda09c66529a7ca51536f5c6ca6b05e6ac1de34ae514;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia7b80ae8cf2697315846253262614611c079c53ada59bf7d982596ff8df770b6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0dd45b65c82498edff9ac44b5b07ed30818dc1ea2af48e5c1394466865f36adf;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I58250efea716c203d1475c4046ca67a47a156f9e4709d26d4b05a29ed1578337;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ica92be8c7303e09b9f549ec558e655816c1d23a39b8d5324060f64a391984c1b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I50cccb280c7d65372645e94b4a4d472860f246a8a6d89c02e4feee7dac903e8e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I726b6a7ed2ab76b049762263a08d5121a597f30ce25a6880b51d6b01aff801d7;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I01d4a1a1123a68c80a967604072ca420c79d4e205c354221591cdbcaa24c4050;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I89362accf0644c192f06b113020d2071f1389e8ddd8d4fee492205db15b25b66;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I702778e2f8308e720ae6aebd003938631b4a76341308834c90d10eeb3611ce3f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4473c0cfd2d569bc671ba814a524058946271eb49a04fc384e9373185e1f4a6b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id2ba36bb60a1673c62e790e5ad15a4fdd49bc397b3cba8e6251a88e63c249091;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2ba73f603d9cb767572f2b2f2a9732e2ebc066392aa85888df87da4dd8b84113;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ifb22aa4df653a2afecbf1dc570c526ccf003e19a0f5972b9bc5ba9458e316ba6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I82f10eef14d4ad82b1f7f8c5d056c398386a6cf790095113a615a8bb6cfba233;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I43fb6b8f15f49b741ef111f2b4a57e5da84af4d6f3ce9b92e0a2bedb18eef4bf;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2fd5dd69a5f551c26d9970d09ab0e26ac5183a0022af58e2bec1dd1efefb139c;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ibc1b6326c8e2b05aef237f6ded855eb730c445a3cb6c7d49293ef68b6ec623ea;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2fd258374a5bda5c58c1fdc6e305789a598fbe70657d6dc18e8878b6c2b0441a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I3a8bec62f5e0501c90baaa2f6f7288929d91d107a2197e1c574428638cd020d7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I76942d3b012aef2097112a1c1adfa2bf986414df19a633b87d2f3c2a61d27351;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie8930f54b7806297e3bb1082b70d74d5eaeaf269112a0d5f82caf5c941ff7a2b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ida428d199205588ecd8cc963ceb39e24bf6f2d004b675f3cb883960e0f089842;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I948dbc4fe20518395aaa5356bb504e41a80332a8adbba9ae4c6d8a4ca0704b7b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I91f0247d07693c53d716345c810ffa0ee8d3f4b793ca8831763f5465db649c89;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5140e483e7397c66b8d4835ac2e465f125e62c4feb9835d7a5f5ea7849def4dc;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I754c4c2dda64bb938ac60db8cd469c6f3ee0831a3a6b6b98e902c1b72663ff28;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If049a08cd46a811753b3637ee0a96207144b0a5eade57068ba5712c3ba23c8ae;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I567c2801d5598a057d5773ea5045f594de038bab88d554ad2c713cf56ef632b4;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6b404c4caf16f09360a848f09b33c16a69029ab05067f1bca94eba5e69701d37;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic9f57a4a1184139b219a3a5e3c554705469b79d3ab175ddc74512ccbfd5898b0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1efde896c2d2e97d2b635b34d6ad30d31a8c855ea5975dfadcf5ea136fa3d063;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2dc38e534505cf47f391eb9f4b090e16136d12619b4fe91cc8029bb5a050689d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I860fff7ccba78c970b447509ccd6de21b521bd8458673134640ce16c6f1ead4e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib83aabc196c7633dfb4a9bcb4b8d06959130620de297f9dff77b1454a8f2f96d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9786358e2588e06550a490e47029ce233b6d39273ad261316c5f730a7ee4bf17;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia23743e423f143b75923bc7b1a4363323d46ace080c8ee9d15ff687afd4bef65;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia01e9ec22c644f28b2be05c8002d4f576e816688e30965ae9f3ef78ca1272b9b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id49eabe82a09acf1b3a3aa3be9bfbc0ff958b96b44ada842e892c587fbddb8fc;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0797e7fab1998d109cd09e4aa801cd2dfe57364a83e9c84bef81be8f59ca729e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I93584fe5ab7128b24b2372bfeea00f7a2bf09d50b1fb535d01cc141c6d6fc377;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I035ba5b524312fb6136ca853695154f9334f6336e5acf5884beebeff72197c7d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I44142c70d3ba4660f5b85d895710afc623ed3470ba85eab3dee5e49a59e1b124;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If058a896104351e61394ece6dde5212381937b7d36a4b63f5e99a268d5c7722b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id8b538e6a6c4a147c7000388923f1d89a193f8ec53ef214556e005218d2c240e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I29e36792da89f6ea79232a191af837f9da3739332265e00d97d40b09ef384a58;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I658f9399a929745b4ba467a1e019fdbe214acd543dd4f5f51a95292420281401;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5e9d25157a8f35aed3b702ea5120ad81de73bafda0cb5811bae0fd0eaf2d11e1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id1ba70174cf019078c719d1d50a82a61fbfdeea2a13e21a1247e567b9266365f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I57f4038fbe1f52bf47fe1cdbb52088b800609231fa2007cb1ff941817005a0ce;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I797dfd66b521bd680024b6e46455d624aa58b4271f5e6ca19fc7abf520f26222;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I592de5159deb6cf98840aff691c78457fefe7ee33d85506cd1dd400679207812;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I74f49d84817f2467b8ccdf03acbd7372c58f1a4fddcce45cb882431b2be20b39;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I262ef0e0ef60c8effdcfb37ad79058672a12fe1aa6b0099d00f1067fb709c255;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib756dd9d8d9a5233fcd368ffa91f5d7d9c8825b01bc26140e5a717d3ce263e64;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic69f5c16ae27a74a97e7bc6fce24e0c868c1e1e5b6a348410853d40bb11f5d91;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1bb2be29dd44258b24a36ad9b1625ead1cf965856f1d9695c62ae80de142169d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0bba5d4133f73c77eb3812cb20554c368cfe3a6ddc34cc7405b33921fbbd9a2a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icbff209e6c8353c58f46c0688f06da0cdf71a95defd8937f2d52d63d387d74b5;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I98234b1225d9d3d636129139d51ebd098c46162cd51cf3530b9c8f8c0f12684c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia628bc749f04b3d12509effbd4e0bc5ac0fadf48a2cd5663e4c2094593870a42;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I31906081d1cabbb8c066a2d5377802f2366fe4f3993b4f749f59d89ed1fe0388;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5ac2c7b61022af9bd2550f824b8e129ca1c336b1ff900b0af785d86e33cf3358;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I735b667ac51f343a3a50cbaf5478e1095cf20f38a650d24285dbb38ba66abbbd;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie511320217185f90f1e4a23ab51ae9686801b09657c714a5bdd9c4e26f070bff;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4156cb61e9e7e8947b6750f177dac22866e9f9ad06d7e45bdad1304988857d6f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I032b833c683eaf0c1c4c60ad831278ab0ed11ed856361be3be59dae656141fb0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I45ae7cee40ada2a73a62a90f141788d37c2a24f503646ce743ae4ac3e43b5bda;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib41d86b318a3004b648c9a1b0ad00bbb144511fd63b1c7648cf3ccfb996686d3;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5ae0ab8d5ea922fff8bcc268c8f3bea87f11b7d6b824787e972c00a9db0be916;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icc4bebb1db4145f9cce0fd4c250f7501f300b6cde1f31327d80b844adeeca1c7;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id33bc2a3f235239565a24ba23a93a90e564b2ddcc7559044ccd4f2e6aa6fdb6b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Idead9dbad4283dce602c05f81e98610ab7f65f9911342174ceff7c95dfa9ddb0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I86a468c8931c4e794856a1c434471a885c62c94dbbc95059bb67ec45a9a722b7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      If7060467d2fac9aee8d69c5ebdc24d515a657bedea3da55d13ed6ed4e3c8e79b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ibc857d78e207a3c56616aab90400d7f0b57c62f4a5e421ee4b5b7ac7bfa1c31b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6aefe769159bdc69fee8e09e46357993c13dd8ec9f059cd51d43944ecd7ce3ff;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I275f7df80a91271f558b5ab22bb6a5b46f01973b93cccebe198f0f3c6e2f2cbe;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icac3a5cc88034cf8211c158a1bee2a04c228afd4eace1b50c7460ad5331ae02d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8cc2be0175b91e2589ee8980b860af09aaa4a81cedf23de18f9ae69d0514c369;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ifa5d23491b028cbdcfd79fdea2e0784f068c1fd381dda7ebfb5d457800e510cd;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia6661480da7ffc0644e0a42782e89f84535952e5f17f2ecf3f1e4cfc56c532d5;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic27b23bf87ceb2ec2d6460321286d798980f966c89d0f8ea42a79a0549b2128e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If4a3892f82907488395a090155f489b67d9808fab6c5f4cfccde65fc41d3b92f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I01500dbf2528609729acf26a24c11bab0adf8cdbc0633527f21644816cfa0dc0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7b2b5024c5f6f54ab62c8e703f603950e46ebd179fc35e2db34ace053564af4a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6db96717b6fe00f1f87347adf69ce2d4b4464faa472ca989bb272b36454e868b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I709336ccea8dfb4b988c870e3d5c854d77a7acc5ff842b9c2c7490be8e10b3c3;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia8cd57b3b123e08e2bc00f82da941eb4431cc816928254135dd13ef52eb9c03a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6ad8cd22867ad477cef7562ef157f85bcd0aeb6ff72ceccd15ecf5c00faf12d6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4fa8db615d84b02196afb2ad926769bcbfffb7c81170387b4d460c7403f0dfab;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If4a806d211914f82ca329f57517b2d1b1a60a8381bddbd3153e78418258d819e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie81813a1836449254acfcf7674552545d2cbc852ee2bd2f37378345ccdfc61b4;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I282657b255db6edb8d72272a04f6c69d5b8f32795992f902cbedae3bffba4a4f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id9fde3ad430d66c92a5aa6797b76ce147e39e4245ea761e36d81214e7a02b4d8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia3f8a8cdad50f5772d19748e82e1e9e0558a1d7973bc2cda424ba8d383c15d62;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8f2cae5483691fdf6ea64a4ccb2372967aa676835ffd4f562269bac888840d17;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9ec9a8bbe81467bd2ec058114005f308873b8eb8a8c939f4002003402bc6c486;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icd8572ba29de1a399bc077f53730492f4e89deb95b9136608da0d029ba60ddd1;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2a951c202348bf2bb4da1f79c63a8515c95484c9a16ac1fe9b857fee59361511;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6eab6bb656dc82d656eea6da9dea574b230f56c6ab898a7f80973183896d8347;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I009b4951ca9d1200c6e7787f401228a9af483223fbb4150aca223cfbb80c8b7c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id802e388c3b33f7d0a0960e0e51da02e7128da423d518a916f761a16b73c17d7;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I3af56e36e8422acbbdb52c77327e09618a7b89e21e35787ba522cb8a322ed0bd;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I47507e717446a9ca85cec7e5fa382cfe435affddcbf5b25d4e74f23a143b02b0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Iea773cc6750944ca9d0aaaf2dbd818c485ce25a1e333978a68333b521404516d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0d76ba051f3db8c1efd9a8f0bd0ca77cb28c7dfd68cf4c290ab00edfedb15237;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5e0342048fa50ff3b98e175c5c8aabadb97e925dfbc34fb7f68376b8eaa3cb1f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I39dc59000bb2e3fcdebec08ddd22a460fad0c09e8b68adc7e72a6e4c3025da49;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie03375db3932197354d4fdbdc800b2b7134470f1622806909963ea424d5fe6af;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6db1df05e1ea3d8011bbd6e08c9d50d91e672a20aa2448167343b839e8f6f888;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I529cffab52c15bb4db9614fb7a0f353e2867564b31984bd2c5551f5a5d407fbb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0d11d2b76d26d33ebe0c7577f5d7bc68ab8f4840deb765b17f4f7fde0a4b2fae;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I3bd4e85424803f9f3607ec830b6c73bf1d273e7de387d11359eae7f842fb1551;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ifbbf33f600185eab85dd2c0dc5ab2f5e0e2cce52373cc2acf5e466a2e27ded58;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie54a4e9ee8bf7646b7e69193c8121ff42b4ab2f266c49916322dec059c92684d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia38b628fe0740039fd44aa0a75c751e1a9e176bfc305a978377c1fc9525c00e4;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic07553da54e29d977820e271e50502264b236c156bdf4e3a654cd948a6d4f726;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Iaeb5b860946e41cde629a762ab6e6ea4a0f177083c9ac84d90ca99fcb90e7c9a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8ba1954b4d7af696e80f659a70d18bea70c37a8f494827a2778c421ca1dd8ac9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ibc0b2c21012904530a727f0c5643b5187d7bb8706a308bdd0de67a80147db974;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2d1936d0e3bc9f6320f1311cbde5d8e855ebeb68cea0b8c3dcf77f3dd63ceb84;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I008d6180d4774d2472158544239ee654e73570389873b54b695946cb78ddb7e8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic0b3a57afcb2e31014f5c80d84c8eaf5f7f20d57abd8e863e6ffe0b8146108fd;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Idaea720265ed96d87e8852c36eebd63e2be5b9768c7803f13fe85e7532b75ea2;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia7f87cbac38cab3ef1ce6466b6b419127464ad3172cb03af43e0f75b9575ff2e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia7bf8296bff6d2322977b0a31ba519bca04a1d6c6f6c0cb5a47e3408bdfac573;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I27a670adbcc49dd11d8a6647a3220c4ac80946eae616e3da78e7a35f5f522502;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2a69131c92e4454ec846c7528679731db69a2aa63420f0f22289d5c0be743be9;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib913fea37f6ef92b53b6ec87dde4020983e78b263662b92008f7241cc029189a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia5fc094477d9d66d7fab491b73a00f50abec21827f63372fc1b7e0bd31ccf375;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1b653b0e5ffe67c25c7a73b1e2fc591f5e57174285113fe2c43ab123799c556a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I41d88c1cdef0448f878686d88600bd254e722761979a244cb1d00724fc1d35d8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I068d321d442274e43788076aecb6c24130003e03ced4df86bf13a33d2ca5e1f0;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I85e825a905ae7dd292f400406048736ce90fa7d47b6dc5507254283662fc7564;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I975a1d7b1fe781bb19e80aba369e5146327185746eb5088542eba76fbd88ddbe;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I80cf17357df8073b050d80de366bbb919c5f6c8983ca87f6606a84df1b92c549;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6668b8618eebf7c40e35e5a06aa3b131a6ea1b668bc36d9731036b61087013c3;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I68a074e808119d0f33d54d3863c907dd5d761b3f6b144b9283e67f956d5932ef;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1b4f3dc17b05ab02ad55643162e80975cc4802ba8cbc4323fb017859b3617abb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4aab61ec97ec8dfc8da6d2ab5898bcdfdaebb0f024fea498a6ecbf0bd15fd1c5;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic69eaf55d245ae896d42f0f702ef6cd804be0d02cfad9f883b3dac30786352d9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I26395ccf79a44d582b559acac5845eae4a01464019f7739b7d52d8c8a4c11154;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8c815413903d61f8d5f9a8abbb8b5e6cb133bcf0e084f4a46ceb98fc67f67515;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie9c493e499f4b2aa598c54d5a5afdf39447612225daf7f9f5b3c2a23b5ee0ff0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6abdbd209c6b52b3d4c69e83d51d89be9b3b8e719e4f4e15f50afdccb21ea02b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4368873c6f3e3d6ba5e7e83747fb90120e80de634655a9d2a97bbee88a9d8501;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6f2bfa7344a4516d6e0b959405ab2c16aabea8d70a454d4eab330ffb6bf9ce2d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I082b315a51a6a180909ea4f576a9a3c8b0550e64aa222610c2e6906ca78aebad;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie7eedf6171b2af8aa5e550f07c6913fc6e02bde23689f5ff9f035b89ea7f4cfb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I23872b1af6db7e455f25a7ddcc050167bb10de0afd16973c0a90804349210372;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia298bc83a87ee16d194185dec24955ca32e85a919f168cbfc79e0724038e43d4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9796589e7a8535d47d56f792d80838aa402e3c235035b517765096d2a6843215;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I78dfe767d8265759b3b1488f6788812b210a952cba86301b7afe8acd0b194947;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I46d39260d96216c08b7940ea3bfe542bdbd0966f5e798321bc90a2a00f64360f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I12a747458626b92b4c562f72f3e5fb63a575053284698acfde64b482d44a98b7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1033817563ce88e3b26188a88303cc6703f47afdaae4d5457fab8b73bade5274;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id27fc6b236852c780351e17ad6e85bf55621c84757b3014ead5a2b9ef31d2ce8;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I343bc73eaaf00a82b2674c8cdfbbc5c6ea52d10fbb9e9453cf4fcf2421b97e47;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic117e33adf22ba594c3e3c03966b6bb0c6827c2c980f6ba1ee5f6ba40da372dc;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1af6f4d00567aa1e302e7d8830d761e7a9a616f5e4e958b264701c476216de4f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I223d1009ee5643d0804f1d58bbeee2c3f61d8b120ceadf46556e379e45ccc061;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1682f44d820722e2566b0d6c02fbf3dc72547221d519ed071e7c7d77728ba21e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I60bf67e044d9694caec17617c4d9ff59b9be7698c17aa034515ab1cc94d6a5ed;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      If0095cd5e911c91331d2ef6ab3866101080b3cabe8d1ba9104b6b5ae5d18c713;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7da66be74fda28e419201be145b24b82c9b29d1155ed00f78e8907d584e214c1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      If7f60dea1e83c3f86ff8ce3adda8214324b2064d06d69ca68477288522ad9de0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Idfaa10639faa52207bae09b46b05e70da4e285f83560fc415e3915d0a0e8fa4b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I3b1abc53d350b3b39e60c3a5725e5a21632e7f0275988b98c1fdaeed5342f9c0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ifc9a7a5a4da00db6f00362e2b2b91e1ca59a65e8e35d66791a13468302dd081f;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7943272afdae80761f8b673788c92e4461bf3de3229f7addec1e54743b11beca;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If453fce64c627db639d688b2260fa70ef90f802d31cac666fd4cd757cd574682;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8417f8f367de885ebb86571786bd964d4a81d6712a88c3a8071c08d13cc7cf58;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1eca2d1c9da79ade1c32a3685553f133098e1e40edd1e8d9c299a961627aefbb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I653822ee3643c81b817be0d9c3f682d0c806ae17dedb0cae5b1aa0ca914e6857;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id3b8c5a0992cfb8a82d0e9857a0a77472fe0435d93e37978bc77770999bc4b4d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ieb917f5db48f3d352eb252f6ce309bd972cab47f09ba1c140f66192b260f3925;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia5acd518b995f7c0cb3e2f5303601027e6195fb82489331aa60c3fc8dfb21184;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I313a01d9fe403e838310c49dc37a50b738025400e99faefbd9b8cbd426edcfaa;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I588a95ce70c7581d9afef4d4a297b619958d34acc8bb75e4d61729b440945a89;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1b81a8a827bd2222ea6820d80d13e537868e0157970625d628f0c062733ec3d4;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Idaeda6020813227d8f52db3ade5daa8152deb71aad3e8cd03094b66b7af5696c;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5615438871373f7ad838fb5e8c24b9517fb94ecf6627c803e66a78f778fe9c42;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I48f239b0c336ab3fdd25e5b7758a5e6c3c0e698832c1f4518d3d1bc6845acd41;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I07f9ecb15d2696b2cacc35c935b497b2f8cedc55e2a661fa57f2d0783e6a1001;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7226b2d9a70f4f716635a08aacafd4ef7a6f5fd31edaee6654bac5577e6398c4;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7fbeac90b85dfc78e20281021fc1d7cc90f9deacb2091ab55ed07f51fbdbcc11;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I14a8ff2f5afad37ef2f9494e67d6fc7df5e0960766ad9f9c46964287587df5ed;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I46dfb75396740f84b7758552420a7ba8693bb1ca5259a67530c588585de1c337;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0b4e726e030569d30af5272062eab7426f9a6c50a8e71353fc19fa3b0d576de6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I60e36bd866a477c35110e2688e7fbb13b0303d210e014c9e151b313d130101a8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib6234dcd7696dadb4fa7903f2da1ddf0a7f469668b59cde104d9fd751ebea2cb;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ibb36dcaba8439f48b18ad2dc8399df26b940f7cd815996635da092d41ee5b106;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I07dcbe17d78ed40700955c3277dc667bccfdb936125e6bf04e0e0ed08eafedea;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I387a4fa48a52a029d2bb0c8e5163f15c4cd55d570db8d89e5f73d7bd6e21ae5b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie14f4f4bb4b43f4c07d648f32e6470bc1626117d46a927a286a64d093110e0f9;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie2ad7096c10eafa6e451ff7793b2dda562b6623b1eaeed56bbad4019662851ac;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I099c775595305f8021cc03ef225be27441e325455935c0545cdc553d0fea3d44;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9de97cb2569312c40a541c0038e02c03024581050590e5677dcde888f4c6c3ac;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9bfa196a8246cf5ae88343b221c084738279254b84fc66495e4669083ac05ad1;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7a55e4af3d00a3684ba08ac52c3dc7dd0188efbb684b859ecf017f783fce247a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9fb047739860e32f32c612e35c96205de22487ff301c0fc990f576bf205b98fd;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib1644713e1c2c63d093c8af3a2be146dabd70cfe25a1a6ac062174576477b113;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib5aae92803bb8df9f7ffc9fe70a6f447be999b64f9d698828709487924cdd4db;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie907506d9949011db3e41c72b9581fb832dfb29f82249768fd9893a3de358b35;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id89ea99f9b791029af271f9916f63681c6881dec4351cd30a7fc9e3ff1b81400;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I678204e14a0213dfa7135814f07e5f6c4d12452a503ed555ca2c20c10f047d5d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8f70e2b5b2ffcd04b7a84ba28ab51f0a9dafd95e4628df8b36dba0ccf87c666d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ice68b876a3b3943637914d8d12aec7fd37cb867f7a7c20be11a66dd85803827d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I21a71d60d8728a63954973b41b85f8ec46e1fedcb5208ea2397adfa9e58be880;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I35e112474e97e65f8e8aa9a4dcce274c7ffda9cdef901ba31801b4daa68888fe;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icc2b71964c3f1484faf865db6f25dadf0a84b62f85a86cae24a8c01baa1ce8ec;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I84992c3714fef30f928dc3330821045f20e176826278d42a9606f2dfadfcb9c8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ief6bd3a84efa60cd8d09e7f71dc4b3b882f2eeef86edace8634b6355a0ce5db2;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I011fbcda61a4f528c38920d0077565c4592c5f6d1a2f5a1a7dcb6a4a734e0c83;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I21ed781b8a01923a17f646d965cd22caccb44b555b8f392387269b9a2ec9b647;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6d2154a30adb0faf296cf58ca9229eb1a298767fccc4a1214092a2b977f7442f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If070967e597fbcb6a0ce8a28166d084e71daea6fec72b92cad9a59d03c2dc531;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie500f9b1405b49a263908c145ee4a337f2ba4cd2d4d784a2acb77068d09d1662;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie0c16d4ccdd2d7d6d9e45d2eea233e13674b7d5a1f8f41877267074f40f6a2bf;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I26997f7f737ba99dcbde55d67661cf9e4efecf397b1ab3ec59e0cc5d8654a75c;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I731f6a3be9c5a884fe93ef383fd933c14af1cfb64cd73fc4381d91d4faa2757d;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      If6181a32c0ba3cb93e47ed1f1279bd4e739882c2905d6d64d0149f26d052f0d0;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I77f33c069479b582cee609a1e4f6255628bb7f6f667e6536333c8e99dac1e08e;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Idb4bd19284288df2a5b701cedcd57347e4f7c37947ec1588daedf3c9ede0a12e;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9288b2d29db5e8dbeef47da923a8ea2055a38ca1f37d4d8ed5d458408b154924;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I4be880e4f25fc41932b9ab9295794ffa2f334ee5338ef0d59894d18918d3e0be;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8e09e68977d9f7456b662b0d7fe4575c48ddf88f897bbda3545f7b1b63d89ccc;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2dacf26260c042fa148fa6c4e97bf878ad2e89e221acc0616141e1841b0c320f;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I53ec51c004b0546b3dd0563e2c294a6c4b95b21301321aaf80c838931473cece;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6cc3662b07a43d62f870bc24d55a9e5675a0e50d923f3b293d7004c2c62ad31b;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I3c0c87041c080ddc72a51a1b6a4fe12cbd62dd40515520e3924dd8cb63728a83;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I670beb5586ec69af20e65eeaa49be81826908f01db21d27643e2561621962b87;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id9bb31b77b580b8375e799bc74c4829818ee16c05c6dad069736736dafa7a8f7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I88ba583883fb596ad6cc6716008143d6b643816e8e694ea5f32ba95f3cfffe48;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5800b2a82f1442915cabe6307e4eee8c6b4071bf852ca93d4a7420bd0e6b1e24;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia8545410ad46518007f6812cf6132f4f4482933818a0fe103dae14b1530518d7;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I40886d5f08de09dc76db805b27c8ca792ccded54cd12ba2e6b70c30121ad9f79;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7018895fda9af57bf39b18e9edc144f8854067ef25800ef8eabe76015fc207b5;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0cd63486c66b03be7f8f629aa2577ef8849fa2408aa41a58514c75db95432892;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ib57f995d569a522f5562976385f777cd6cc39ed15491d0ad8f88cc0e908c326a;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I8dc1d4da11f5cf2226f4d8211654acb056d8fa751da8aab85dc14664d72b21a5;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I35636bd5c56cd95d41880b5c936108a3ab7c1517a8e09f76731b2154d39c87f8;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Iaa67bf8b75feef8789908b65a38dd8124db04184092d5a584054726339440c63;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I84280195e0f72492aadcce8eda907d5de2e05dc16b9c5ba1fc2f345192ade355;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I845063b254fc4b71844ce1e01433e1d8ad7e176fc80530a73ecb26c31bcf8bf7;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6532aae67414dd9e03b874fd4b6a321437892a7d89bab17ec2d5a684aa9ad55d;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I51b1e937ea9e8b9d8f3d8c8c66d7f69b172137911df42ee5fd10dfc5d32bca27;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I7032c41ce2651dbb03999e2120193d71ed608e40ac2d51329837f3abc0a976b9;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Id90613f9d2194b97066ad1f5247ec5becce3f39f02d165502d84b92178a02948;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9a800fae8c9498d12065155e7e781ba817ee2b03ea6540813400bbe438f4691c;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I38b86f50ae5aadaad749bf30610fc173dbfebd9d3c9d91147b1b3afe8d7f1004;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I1dca7dc76f83994b077209eb2742069045e743b6eb763805cbddf87e6a8fcc34;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I12d2f80160672a05ea5c1aa8b8b52b7ad7872b05584cd462f2fd449b06326ea8;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic16409f8fa42d6ac05643c3943352c03f19cfee0c3068e96d6ca3630b8f2cacf;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I08cb7d15d8198cd0c19dee6c97c2732b1f72f7e00294bcfb0887c25cb0951701;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ic66f776d5d728142606f048e3cf27e927f094082fe1dd31f90e757beebd5b5e9;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icf9ebe6aa27457ed3d8ac986d9dc8260bc590e8c778585764d6021c62b1f9d5b;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Icfe7c47d401f26676f3f8f13e34894792fff7a3881d754de5b4ac1130cfad989;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      If4d6db4bdc3cf9677389d183b78d9ce032dbeefbc9c6374296777d351a8d958a;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ia6852c630d3d698cbe47da7b990ed04d4e0b995b3d765ff6a8146da11e42dea9;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I15ae50aec5944edbaef4ec461dfb5ab01f597a46233c643d7139247b8bc2f6c6;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I5e5d78a5f1d49833052eb3e84c516dea9f05d6d49879c593f5e0b9745f84fde7;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6dc76307fe143582b214c945a6c0a35a4545c8bebb622615b3ff784edeb2d0b8;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I6454add174b2968c545e831c5bacd6b95b351b7d68448b3fa9c2e5476a8cca35;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I831951ac212604dca0a254f80af9c1bc9a941f743abf321cc91063922eabd175;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      Ie062df11427db764a0e09705579e134d08f4ed2a027e913a43495db5d5fb9051;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I0d347b21cb8cd8b8a0fb2e002b97a2078bbdf1c6e71a0e4b9cb022e2a0db8de3;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I2a2245385398379002074dfa174bde148f97bb3bd83073505b550c0c0bbd1e65;
/// If852628b048cce63ed033baf5d97ea58a853f438408e0f7943a317470d67c426 I0c9618e9849a62c68ff5b0e62361c05f4b70b181db1ef47eed458a17f5f4f3b6 bit
wire [1-1:0] [MAX_SUM_WDTH_LONG:0]      I9c8cc6c27c1fe245ae54ee4a9dbe2f5fabe4c675abb8af6a49a61e6076233e73;
reg  [1-1:0] [MAX_SUM_WDTH_LONG:0]      I862f2564a9e7f99bc8370fe12c1a5e57612d564f1606a21f6a468d558c23fc5b;


reg [MAX_SUM_WDTH_LONG-1: 0]                I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6;
reg [MAX_SUM_WDTH_LONG-1: 0]                I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac;
reg [MAX_SUM_WDTH_LONG-1: 0]                If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e;
reg [MAX_SUM_WDTH_LONG-1: 0]                If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975;
reg [MAX_SUM_WDTH_LONG-1: 0]                I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85;
reg [MAX_SUM_WDTH_LONG-1: 0]                I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5;
reg [MAX_SUM_WDTH_LONG-1: 0]                I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55;
reg [MAX_SUM_WDTH_LONG-1: 0]                If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93;
reg [MAX_SUM_WDTH_LONG-1: 0]                I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6;
reg [MAX_SUM_WDTH_LONG-1: 0]                I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727;
reg [MAX_SUM_WDTH_LONG-1: 0]                I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733;
reg [MAX_SUM_WDTH_LONG-1: 0]                If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c;
reg [MAX_SUM_WDTH_LONG-1: 0]                I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84;
reg [MAX_SUM_WDTH_LONG-1: 0]                I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc;
reg [MAX_SUM_WDTH_LONG-1: 0]                I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7689b1f287170d28fc72712f5ff2fd209108b000a63e268b12da08dfed6d60b0;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic114200c11d550dcee2bd668ffd91dbdd193a00571dda2d6f99b4985ef999f83;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2090cbe74e266e4385d5075f2913013cc38b26c5332d982cabead5dbe52d7775;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7802f219761d40fb4b24650bdbbc6faea69cf01618fbddae575028e96aa7c627;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9e11bb32c337ed1d87274c3040deee6d8813fd3f6795de87aeab9f93686ee409;
reg [MAX_SUM_WDTH_LONG-1: 0]                I08382faacfb31fa012c97cbde6527792abbdf2c9124d886540d385dbf39e24a7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5c8ffe997fea9d77126fb36c6deb4f9b9c9b38e6aa562b574011ee5915a00857;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6f9b56f1fa7e83cc6acf75b74037938bcd08ba89ac2cb3dbf4df512fc9d521f8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3ea241ea179029fe0c486fead3909ff2c05b2d47e4484549d1d521a4f891a9a8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6f9fd1c4756d8d1250b0ed96355e2739d3bcdaa3603b7e1cb5cb0dd0ad5985e5;
reg [MAX_SUM_WDTH_LONG-1: 0]                If084c3e6863c87018f76e95d715c83cc83dd85ddf7664f98c6ff35e8a0ea40d9;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7fcd9ade547e48c042200e4bae7d4699b326df8a285204b7e23eee2a019cb01d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9207b21b45d4265cc52ef02ed257ea78cc5a269d98165b2a7714a25b1c477521;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4322d4cf469c3caa560e48f6eb1fea264c42dd76b65977c24c676681518691f8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I924625bbe810db6c8d5cca4407571d5819d0f7361e2d7f1906bbeb822457aae4;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3a01e4ea96fcd387a6bda68d7d07cd6b4e89ca653c798f08ac8402696b42a371;
reg [MAX_SUM_WDTH_LONG-1: 0]                I96114d8145aafde7f8f5666ca2f6dcea9ddfe9796f2e3a54556fb1b23fb1a331;
reg [MAX_SUM_WDTH_LONG-1: 0]                I006672e4b2c9c693fe5b05655ebb6f31e96ca8e2c92eb488cd28e5a940e49766;
reg [MAX_SUM_WDTH_LONG-1: 0]                I408f22a4a77906024a2e6ceb970b39ba9ca76300fb2584bff35e37da452c6613;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie84e7eb709edc06e55ae27284cb93a0c656ce8559679c49a47c7f03f0d64fce2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I84fb24aeaf533382e57c00dd73683ce0e4f5f33a0e7a3b36f2ab00732891682f;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ifc8b49d8467101e2eedcab4b6ad6a73e4f657c0e995ccaee5dee276a5ae916b2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I001fd8ecbe068f57df7498db3f519cbb5a65bc5af187f1d34b5eab3df45447d9;
reg [MAX_SUM_WDTH_LONG-1: 0]                I11745815606a2dcec9059a24625e93a31b0f15d9b81c97403905e00d3fd64f43;
reg [MAX_SUM_WDTH_LONG-1: 0]                I37a341bca6a12362e49dae8435798cd8e7550a16cd506a7f852f4223088bdb4d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8ab2f0a2c9cf1f1e0401a67f3749b106fac7d45293bb9648325f330e3230517e;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic6ce7ef3f9390c17ef23e718bce985f168504ddff0d66e2babddf08b37dd2819;
reg [MAX_SUM_WDTH_LONG-1: 0]                I26c16ba52eb0f661ca599263265d1d0d7e1f155b4afec85407f3ece6fff3c391;
reg [MAX_SUM_WDTH_LONG-1: 0]                I31afedbc324d4ddcd04b3ef766154a6414cc6e31eedb0ff24b40698430e84927;
reg [MAX_SUM_WDTH_LONG-1: 0]                I807fdac75cca555b8d81d1b4d7e53ae7cfa0e4b83bcb260cadae218faed4f781;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0f8a9c8deb02bf990a6ac2ac0569f9d0ad9f167d7c18dc70ba544912aed4bf78;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib3e6663aab02fdb649843c552944b6e325240f5010acb414c311ae56e78f8459;
reg [MAX_SUM_WDTH_LONG-1: 0]                I41339bac55a76a05186d632423b1fef8173940f0cbddfb64c83282af5cd04cf6;
reg [MAX_SUM_WDTH_LONG-1: 0]                I28fb4df9f762474ad496e8689f21d13bcc5bd4fd79190892b78409a06720e2f3;
reg [MAX_SUM_WDTH_LONG-1: 0]                I84ce9c6711b257cb8cf2f09bcc02e0f03490605e543ba12942207df6fabed5ac;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8f3d31b6843ca54e80e8f61be651cb7788b43302b001d791357fad349785eb1d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6fb6112b591f6f1495935e422361833f041f7231996d88a3936b5da186e4c48d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I959de6064e6c31bf0d18c2d6b4c274ebd5e9fadd996fcb32e695047831716951;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0f46fb1c05f0f882ae878e86285077da38a459201c305e13fb4925ba34eaef8e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I99e249a8eaee9127d347ab629dc27a21d5b55d2826c354eaffd9e6fec47b1043;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2f779bcb2996facec77594ce5efd7c78acaa443f2b6ab3a5506ae96dcb986b23;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia765277dd8a5fbb2a65aedce2934fd6c4dc9daa4e0b316604f6f137f19fd5d25;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1a47d1294e98ebbb0493fe3cf7743d1932eac70fe9d2754367a51d9a49448d12;
reg [MAX_SUM_WDTH_LONG-1: 0]                I71c11e07942c42d17f5b85b1da8857e91f789966944c1e0948bf5f0285c91079;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id810b154e951f2b2d0b8ae826f31effa4f39b3a0396d446ebcceedd7225c5018;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2a96d9fee197ec3bcdd50abe43ee0d3992f5b03db5cdc958771ed812bf3a0b4e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I280a4a7c5231cbfe245c071a856f7d1560c4154e9f9a4c5fb6895baa2f4f5871;
reg [MAX_SUM_WDTH_LONG-1: 0]                I01562027a6c7a542ae356bb1d0db0dc55b2094f3470a1894e67a3b7fee9e4361;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie3eb1aebcdf48fc8f41590f0e9524e989193fd14fae379a200c20d1fd3755db3;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic585c7a7014e8bff08f28b2d432e9783bea57ff5b456d851503a2c3eee80a768;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4f0a460fa116f5a45cd0c435e594ccc7597b449cf5205391a2dc6e977f4bdeb1;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib7f3bef766d8e66cc9002dbcf3538dbe974b70de4d7a8a3d9cc3bfbe815841d5;
reg [MAX_SUM_WDTH_LONG-1: 0]                I027d6136f1b64e5e2f94af338f8fbc0ef9fdf8dd0a2d58aa0eb6879557361681;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic62f1d181b6452f30ab2146b4e43113b2ca1bf21962f686be46f59084d39fa0e;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iecddbb8ccabf830117fa8836a6eafc8dda6fa463d9c907ea25d298249bd066dc;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5a2b6e5bff0ffadb36a7f02dbb3cf48ffd37e6e29ef09200db12ccf9fa9d8450;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3a9d955359963dadbc16853d82bc2495f84c37d8cabb868a144c5f24d9edb2c9;
reg [MAX_SUM_WDTH_LONG-1: 0]                Idaf457dba6ceb8f056ac34d3bd84bb9e9554c0d55db8928b9b48692c316e6fc5;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iec8531839aeb35f1c356e474abfc871d1ce889c4aaee1b37b272dd9650fb6981;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6a320bd601e721d94d7ac0aeb59e2c81a0a9737d2f7b49d668369336dec2ebfe;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icd9be4d5172c268eba385d2cf858caf3450d81a87bb90fde24fccae0d1637d99;
reg [MAX_SUM_WDTH_LONG-1: 0]                I64227cc72d5c6450ebded626fdcdfd149c8e29dcd6839ad76b2b9a932817fdf0;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic754b281b704937ea08e702dcb74b7175f8901b29809052424f867a6685c1d41;
reg [MAX_SUM_WDTH_LONG-1: 0]                I861b39dacbc8ae1c9cb21a407a53608f0d5adf148148ddb8c3ab1cbce25e2497;
reg [MAX_SUM_WDTH_LONG-1: 0]                I994137ceebfa9f1bfb6f3342c02ef25b1a5e881f6fcf6c2e7f274663b5b4a3ba;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5193db4e129f33dd7cd8691b74f52f030a066b583bbe2d9a4a6e9962f1c43280;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iecd0fbf7643812e36e8d17ed6782ecf4b181df9d284988b1f416de07cdfe6095;
reg [MAX_SUM_WDTH_LONG-1: 0]                I390b2f0e16e0de51443f9cbf8ae301009d17581f5e20ec4956a8e95ede2c0822;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia733b3c17807a98828719894627b0a1fb161ffee86fb28c11d92f5b185a6284e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6b87b44befe3363656697619cf3dd967526646ced0f90813c24c960ad4d57d5f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I29ee4a3cefb214cdfe60e6907e63799323eec92930d4a48797c96a7c1f3e3a15;
reg [MAX_SUM_WDTH_LONG-1: 0]                I748cf7beef2ac47341c77503d0042b6e1570248031f1d9880d0bf14969378379;
reg [MAX_SUM_WDTH_LONG-1: 0]                I559b90a32f7cfdeb35bcf30683787c6357460614330553ffd4f5732cc03507ed;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie6d770decdaac3d75cd6c9eba7edc89898bd152a7c75f43a464a47c9994c9a87;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6541e01880f3c658b3404a81e96fd03b861ba4a26ec927e9c2c64aa9973dafc2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I184fea1e133f0a5b9b8a88926ebceffbb79cf7816941eaf9a326764d876c924f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I78d3ad872172f1089358c601e00c98f526455a961f30bfd6a966e8d8bb6bd098;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ibe18bd1138dcd8295a35b807d811d5b05b07df9efd2326d0cae0cac6589e7bbb;
reg [MAX_SUM_WDTH_LONG-1: 0]                I68fb3ebbcbcaf18cb81eeae19529cbcf7fe4175df44bd847d87ba9675ffa862c;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id2154e04af88ba8cccdbe100e1c4e4bccbffee35bebd3d43f9229d2915bc1deb;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic95be152c428a61c5e57fa5a5e776b9341efe9f2d08c73fe0a9d2663b0a974e0;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6e7d06d6c6a765e6994847af070c889f9c7059754ed634122e0204f750919234;
reg [MAX_SUM_WDTH_LONG-1: 0]                If0343bdeee565245554859329a0188f1267cab02c325fbe93d4df18606760025;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie090cc0a910baacb33f7e858eddac0b221b9a5c567ebde9bba44380b06e8dc29;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ia0e41f1ae6bbe04c95f97b4d03e31d86b4399463bbd9fb5bd714b9c2b58bb23f;
reg [MAX_SUM_WDTH_LONG-1: 0]                If4a86cc5d7bf6b2552861b330822e6bf86fa60debb5d503d86e081b720f3432e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0d2ad8151436f1c3336aae018a92e8bd400452c12972fef401e7ab55030d285b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id2881f7fc5d7a68a4583d24b1a8a9e09928ea1e5e3ec22fff19d4d59e12a201e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8733749031c60ed31e2867dedeae4f9ddd4da169ff086c567288ece5da43decd;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9180b03e001160fe9a51818e7641c427a35e0b2cbeda9e6bc0e32878bca05815;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2f00eb344711414f5f6efe7eee64b5690b4610385673a7186711075eeb319cf9;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iea8f3fa357088442ab8048febba14f1e6ae367c6b1a854ce0b2c4861c4a2ed27;
reg [MAX_SUM_WDTH_LONG-1: 0]                I0d3923859952e0ab6d926924645383b83904ee287f1783cdaa7f314b171f4171;
reg [MAX_SUM_WDTH_LONG-1: 0]                I45f444d890e00116a19e16e3c50c555419e910e2413c0277f62032d6ff66ca15;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic67dc4f0898ca883d489eab901e11caae2adbe1c1c502ab57f5366cc26d4d335;
reg [MAX_SUM_WDTH_LONG-1: 0]                I89150482cc550af995633308cb14fc4aac6984b8c5bb09ed4018e5692f8866e4;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id4c7f10c8e46d38df8e36571905e342a0b283e8badd00d3e4081890010c25f34;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3c6ebb6c57609827961bfb1e39059b0805cec40a48787adfc9b2b138a5012c9b;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic8177ee86d033bd8ab95b63937a4f80b02ebbb66d4c16d84c8822d133e7cdd0d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I65cdf21d7c52f9a1fd2d4bb265a678e8b543e0dedd9fdc5cf9e12ecf756e66ae;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib047d12eab2012f21895617ed9bff57a0678c2c85235301fa1276f99ecc8625f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I4864402239c958072b187da428e64688ab13cd5a3ba940785ac5086f81c50e92;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8d03bb3beaf84d3f94a15648cd5536d5f14020daffea4160bbd12426018140e3;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id3b64ab87f29683b9210364e13398a54c486d0b8b8a7a5ec6f15c29cf752b5cf;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2f3b819fb1f865426e38d2b39a1a4a8ea0560e0888f19913e2393d416205f3b3;
reg [MAX_SUM_WDTH_LONG-1: 0]                I23e7ddde350dba3f41b08c523c29dae580b57e09b8fd9d35af6ba3bd4b104b6e;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ifbd6430f8434621a650f4942f3be3669bfaa802cd912188e4139542d2a64a511;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1cb9b876fadc25322c3f466b101084a68e5a283260303beb238d55ca788523c7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9bd2fc6de34fc3d410b3d5e30c2e9e811c7063afaa6888afd119cdc02e39afae;
reg [MAX_SUM_WDTH_LONG-1: 0]                I9e9c82e0f8d919f8e2e03046a1654698592da05002140ff69fdd551598618d59;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic9fded9a702f4299431ec45bc00c9111907d62279133f1a5f62e5f6527823aaf;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib95adef89f659c6d98e43f4a9c43340a0acdf273ea6bfea0b8e99f0751c250e2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2f3612471464f3108bd427b6427c8fe79dce2b8e23dc4bb74cecb7e89a3b64a1;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iccedefdcae7039447a6901e1cac8bf962a9f520d3b343c2b00e654c7e11a24f2;
reg [MAX_SUM_WDTH_LONG-1: 0]                I8252bcef404ae08a2a748c98d672c368fbe4187f26e788e54d93af9077f92a20;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iaa2493521eb50d228c5b0619dca5c86b89a165f9855552ce98021778cc196f8d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I69d7f0497be77c5b1457ccdc35789d454bbe83f7d9eb458527d737a2222c7796;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2c40224a96616b7749f39d78a0c07514232a019bf2c9ecd7340560f5aa5ce6bd;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id95e503df18410329be5e7761b6857182c75f7d2b0268d0fc377a415c89cad3f;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5cca65d1f11141b49a1136898dac8226cb1ec1654c8b8846471f1e4c36bcf3fc;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6abf4748a0be2d4365fd1d9b53a44c3183015e1bdfb9a3f671eb5beed231eda1;
reg [MAX_SUM_WDTH_LONG-1: 0]                I56bb103437d88864c0ecd5bea1ab5a0313fef2b904c52adb559e19bef8f716bb;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5596d8fa3572e105a1618deba542906f0ba5acef8d7b0a48d0fe2e4eb3cf7481;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic00f466513895a54a6974af570c7bd5aba8c0ecab5612798bf512ca88f27081d;
reg [MAX_SUM_WDTH_LONG-1: 0]                I456f1fae558de9875bb1f76cfbb1840945f61ea1bce9c9bbcd0ead15d4b2803e;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7b2c627cf9d530af8ad8ebc0d3dbc53988ea1819d98b5e36e1517e21cc954782;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic61cceb25c811577024c75e771c53089a2adb9f80e6a622eb82f9d8e5bbb6c16;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id8edf0b11a998a6c5737c8877c9b203e44c777ca9ee01cce63f046a6bd375c13;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2813295228131e78d6af31808dc1d9a6f712ddc60b2629d5329dc6ee2d07c9d9;
reg [MAX_SUM_WDTH_LONG-1: 0]                I6736fca4e33cbc58b4658d91a401b558b1fbf9b3496e1830a8d7b4237d0ef125;
reg [MAX_SUM_WDTH_LONG-1: 0]                Id66c49fe8c0d931dab1b901945cc3926c6e7e3d220480a28e0099a0656241a03;
reg [MAX_SUM_WDTH_LONG-1: 0]                I1d8a87a805073dbe04ce0f76953a234bceb3e6027b2a187071b492f644843715;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ieb9ae0dc5ee16583e8d05536052b61089e8004344fa0e3fdbc88c5af5119f293;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iff41f572ab79a4cc8e83538b32d4861e88ebdd0a9ce51555053943225158c5af;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7f8fe2415810e04fccd129edfe956981aea020e4b24dd85d59991f4ef0131380;
reg [MAX_SUM_WDTH_LONG-1: 0]                I5eafefae338dc0fdd7610a7cc3093d323fbd397263d3c8b7546bf540e77d60de;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ie5d6a774e706204102b6a2d413e41c538f5e61284a19c7a47c42e356ea77d072;
reg [MAX_SUM_WDTH_LONG-1: 0]                Iab62db2e5fab6a7735067ea4afe23d7904f71c5b92219a1ea7848fa358da3cdd;
reg [MAX_SUM_WDTH_LONG-1: 0]                Icdf027acf32cc766a4ab1f19373a58cad87f74c1ca1791f66e958de6f18803ab;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib087093eca2530f923f55a4b4cddc83869730b169ab16bf26f6378b580da58f2;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ice19f7340dbb41a6b126bdae27e69b813b5d6f73ba4db6ee79715328be678511;
reg [MAX_SUM_WDTH_LONG-1: 0]                I575538bdc858fc8c843bc6b68625f1ba5fd33a904937071914caccc65f324a49;
reg [MAX_SUM_WDTH_LONG-1: 0]                Idea12ce0edfa5df65e47f6496f2a457a03907e9d62de2cb3797ec2cc6c5adf07;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib368839377e69cd28a997a22724c32efdc8820a04f9b5f93d9877bf398ec6e61;
reg [MAX_SUM_WDTH_LONG-1: 0]                I67be614a904dd4d47457ba0dc7a19b2e9f8e4231797917ef3610aea55d5ba3a8;
reg [MAX_SUM_WDTH_LONG-1: 0]                I7cd598a52037f986959ad3f02b4b2783a613170f53a7e49573c5da74f1cbf614;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ide70b17967ff52e323b4a51db51e71445ad3c5483c745b2cec2cc338e5f42f6f;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ib28a3a83a3be0baf561a184b6de18de0c4847ff892c403bb9da441f017dd5efb;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2416ae27b898336a36264980b371003c06275245f514135d0adac28d88379cf7;
reg [MAX_SUM_WDTH_LONG-1: 0]                I2d58b3296656a43e75a58883e59a576c0bf73dcd6bc28a939582be7ce0a0ffbd;
reg [MAX_SUM_WDTH_LONG-1: 0]                I3f548241255df4c4a5a8b71a4352ffad6c3e5278c73de2b1afd1a1f1f1f94684;
reg [MAX_SUM_WDTH_LONG-1: 0]                Ic3ef9d69272fb936b5ada08c6eb60ccaa6acf7b139689e5cb44e0ab76c0ee24c;

reg         [ 0:0]                   I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iea34a791d9561118f20388c1982e96791b9c45c8d09efe2e56ce981faa134d13;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4c8eece46c2e28444c6f5c37e2e5554529d6939601f8ebc810fa90d8649ed6ee;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifac89ff7eb9686dcc27ac30cf29859815ca420f6432a51b6f402333f0683a4ee;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iddab3676c92e4641120c33849987a24c0d6ce40830d17459f0535c40cc1bbce5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0136c7d988171747d52abfedc779c36c470e40bd8043ae469b0c1beea8a077ee;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id1218ca0034b49373a64117899424a661aa27c96a30d3ade1da1893fc2761be3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3e76241b601228fc46605a51baba2f1651b23918015bd484399022d97f09bd92;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iced807c14e21b11607cb94ee75e9f432fdda810c34b30a39aef1e50f8ab0e30e;
reg         [ 0:0]                   I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5ec4520bbe75dff595380b5e3dbc662e1e5193efc9e5b282d68a1bf00585f9c1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I107c1cc34b3e7fe3f69400b3e6f18745b97d257839df7315d1f12f3cb9256812;
reg         [MAX_SUM_WDTH_LONG-1:0]         If0a186df3c3fa86b38c53f061c5f78277ae3d14992d047cc5594125a73b50dd6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I16f0af67f0951998267a540be535b5431ed5e6ffd14355109089885e42fc7e38;
reg         [MAX_SUM_WDTH_LONG-1:0]         I25c23909ef7300400c6ca2484a36d95fdd5765d0ab9f816f2b7eae40b2896405;
reg         [MAX_SUM_WDTH_LONG-1:0]         I29c0576bd0d8df0a78aee42f63a6007df95d1b2cabb7424d322627654b6a0bfe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I06f14700638e4bccddacf4896cd90e26b33f1388f0a21678bc35a81fb8973e02;
reg         [MAX_SUM_WDTH_LONG-1:0]         I07a85d69a58e9ae8356b7758dc0c989aa6bcd71b408c3c7770d0e646bdd5ef2d;
reg         [ 0:0]                   Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9dcc9ad0f4591fe0ea9c5196fb457aaab567f5be24fff2b29cf4e61567811938;
reg         [MAX_SUM_WDTH_LONG-1:0]         I23c501712a70f0ada92c78d2c0704b55e90588bfea60dd5c3d6dbb0ba70ed009;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8cc4346951815e7dd3951d1975e1d4529332c497689815c86cff1a2e6bd98872;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifb944e4f518bc9bee1423b4c08427b203b24f130be8430fd7afb83bef7ba0d2d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifcb9110b05d9709662dcd3a0c985290be9f283f2b76d0a82a60b59fdfae1f116;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4359ce5cccb720df3276f0771c774342c0e7ee09f4e356283023be0a60cd1115;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac34667e98a93c9bb269f6dbe69d4148df3a55d9ea25098e7630a36b5ab58138;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c29df9d670f78350175d3c013388fbf48c167f3cfc7576f8d56186e227ee2f1;
reg         [ 0:0]                   I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3b58ebce4a4f16f7271ba1ae7dac9dc9977abd0c90030d9aba39ce0c5d604478;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0a8e687a253c1e072e5d299c180b344586ed28837bbf2b20a2a737dfbb904ce;
reg         [MAX_SUM_WDTH_LONG-1:0]         I857c867fb70f76bc0c7d09b8c34d62fe9d558eaf96766b58b776793692b63497;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3c98ae8ef287ba03079f7fd14ee83b588b02cf1b02e362e12737c93f35031230;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaea6828ee218d24373cfb8449c584b5806a1a815d7ab34c2a39d76dc3186ca3b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic34d5eef3a8c9a0ff524b6ca5d233209869368afe0266bfa94c6d159c3b4b97d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92306fea80ed98e3391ee19be59721f0ddf93aff9c5c85a1c03942ab1ddc0b7b;
reg         [MAX_SUM_WDTH_LONG-1:0]         If38b0396ad61a4a69acd171a8474d2270c09dc3cd74273589ce39f3cf9c2d9c6;
reg         [ 0:0]                   Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2aa525f826749dfac72e0a870919582cf43e69ce68dd68555201ca204fad6ee3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8e300db9fc7aee834809aaf20ac393fc3d046ffe391d61effac8eb11f7daa1c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f4e6a672481e296d10f94ea345bbe9babcdadc2e3b447be67ed1cb4c5b5b010;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id1d212084a29e275b0e589f056235a0f87097cb4fe96989ee3e2e8b44b8d14c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0df196e9a75907dc29b66b17b63677adc1d35b6b543dfb5ab01f7beedef65a95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I45edda32704ad01d8fa7f3baa6e5836bc669570d223d634ad149ab4580abd625;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3e1f15e4a1a4c0522470cf8fb86314da400e3e882c97731468b384e9d84e739;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib8ae927e56d694255bb5d70c5a6602b13e582f7ec4b06fad5c0f1c623b9bd64f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2956ab41e4cda82864182a110ce8b803793f9e0dbcfccfc439f0e473385d9746;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id5cf825b09ae8cc8c7c63eec98a9a37fd15767b0f44364dc17e6abde6293a711;
reg         [ 0:0]                   I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252;
reg         [MAX_SUM_WDTH_LONG-1:0]         I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d405f7f9d952c8a7ca9daf1fdf591b1c0108a683ef3084c8bd0a95d7ce42788;
reg         [MAX_SUM_WDTH_LONG-1:0]         I88d3389ec9d452ba7af534f1a58d6463b08369c185e66a77bfb6604e6d201916;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0d869013e0ccbc57f7bd590ccf22dafd343f209d7a547f1d24b105b31815ba18;
reg         [MAX_SUM_WDTH_LONG-1:0]         I707948c8eb9a0d646b7d61a3b86b807a4e9962d5f81c582212a6bc7fc58e3c0b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1b8ba2fabf6c4f6336045bd785ae8b52ff275740fc54346295ee42b9ba530a1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8fc3cd3e94bb31bff1119828a5ed77af969c8ae0ad80901b9e6303491db001b1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70a05485fe3663a0704c166ec4819fdd34b5b705623ae6f1c76a783449f04af6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iab0a5fa6bdfbb14163473868e4651dbf1098141c464648018316844fa71bd877;
reg         [MAX_SUM_WDTH_LONG-1:0]         If86295d92e67aea78f792b994694f74fef76cca427defd79e2368750b480156c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7c78ad362cb79bd72205c943398381fa981d5b2e995582c7b16089de4bba9b27;
reg         [ 0:0]                   I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5a70e23cd0dff70ed6ed5b227d239f56dcd214cbb2fdb0286c2e154f4e450ba4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia7ac2e243e12e18eb1233f947496d37da38950a0a2db140cd51b6e3ea075848a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c9e693d898458dc309fab7b6d2492d5b78b53f9c89ef8e7bf3f8038972b2c24;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iea4dced4cd8775da052c065ef31c3abf4aab1d0b2654d5f7e904bda36ab05ec0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5a5083c658290744b00a18aaa5fc88ff90eb17aa0c06746715f76592608ace49;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5e65da8fb9465ec0e386cc33ac36903a3dee2c59151adc9c83091591a0bf554a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1911ec0cf18a635f5d524a57281219443e1eb9eb4cb4f9b5c5f07dae014ead9f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I09c8e5480f9759a5e59d4ef582789a986f66929ee1e1cc030f6f1a716339d4d1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I29e4efa13123958a82952155cf24212b7f04fe94bf1aa7579617cabcdfd49d03;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24cce2dccb4540ed239adc5602a5cfb9a2a480bdfa780124b0d05dba8946730a;
reg         [ 0:0]                   I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icb9ad5b9e222f215f848ff5fee922a8dc526f16eba35decb2cc80395c848903c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I181f8d112163d3cd54f1842ed88acdee6575a19ff24c4702f463ec4642361196;
reg         [MAX_SUM_WDTH_LONG-1:0]         I39c3950d86099683961f34448fe235f94e87f5b7067a39abaa69732a48c0ba79;
reg         [MAX_SUM_WDTH_LONG-1:0]         I456e1a4a9412cedb175a75a2c7b65837b127c5f2478a8bad034592dc7db84079;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id5d890ac1e6399e0071d7e3ae3f3f6038b5dbbd5ac18819fbdb425cd65d23aa6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id616fa98bf8bc6050ebcaa718c98c6dcac9ed2895a71b3a0d6fc42fd71205959;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0e86f93ab7eab1ffc76fcb7a83eed533ad27ce0f06a15ccdbaeeb4c0293317f4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie517400824ee7e75e8f286ac888007dc57c24fcb6707f0b369532fa6b0a96b4a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d5e1e1c63d137b4924c9e478035c320ae319e1f2a23433b9eaf3a537db29c2a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I93f155f57d9443e4b03255cbc0718355e5bec200a58bd83eea6bc11ed564ced7;
reg         [ 0:0]                   Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e0a468c76cdf4b3b95812da2dcabdd9992c595254d9c0a02d815dbb310c302d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f6ac9fe8ed957551d29e18ea194077943be18e78174e93c0ff4f9d3dac8f657;
reg         [MAX_SUM_WDTH_LONG-1:0]         I46d9e33c21650fad18bb70da588abee2fe9735680d0c187331e081c111bdc4af;
reg         [MAX_SUM_WDTH_LONG-1:0]         I15d1b221d76c92d20200cadb2f0bb529c3b89164d7f67774ae33b2a01ea39fb4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f76b9ab604bd37a481f9327251fbb99d28272bea9f03133a4d1f97499a2b4db;
reg         [MAX_SUM_WDTH_LONG-1:0]         If9a6c15537c6ae15c785c8729b2c059a320f316c98f777dcee42050c46990ce5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10f9d40381df04200ca994a74c8a8d70730997334d739548351b8bb93dc29a53;
reg         [MAX_SUM_WDTH_LONG-1:0]         I11b57b318e1a6ffe46a449f5031d9517c7b51452160307f7c0c414cbce227277;
reg         [ 0:0]                   Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7b41563150c1630c478200a5a0a08a7809a1ae2d161450e63f10f4629308ba45;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9e477ebbbe435cede26f2d18e939f81f8da88b0089026282010e0f60e8d3e89a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib2254e933b3358a2febe2ee78bfa00d03502945608b8eb00f8b921077315df0e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92aa5d178a20d871c5226ec40b3c94942f20c06ab5351b9f0bd08586022f76b8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9261ce4479f81cbaad6fbb8ee9c872d9dfdab45875f0af6c01c479990686fffd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7def5551ef03ec4cae6129877ec5f900d6d7edbc6fc66f3f80de9a23b31adadf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9e2c2192b5d360a53c35daad843eb9d5e18e850305732dac35c9213a45ca5d05;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iecda880e0e0336e9564a1eefd20e2d22e0ee56f103a90a56427a0af52069511f;
reg         [ 0:0]                   I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica0e4cafeb0b7c9e6caff0f66b45625890be48216b4a25b0fd582a72e2def407;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibdbea6826ae5ea65408f48eac06e1542cd2b3b0e1a4bbeba724c85ee552f1d6b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I67619c07a6d53459465f2d77929930804aae53cbb52a97de1d849e532d9ce5cb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I555422dd30763e140e02b9b6385eec9ea18ed35842a4eb56f68f861556d50adb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib6b064fc5e6213c920e8d2207427c6c27622bfccce85f662b0bb2e677990272e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e5e6e223f3acc5d6f776796e0be8f4806d5355cbe795331b0ef20ad3e12abe9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1a7d235bf70814393dfca5c8eaa078813b915fa814648adc0a6b2d72e24d1d52;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4536ef4b6318344733197809b7d7c05af0bdcfb40818c16bbd525cfe55e1eb81;
reg         [ 0:0]                   I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic4910d74bc015f92940dfd059f327ed96a95ab01a170d3d00bb266061a7a157d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9022439743896e55957c8ec574d3e2e14f88e6baf4b65c4126cb39e589a92da3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I52412770a9e85565ac24e94df63da66b761a5e54ec1bc8c5c8b07b621a33a164;
reg         [MAX_SUM_WDTH_LONG-1:0]         I43c4705413499cb45c94379264ecec3fbf0bcf83aaaaf0110c9f13309682d21a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I815e9a6b98dc1542b276704eb99ea559b4b34a16131b14fe631575d5fdf64e66;
reg         [MAX_SUM_WDTH_LONG-1:0]         I462a0b49cb7c2a4940d2befa6f37a5c2aaed3a81d20ff47d528b821f8f9dd245;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5f1a06fb6eaeb2fa30f132d4fbbf98080868dbcc827b35e3a3a75945cfa97ebc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie6a253c0afa00e08e20896c2d4c77582cd8c24ba00c3363830f057a7f321eb05;
reg         [ 0:0]                   I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1aa2c1de85f2c5fc04250c2fc277af4c7fa7072d9c7946dc8f6f240dcfa87c2e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I61539a1a79c4785262e8d239fd7e9f5d8e7f8fee2526fe7b4057795b6e5a657b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iacd51e59a644b3ee8d3b73b5c6e6b6b89586e869487aed8e8c3c6b86c5e82135;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3ad491fb952d351e2ca1c3b3994976b3dd273509d86e95b341f2b609175cba9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibf8e7c032bde3ca68321b7cbc2e86bfb0352bd5c21d5da458b3f98d751b3f504;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d9675ed29efda87fa20ed542d67c88fb1782698b8879fc28e908d27377c939e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6292a3c00e5ada17538f4bf8df9a28541f5d080a806e8104c49a89d94abe9ffc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I96289ce0db8e685e23fe7fc2b1a700a4cc2d1938225bf444c320d7194f1ae820;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1e20a0a29f77c9e1e9f5d4b6938ea3dbc0fd30eff663b54ca2a3e255b3075c9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id5110d84643f22616230397f50ceaf2f51e6c46fb596eea856ad3f29c4385149;
reg         [ 0:0]                   Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10b08e5e9575d53b3c52e32527e38bca0fad4f0ed25bddf20bfd1d454ef836e5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9473ca20629c79a46dd6db402744d58ce1ad19d823d0f3f9ff6988c22f02dc8c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I26657dbc109dc227769ffb9fe0418b97e1407634c4cb9d19d48337861333cf76;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0867129ec512051e4846e12f23bb824b363561c6e2511511bddad44a934a9299;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaa9d2267657be14e58cfc2369f00ccccf2d09b8711e2325c11eb099296260046;
reg         [MAX_SUM_WDTH_LONG-1:0]         I08db08fceae6dac922ddb30dc8c5d2ad75fbd5b6aa2f24fb0b42216c988e8881;
reg         [MAX_SUM_WDTH_LONG-1:0]         I835263edaf6c3692cc0dbdcd536e403006ebb5becaf77abeac432c98f2a2e261;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic6522502026653a983fabdc7a97f3a61c6478884ceb2dbe7a61669f09dec40ad;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia9b3853d7376f2b3ff71063cab059c2e5b2b888b4bdd3ddf38c5b207fe5978cf;
reg         [MAX_SUM_WDTH_LONG-1:0]         If869318b9b2eea76cb0f28203ca8bca23b5493b21f9dbf176915a73fa7383cc8;
reg         [ 0:0]                   I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f1a7cbe72daa5437fa96abc25ece5bb43cf13aa018be3537e107fad506f28fb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iffca3b5121937820dcc59668b1027b5276cc746cc65b3c8cee5adf9be0e4f33d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0ca8ee6c12c754f4b5fbbbc35b5edf976cd2f3a819a967d4f7808544e759058b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I09701bbd76150af027015cfe8cc976f8bea0834c8b3cb443f11baef2e0799636;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7225c329ff4c63f38d638c6647b92bb12ee5063dfd2f1bfcabf0272878cff77;
reg         [MAX_SUM_WDTH_LONG-1:0]         I78da05b970dd2ce30b2503f93922c4281e5daa812cb0aa255120e75ad946cb4d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a363fd35ab7009f60fb2c4f96f61326c370defc1103deedea40bf0d0159256f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I806f8a32e68e72b07ae9fdb26d41ac1a42bdb0fd4ffcdee68fffd430b0b007a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70c5e2d6271591901678b8f0e488d737b3cb603b8b8e448024cc9d7e0deba259;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3546a9ead1e1b810503b6521bb2c34151dcce36548225099755e87bd323b21df;
reg         [ 0:0]                   Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5466c771c60a3618aa4866c2b07d5b586e7d7c70934a747a04273c3367ae8abe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I83d8a4e44b0c8c27a4ff0338985fea545759f3660b941608878feff2c4208c82;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id4e193d0a39e2ff4ab10d577523c3d264b54fa0a698b4ed0aecb5ddf075a4acc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I779445414027b5e440b1075ad92e9c743a919e539757a4305d3985b57cf1ea50;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9cf43907a8c090249537efb3105ef878ec38cf189b1848dda10fa0934cf6f0c7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I946b706dbb3722bc8069bc60a27d6525a81955d0b22d8c06d5730b117bd8050c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifd3de8ffeb5f4768dce5d08e6e10e4afda032d8e4ad7e88f63c50adfbe81afbe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2325959aa541dcc2298076e643b12a8a9656b31c28607ec3204bcb786729b88b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib8801db7c3d797fee2cf63037daafac592616e4a958094ac2d7a85bad398c437;
reg         [MAX_SUM_WDTH_LONG-1:0]         I64e64024cc00dbd7a3a826c0f9d82dacd15415b344d86bda10ed4d0142fd592d;
reg         [ 0:0]                   Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I658d4c16a7bd3c6d82219fa10195aa78c15698af2fa5f3bbde967e29fb4fa8db;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2e7b8e10124f284adebc18b9edb14644f54d024c862e86b76f5d4b04aa2bbc7f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1a054e117ce979becaab2b848f8b5874cef5611170ed854e8536c94d310b3ba7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic15c7d8a56833e13814c297cf7982b48a42a0d89cd37c0a67ba3c3528546c240;
reg         [ 0:0]                   I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I79f4cc267149652c039a1084e89dec27f52317ffdd1f4e813053380c7f38982a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7b69470ac56b2ee8391293d6203e4fb6b7a3a605f38fc684f2eb1ff49faaf1fd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a670a21ee5fcfc5f08786bd903f1da0c55661633e25495ee189a3dd55244f0f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cb1d387b00274ba18c42d1329f0bbdd5b95e586049a8230d94772d73597b47e;
reg         [ 0:0]                   I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3f002730cfc58d827800579d570d0433b30d2f387e44b0641fd4004f52c01c27;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife74c161a8f2dcf48e3a3b07d65523789eb2aeb2cc2aaaad88cfd91683069b6c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9bb3d89cfaf62aa40cae73b77d1a1ac2999465104de1d7c188918432e1a17c80;
reg         [MAX_SUM_WDTH_LONG-1:0]         I82aaadd76fa8b5e7bd489cced1bc3b825f8e281accbc496474db7c4ea4d1e1e2;
reg         [ 0:0]                   I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804;
reg         [MAX_SUM_WDTH_LONG-1:0]         I790d57f4f5730ea4166cba282bf1350f040ad2bbdb8863311b0f753991858960;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f9bc5d4b3aedfd4e192fdf7774ca874dd2973d41203f33deb2dfee1f3d5eb90;
reg         [MAX_SUM_WDTH_LONG-1:0]         I219aa384cadf0adcf51cc6828ca3dd9781775e7e7986955e6dd5074ae6bf0887;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia682b7cd027239465bf24461fc4d88457ca84c607032663699d76d58992265e7;
reg         [ 0:0]                   Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie226e795a9a67a0d9984f30a164ecd2aa0692100a18a77337c2efae4395ff952;
reg         [MAX_SUM_WDTH_LONG-1:0]         I393c6e437a6f283fdacba0192edc09f7a8882ce8c6516d0284b10a6ed2a43a27;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8ed39202419d4320b8d1fd945da1efe6befa43abd55b3ad1c7917b0587cc3950;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia66d77f2baa846741b30c7f9b8d0f770d488b658b6d2ce6c265f8de5dcdc3af9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I939a2a515cd6383018b9d98f9c3b748c75abd1beaa52e26c273eaed8978e9372;
reg         [MAX_SUM_WDTH_LONG-1:0]         I66a18b0e3441516bc7212f5564b7d2e079b7a73bbc481c67c4b357fa3a766f4f;
reg         [ 0:0]                   Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6e91dbdb1c31ffd16d890119d91969004497b13d180320f54a27b001b8814f3f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0b0cb7147d168ab10e2a8d7c9c839e509d8e967d163eb11c4afa8738c06a266;
reg         [MAX_SUM_WDTH_LONG-1:0]         I54327a37a56f54ad389401b3e67be69eb0a6ace8d0f5ef507f5edfec4cb60f33;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id6ff08336ff69aeb7c86ff3c649c59079585a9117b8366ff1776938c76509345;
reg         [MAX_SUM_WDTH_LONG-1:0]         I74cae7d7ceb41afef5f215f9e99e5ea1ee0d38efaa91800a240a26b49dec44a2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I73d3f78f124fc07e4dec71f536f875a26946b68478ccd830fe94b24d6dc73f0f;
reg         [ 0:0]                   Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0dbbf32467809debc31db520a1d652a39c6f32927d5fe8e7bd87a0ccaf5dcbdc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4bd4faaa74b900831991b7a4ce8511a5bb45c1ba413ef0d2516ae105cc00c740;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7252a8cf8ccfbfa3d707c9f2ff6b0edab9675a6e54f6e03a8cd7f06f77d2eef0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8534ec2afd654d78899e86e2eac05d7f62677fc213d962a50b1fb5d853c5b966;
reg         [MAX_SUM_WDTH_LONG-1:0]         I07de1ee4eb883d98b9baf6d4b08768203be9277a5780b0b713b054c67b6e9362;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2dbb829ee8781d23865b9bfc192543f10ab2839afd1a8f8211259f1248d89f28;
reg         [ 0:0]                   Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1c85612795fc824409767448d6770bcca93caf10fc2cd8659a98eb808c878444;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib2c9dc402fbacb1f26f72f8b1f1578f70d7a69d30751d4e4661514a819b1a974;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9d10906535c09c58cb10aaa6c3ba524ec6f2bf3bbe58da21edf42dc791662b04;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2cc9acaff65bd5636a9def070cb29149ff8834daa39d18594d09d6156003739b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I478e7d5b826a54848c89bdf12a8fa4b7ca31e387d033563784c60c493cc633f0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ied5920560e9017a8c035f2d6b019f9abc3c8ac6dcf213cd3e422f92510ff38fc;
reg         [ 0:0]                   If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115;
reg         [MAX_SUM_WDTH_LONG-1:0]         I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I50780605e408ffc7501e94d92284899a4878c5721680a9d734ef276a4c9974e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibf3bba34d932e08687d92505ae09625c8c1cfa5c24d3d52273050b8186ecafce;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5af920c58542851ac5891f1f1dce969c57e1e7cd12a302a68528c7c02c86a524;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8559dbc457ce562bb8447f1227ae0c59f2566cdd93fd9051488863bb3e4aa462;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3aee441136da868b3fc343e6eb88d4a48a636677bf1188261315fff1c8898690;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1aa8aad0f4f034c292c7799a12e5f7887263752b5f11909fb73b32db7c6d7263;
reg         [ 0:0]                   I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I559ba5b3899cbbfda28e2b04083c4958d942ab0a8577e5e7b9dabc58053b7f6c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icb53fd5ff0cc1bb11f4efa51be8b18e0455037e4718b955718ffdf5d6bd24dcc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee6c6b7151a6d52632c5dd250c0fd5c866ed5e07c96d8ba7ed0fbfb13b5cc9ae;
reg         [MAX_SUM_WDTH_LONG-1:0]         I54cea20aecb1a113601e099b4a28a9582e143bf7b257df21a059c2c561056024;
reg         [MAX_SUM_WDTH_LONG-1:0]         I127ecbb26b8b54be69afacba0c7c900d1eadb8907e3337013e771e8afd15b8ec;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib655fac982e2ba3b34f9be933b8da91c7416d2add55a9225d8354e85b51c66d6;
reg         [ 0:0]                   Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26;
reg         [MAX_SUM_WDTH_LONG-1:0]         I066453fa3220e314882976bf9b0e935d3cd7f5233141a89a6fb00390d245ed9c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc27708504fa373a81980a39fe27a732fe8ed4d3e67838b787c8d633cd1134f9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9dbb69baeb72fc989c784ef8b69a50b8acd0c076fbd3aea250967efda14c7ff3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3027ef5a77a2956cd097cebac4348dffc636fa06b156a08dd403916fdf42d957;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia0f10f5c6d9dc1cbb77556836ef659a542681ea3f0bd54d0edbb2259e14e6c0a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic81c2a6ad2dd6d624ab25855269124b464c2d5dfa31e41fac639a888994a2ea6;
reg         [ 0:0]                   Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifd84bbe3c8b82cd5fcde5db6c40190c17411a69c9502007d0392efb1b0507c87;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4ae6345c74a23a9713c9efd40683df95cb7d8f18163ecc526a0188b17f0ff54c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iccfe7f8fc79fb4b135af4cf2a698e9ef2614e7d01d137304a0b51502ba34a79e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id99854c623c0f1fca0e55e9b6125fbad754c4311497cac1ea4af1471342b7f15;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iffbb3bf56ca327afb4dd8826363aa655718ef15e14e5a6b9e55664d0cfc76738;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6f62760d6931ff9476617433db3f760557bf58b267224286d0f1f38777f1c19d;
reg         [ 0:0]                   Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99;
reg         [MAX_SUM_WDTH_LONG-1:0]         If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib5197b3ded0d4c6cfea1aa9572fc7eb7b3e0afc3b5afff40dc48c2fc2d06ee81;
reg         [MAX_SUM_WDTH_LONG-1:0]         I421cb52dd669a636801d3709f62f6570b289aecb322b1afd2ffdcbcb5f1377a7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44643d87119bfc715397cbbd514f7a75934db3d6fb8308d0874dad36e6ff0969;
reg         [MAX_SUM_WDTH_LONG-1:0]         I016081dfe95a2bab40513c2f55287a990f0b79588fe1b8286174ded6b93bc278;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib70f45a310ffb94185cae456609a25620a223187f0c4c3a9f8c5c645054ebb96;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4e13170eb723e9bca567d19c25b56d782987da1f75c5a54ab26d0b1538f779e9;
reg         [ 0:0]                   Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaabe2ac34f3411032dac139922cf9783f86937c5d525c8730c8ccdb257f94f2d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaa84c2b3b1d95fcb9ff86fcc68a6049f2c0c0c34101bf5bdecbb6d72bee244df;
reg         [MAX_SUM_WDTH_LONG-1:0]         I79cc31e6c010fa8eb54cd33d70364720a3290ac19ba06f27ba05b1bdf24d6314;
reg         [MAX_SUM_WDTH_LONG-1:0]         I045079845680e722358f1a61dfed5b3758b7d491231d08f6f6e674dea560885c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I43e364076c55650d4376369dd211f84289220dbda754e9f3475b5d1310d66659;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0b9df0d909722adcf9aa8ee430e388b6f201b7f66e12c3cf72b4751fd4249b6a;
reg         [ 0:0]                   Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iec9a71f06ec498907631c7b9709bc6461d2b77efe8493e4815501c56083727ec;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibe52a5b5286c8d781c590bc26cd000c66c7ab759989f65c747574503e47867f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I55d30fbaca443183b73eb12a611cece679d3b08098711ee7a74767fdc25d8ade;
reg         [MAX_SUM_WDTH_LONG-1:0]         If20f8ce49f49f296f4747ef4388ed862862070b059bc482233542b99c18d7373;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac1ca36a507d9c411a740df9fea1934e7d8d64695834a37eecb2cde9d03a9204;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id62572be7c49640d6256571053ec24877befc584f4518c67f81dddd33afe02ee;
reg         [ 0:0]                   I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25;
reg         [MAX_SUM_WDTH_LONG-1:0]         I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8c5856de3a047c2d8cd91175dd65f574230329e0a98bb369bc2f1efde176aef5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic3358b7d409c989b0359b4768845d172ff09d2c61bf9d17e51d0323a347dbbf5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4bae23c126c76b438684a2e720dd190ada836cd8aff3a9f217f8fc93dcb5941b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1c6046860b8c1def57621b5c2fbdeb57b6bb9de1195675a875a1a028ea2cf881;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6f58751fe0a0b377048b39ff9ed4d073ab5205a2ec8c36b93cf8adb44ad81d4f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia43a684b6db0d7a69334ee35b6e06b35546b75cb48143fe9e7b54773b8c0341e;
reg         [ 0:0]                   I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0d2a131e78e3e0c36dcc971e7ff76990cf1d19e2d90d373db2a81750458bfcc0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a190a23ac0ecbec7ef85c968ae10b90f7f0d9f5400aeb74109b51caf4caa2e0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I97576b987f44843040444751f4b37c3b5974dfe60b4015dbac8adb962635ed1e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib6bcf064fff2ac3dac1a636d200459bce8d2240757710aebf6f5ff055ba808b8;
reg         [ 0:0]                   Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iad4f04d003ec15a32b36b0741a3fc3ee341e7d02d9b7d495d63e26d02d5f278c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I71245defdd1d5a15a8c64a0c1bc585fb3a5acc2f6427408b4c526faf77e5668d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9ce7dc815e30f744716169eabc1fd21116601a539776481e8f75ee17262c7fed;
reg         [MAX_SUM_WDTH_LONG-1:0]         I19dd506a7468a183410e0bae3025af7af57306a264f0043f2f9a0635a3a5cb5e;
reg         [ 0:0]                   Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idfc570f0db8ee7ca88a35b7c9ffc2306308ecc26877a75c31ccc436f1e9bdcc9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4e3b7e54b82af833886fdc3ffcb335189bfd516a758fd9fe96a0f4dbb919ed11;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92b84a136bf952296131c7162a68c4215e69d2cabfd345b29ac1c0bf22585921;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7203b0e25219256938283b8d39adec66610804f8024a63dd2bad2ca9e9e01a10;
reg         [ 0:0]                   I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb;
reg         [MAX_SUM_WDTH_LONG-1:0]         If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8d5085a98240b391006667ecdde09a3735f02bebf47c3ae2e3f4983183111e5e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I793fbfdab6a3b0b8951196e0a8a76d4844094cb64802cd8d50bc2b7ffbb0d937;
reg         [MAX_SUM_WDTH_LONG-1:0]         I62a85956a9fd75b6c1d7f93f5472394fc8d0413995f21a8eab042ec0268e63fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I64a047649ca6b299cf603e326db494b30d1eb35725319f172957fa38f00150ca;
reg         [ 0:0]                   I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1da8e393ff7564ba162ca784da6731a8632fc4f6b34d907a52185a8b6a59a2d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1c9e95f283090d633d1a8deac1211672e46383b70ec08ba60820f0096fea280;
reg         [MAX_SUM_WDTH_LONG-1:0]         I066d165e686a647ec05e381773c53d7bd83320b8abd57693dc5dae88a01fd8b6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iba95ca83f9a8247abda33f9ae9bafedf0b26e6616d5bfbfd78b02637f6120c00;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie4936469b1efc82d537631d9126581b917e052838c19db1f8fb4512d7352f6d6;
reg         [ 0:0]                   Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7dae66792f1ba5fc8ff7d7541e3c9fdc44b001e3103715d98c57ddbd35686d37;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idb01042afb3fe35b5df33f4a990e8d512975c238b7dc146f8c60fe42178a232e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I81b03c11c47391653037bfc546e4abce946e244fe10d6d3746006dbecc9e6dc9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44dc65b9b972b02070e5bac23ee64e568adb39d61d0f3ddbac27ad0abf453fde;
reg         [MAX_SUM_WDTH_LONG-1:0]         I53ea37aef026e5dc7e966fab827b86b9a180b1c64d53801e51d7f2c66c729cf1;
reg         [ 0:0]                   I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7147ae9d3a1f4fda281c89a81e01b66d9db82d9e8f609e313a374cd5aaadd687;
reg         [MAX_SUM_WDTH_LONG-1:0]         I550a8278e2a551834175e8275532965c7204bd2f4d021e0c087eedd5a3fbef93;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5b5d22613b68a9bad72ca89d654b0a7f9d21914b3d596af6ef7de32b98e66e9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I749908d9a05ab10736825bc8f1db4b879d94c4cdb920daa9aec231b8b2a26dbd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id85f8d61522c12b51ada0a5c2f8c492d1a72c4d5ef88c99b2b5ca0c8a885aed8;
reg         [ 0:0]                   I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a627bb2c8162e911b06414d590ddfb19a4b1b84d0af6c65f451bcb6cb4978e1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica888e39630b6f3eb799326d4046056ef55883125634fcbdf6c36133ba571b52;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e0846788926a4b2a76f01957b236d542f43fb90aafc16a952cc502d83f31cd9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I85ff081ed2d76aa65ad78d86b7804ea0f8822cd35f8b14612104ec232184c5fb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2f5cf926d3a647e02544e7839c6e999a0798aa5c810a6031433237932e96602e;
reg         [ 0:0]                   I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5f43984a17fec9b995aac537cfed942b8c61fcb134ba29fc82a41db44d46c820;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a97a4296eda318163fa6fe4417e08ad1963bb488a6bac31f3b3b6af9e7ab213;
reg         [MAX_SUM_WDTH_LONG-1:0]         I439b2964d8e94fafab2d3cd19e72728d4e763624497e8f44e10a8be796d87a31;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6476bbdf545c28c272dffa9640a8a640802826f625e7963386bd6b5309fb3588;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie4122a78fa86e3e8cc54ebd8e3d1433ab29af18f8d6683a4eceefb4108faeb0a;
reg         [ 0:0]                   Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1de838959290a975e08aae4a25944f707aa1ed044defb47058acac42075cb7ac;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5175fc2784d1f63752e69a808f26af8fddf78fb8ab1a897fbda883f056debdb3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4056a6197e1723e278afa54ba45c2bcaa2766665f2d405d7f11217213f4af9bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I913a4d3bc811c985c378f0c3ceb8cc0d03637df817266b2a5009fe4e96362cc8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I594b5684b4713ef793ee902ece02cf083e909b95354d67c351748b2b1ee2599d;
reg         [ 0:0]                   I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936;
reg         [MAX_SUM_WDTH_LONG-1:0]         I84f3d2170c4ac381738a10ae95bcb1a102d86d6c96bc9c0eef4a682237cc96fa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I386f960be90b491237062d67c19264f36bff56381c3264cd7942a395bba04e72;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id25989c592a2848f8881f1ea00c42faaaf70c1571f602311ff1bad99c7cd151c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie224e49b46cb25ecb4a8126eaf672bb12181bb28cb1e7cec7eccc94403d72b09;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4e51e76c5c70e114f648c8715d629503228ea3845a66122c7da381e67e805912;
reg         [ 0:0]                   I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0261480422708e60435782d1ca5012495ec5345a3decbbc9815bbdc2ac374b42;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4c4a1c399094746d92937b66958c6695428a7963aa82fef3c8cad424289612c5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic8f4e82cc2d1d643e87ce3d6da690336e97a779fb6fec983608492c39054b09b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ecbc44de1811b06b96aedafb731823325898269d3f4d57a164b63cede9bee6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib23e10fc2319b575483f38a9a75d9a8b55d394fe0d356c89478844a16504cfe5;
reg         [ 0:0]                   I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5e6f080405681748ecd82a9b555257d553cc1dfcde4ac5f470bf1d282086b3d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia50f5ef4c28fc1650d46ad29de2ca34971e271c9248f06f24953db1d9f767faf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3bd09d09f4fc3bb758f3c1f36925e9f0504fa342b2d80ee031e4c9665fd4ea90;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie6ffb8ef3481ecbbf20e52ff7d04f51a024049190a3aa838c398f71bf1862115;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a6117b4c4c11077b066e21819d7bc164de5f4060d1c12f57a9751afbc6fa59f;
reg         [ 0:0]                   I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I96bf467638c2ab6963f57f29caf1efcda6250dad69e87b2833c6d094112a6731;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6a9adf149ec3e5da62c6f86b4263910048b212f13e52e6b680386feaab5126f1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie8947b0e08f05ed4ed4888467fd64bbdacfd30fcadb77185a75e53a60bb78877;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a66315056f6207395e960b11c230998d50db5a65f8414eda3a59ad04784a571;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0f1690027b69262a948ece04cb1de6d4d7a358e60caa676760118364938210c9;
reg         [ 0:0]                   I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I97771793dd6517655733e9ced45e7daf0a11abb8377c42ad9710c40651558e6c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ieac377a04bf039ea4d773d3e6e336e32f2cf37f375d79bf0867b5e7b7b269254;
reg         [MAX_SUM_WDTH_LONG-1:0]         I887deded16218f24dd4ccc29a870e96b43b256ee62e0bfc6ff19c01fbe5b1ddf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2b9966a73da68558c67e6cfe373b58865794a87b39dec4065056da2258197341;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6ac7d8576312302a7dba1bea496c3dd7b20faa3bbc8972a0e231f4e5ae3df8af;
reg         [ 0:0]                   Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5290a020c4e8d95084bdead6e37865decf5c9f5410048322c1f73361bbb49ef5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia2fc1b624f958681d009ec01ed83d41c0e26c3c16ab0fe1e3ec4db7d0988255c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I33974096440683b354b7725f26284e9c76a7d5722885b7ad9adf8630ccfacc79;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8de6b3b4abe26905e4adae37762f35b8d1742281e0d0c5ba45a0531020a073f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5011d2823a3b17fd74435029ee1469e792ab5a74fddd2d617c4d21b401781c0;
reg         [ 0:0]                   I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib4de4fcc7d35169a59e36a3af71a7832f967b7ae3c530c07cad1585784f7edcc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ica1376e18c562fa0863404b998af3c4e320f52008e7287b730de37fdb58e2dc0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia6251a913ec7fd4390c5330bbc9f4a983a37c274495a16d05dc96501050eac19;
reg         [MAX_SUM_WDTH_LONG-1:0]         If46b3417b1f584a8866028e97e62402cf411792fdddb34faad96f0808ceb6d89;
reg         [ 0:0]                   I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54;
reg         [MAX_SUM_WDTH_LONG-1:0]         I68dd3296bad4509893f3569f8b4e0539af4364b95ceefc0f95e3dffa5b90ac1d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e32c30199d506efaf13a091029320249c5a524f32b0e55deacea536599a92e9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I97f44fd7abe7a43044027a60cc8b9e88d1c474e613b30fb092267b7d8e0d0748;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic9b7ae6f6993eeda2a7297af8e3a9301da5055c1031f82fd99451e607ef70738;
reg         [ 0:0]                   I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idd55fba0f9374647ac6e708497c4118c4493602ebe8f342e6ffa87b496fb92d8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I94a0208aa6cc55e3ff0c47d436cdbcccce15887177af919270ddfe9096a0a7fa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iff2621e7d8b4bb5de9b649f5424e482b9dd4f01bb7c5609ce8eb76766e301d6f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8f5b316fa91d4e39b9eb94d7d051c81e4e95dfa2a2761af7970ff04e6ad1056e;
reg         [ 0:0]                   I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cbe0e864523810adb559c85aeda0f79a1dd57f819e9904d4635023fa1a689a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I03c8aad8e9fa3cbae4ea5779a2db031113b6bf72ab3df44995217640c7f52cb2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9f9f7fe2510dda62df0c857cb4ae9430a8c435a64bf84a6d94848e53bea684f0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie596b7fb4376d234eeb9946c5e2d5439cb738fe881235324c8d333cf0283adf2;
reg         [ 0:0]                   I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44d6eda047420415765497d6523a69b8ba7903ba7a76658dbd8f84d079bdc416;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8677eb1f6f7ce797b6e713913227fa9a6d2953074c6b4208dcd3a04a1769b3be;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1df660831634377e177514ff041dca7c173c608c37c0dec5233ed65899fae519;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia5900c9e78693f74b25f0c17c8dd79a78f7187cd79892df701f93314cc71963b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie8edff06c26702bf20142c7cb6eb605bfd52076483bbd6e941fddcf87518f184;
reg         [ 0:0]                   I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id858a113ed0d9d3e0b3b3041add0654aa217c3781cdcfc32a081422edf6c94a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I63688514e288f5d828f22310d609beb495c809315db245d6cb783e02d21aa354;
reg         [MAX_SUM_WDTH_LONG-1:0]         I402c6bd3528da160ede7f8c92d97a0c27835b1fd267e14fb8d92706f13719570;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icfdc65f513f27d474c48d7fe42ed9134e668a9b706d011dad7025214c61c5c6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I59cbaf9b106eecde3385e8d646545284791f53e64fef5d89e72699fdf9d66786;
reg         [ 0:0]                   I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528;
reg         [MAX_SUM_WDTH_LONG-1:0]         I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28;
reg         [MAX_SUM_WDTH_LONG-1:0]         I80b1e51f33d8c209746c92f8e1d059c87bff5b4f169bf9304bdd30f96c5b1d8d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic36894855099edb8618f29e72154ee32f3f130987bdcd435cde2f87ba39aaf0a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I676598186f1a742ac68bd8a533c205b9b5cc6aa540b0519a995388d5db421574;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2212dc39f8bda130c6782e104418cbfea3d2089b3d0fc700e8acbebf1fd9d296;
reg         [MAX_SUM_WDTH_LONG-1:0]         I371e726b1f426a879388bc0d28dba55143a4674655374dd183793fa42b8bb67b;
reg         [ 0:0]                   Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie412b52497a49cb060e42e15db8793b4af98294d202c14543413a6e30de8fe09;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie3226e6cc2a926d44860fbdba32984e2c3a007c1dbc172c3765cecc6bf4efba6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7be3e45435a982ec33d6b56aef2c5a81f233859f8312e4b328c0a9e8c11b5822;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5363dc622b9c481283f71015f9fb2a340bf5f440344dcabd8adb4961a89bb36e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I194ca19f61c5d4e4df1e7cb9398ea02166bb2f231546f23d151370c7bd533425;
reg         [ 0:0]                   I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iabf25360f3e96668f6ed500de6bde88342e176aa39205579d171adff86c5acf5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I67a8f91668c29b02c6638bc4cfb4d99364679a1e19ae54b6928adccda64333c0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idd22bb99613e9b5b2120390d00fc41e25227523bc60e6d281f9ab3e0d9eae0a4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3234917db6bb05ba543d97c095bcbf419df98d4fc7a64899f340864d7965708c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I111227fa4bd1705699775e2dab468800630a0faca805bac5a9bc6d39e3e0c721;
reg         [ 0:0]                   I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56;
reg         [MAX_SUM_WDTH_LONG-1:0]         If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17f10c5cfeb0d1c9030ca3b64a6cccc65dc578fda6a627ac3d0d0c03aea66041;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d431ffdead0e5f6add0bec3d162c7045953e597d33fde53a111f929f278b8d6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I57b332bb53fbdc45a8274e8a6838c2d3722677a6b560c2379ab92e225f4aa64a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ae1dc3a3f40ad8a03dac4c2c2b657d83c3522992ba57052e238fbc8b836af26;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0980470783afadbf12692805326a5b81079ba76f1c19e80bc7f0a30e73a5294b;
reg         [ 0:0]                   I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4;
reg         [MAX_SUM_WDTH_LONG-1:0]         If55dc3c3f903107602154e84ff4739788ba44ad35a05bdd8e2987d02dbfb165a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6aee7f7827cffd92b9148e455718c252b04105a64b8d9c60ccab52ee1ec08e31;
reg         [MAX_SUM_WDTH_LONG-1:0]         I619b017a1e80738f224764b9062ff6a3b9f2321eeb8fec5ec95573033d33a9af;
reg         [MAX_SUM_WDTH_LONG-1:0]         I812fbc992824cb1e29cc2c40421e63ca06fb97c9d9e40094473cacafea5f0e0c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I925edaebfbe72a77427ff9387ca2b955f2eaf2c3b6d76bc14f6acb37b4f98720;
reg         [ 0:0]                   Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5842c1f6bd94143ce3217369de2df9d5f2035e55dbc619313375adc7bd97f727;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2af5890840cbc6f131cf8cca27929dc20330f4248a5d7b5071de85d941bdf2e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I01542998e0af4239394cf341547e6dc36ea36f77aa1f2b371a6f915e99846f20;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1ac783cfcbbcb2dd26bb3b2a766481a364b520ff970a1ae49f52048c0cbc228b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5ab65b455c544d54467f0a12db6ff74521cebe6cf47f583a02508f73674f5bca;
reg         [ 0:0]                   Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681;
reg         [MAX_SUM_WDTH_LONG-1:0]         I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id3731847bbab8d64f89de08c1fd5a8a089de6eafc93e0a079bb7e0a990d3a010;
reg         [MAX_SUM_WDTH_LONG-1:0]         I519df6e33d8ef22d52e32b8119be2aaec1f50dbccc5d79dbae0f55ceb6cb8f18;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9b4f99332934a592b74d60329e811e336cbc4f6af94e1e7585e47c8096b05b3e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I513af0998e26ce841c280947d55c670808280391fcd874412081722d9a9915c7;
reg         [ 0:0]                   I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iea8434e90fef04642cfc1cbec886240547c066665e40258a1412ba69225faef5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4fbe4e6bbc2d22f919e4642a3f6e950358f3ad9c6ee0d7997ed355969a8023b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I83d1b40ee8296b6a8bbf02a87c6f077c2230f2e8875c679642386b74c055dc49;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia70f5a20618894e74f792df1afb11ebd1e590400cae3cb09cd1754416a26bd07;
reg         [ 0:0]                   I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8b2a2914ad57445d7e6409d706a2d5c9cdd01b8f7163d153c1647304ed71c1c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibdb714449c61293321fdff34d19ff92c2a66cd677739a387bfbbfeb482a17aa9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6640a4310bb1a9135eff3995cda6d740dfb307d44c62603190f7cbfbfe285718;
reg         [MAX_SUM_WDTH_LONG-1:0]         I13d152d9c14bf7e9d0d71bde2846f80bafd4553400bccebd37d850034d62514a;
reg         [ 0:0]                   I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3c0e2c1dc0aee993679368343156a72f56d55c38911596cd28c13fdbc68ebe53;
reg         [MAX_SUM_WDTH_LONG-1:0]         I76208cd61a51a2330f9d46b67e0b036db6de794a34a380a75ca6f60439344546;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib95f8920a685d0da3fc07ac7ff3a19ee1fd5fc65dc4b6db141a709668c2d579a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie5269d77c7963028196afc5b429c121674eb881ef85f0c30e06bf3e0b5b3a7cd;
reg         [ 0:0]                   I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ied5144deb00adc8fdbd1024c051f87a6725bd5211f5d24ed9d965ac7bf0dbdab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I604e5b545ac6c440263889210560ae82bc9dc0f3717b456ea8844cdad1813c2a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie802b6bc444bb7d279d93b810491f7dd483ceaa3c122368578579700a1723669;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17e1e63cdaf581226fb06f909c0c75f2ceeaf45e1ebe93127d22a0ee6ca7e8b9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib106ae5d2b37f2048bc3c493b80c76048d8b5c4e1ebedf0cdcc6bf20958f39e9;
reg         [ 0:0]                   I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6da36192889d17f86e9b385d553a116e1315dd88657c56f92f4603cb75e6de4f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I48595b1f5633b6439ad79fc3c53fa5da509c15abaa66b7b6aae7fe56e8b560ac;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7ff33f6abb8c5ed6800e5c1c58b974df6d1359987f819291202ff2413494aaaa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I914341a688ccdf40369a1abe1fe5bf72b3d5ddd306f81d3364e2ed4e03970149;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3e201da437cb62d4d6db5d7fbc655eb26c3a1d49dc3d7ec08b65b4979eaa76fb;
reg         [ 0:0]                   Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485;
reg         [MAX_SUM_WDTH_LONG-1:0]         I59be2b7a5e95aa90e3d27275839badf750e2f713ff498aaf28bd202039ceb029;
reg         [MAX_SUM_WDTH_LONG-1:0]         I634697ab8c90d12c2b2b2a65d6545a8de51ddf645111a26570ecbdafe71644f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I300f54df5ff39044592d1e17773b678120282a58df676eb35de5794a0fe9e562;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf7a27915130178e3aff7acb7a945422a7955b81a491f1579d88f01797270738;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ida7fdf0874cf846834b903eac34741e8b445fec4ac30ed1451ad758a50d90aaf;
reg         [ 0:0]                   I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6ecf3391cb1fa3dd5e19dee9f9d10088818c528a1feeea04869723baa4e0f2ca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a0182d704153bcdbc1bd5927e4a45326e90a16a9a962183407f29753db6a41f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I044b0c28219d5422e97568291ba0de670fbeb09c83f1eb2943afe0a4be000651;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia82e0334a1b24c5ff4ee87a2d117c3c7301aae9a45e4704b36436f166435ac5c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cf673d7825554846ea143f7954ebee1453bd097d3051107dafefd72ff05ea29;
reg         [ 0:0]                   I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3972965d0045633d150172c2debe5d89bc8aefb8473b1c697d26accceec1b2b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic4b7ca6006b1fc68a4e04414ba1c587cfef6136c1ce1702fd09cfc264ec96920;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib4e8f9db85c1b658d5be48822318c0688eb41b8d011aa69d188be0680d53de8a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic95ac5beb10ecc57a9669b74ccc04b6d5327b39b5a085d6937c1ceebd9cb480e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I32d8bf76f6a512a10f6231445299d254d8fb22c51f6edb2ffb1c69b44804cf47;
reg         [ 0:0]                   I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I100ae29be1331206365e7953c6d6faa026c8c4dd25311560d51afdf2db866849;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iab0de1945cb02c4493fb064c1efb72f4e5a0483452c5c29276c4c7e1deb5087d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib13e8ac762b6740072f1415df276b0ef0703a282b8dd7268638bbdd370a05e90;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7b4e445b2a01b541d52ab461384c1bbb27cbd46e82cd7c401f4350a5e468d237;
reg         [MAX_SUM_WDTH_LONG-1:0]         I70948947c6b4777cf695a6ac2097443bb59059da06704ae1f5c84b42144e4a54;
reg         [ 0:0]                   I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie5e4bdbeb1b832d35e7974194a251885c1bd525aa0c434055cf87fd540b224d5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie12a5b8c714d7783eb66355736714fac95237a0f821071b9b379359f5d6665f4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1b5dfb756878da24a1f7528fe4a866bb750e2dbede6da8548653167c555ea8b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib07212f6fae72454c08283293951d3fff4ff77cf5455f98c5a85218c07a897dd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8af68a180894ba478298d5c06025d929869476ca01e3bee443254dc410fa10e4;
reg         [ 0:0]                   I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9455f55f4c34a937845af7d359cc07d1976a1fb4f3a9e7a262316e137b241b6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifaa7c357c28b482e992040ba6eb62623f7ca590303fe66b20480f8eca1b79974;
reg         [MAX_SUM_WDTH_LONG-1:0]         I48fe5a4d8cc9de9df457625de0ccd81303342c2653cb9051ac93358c46aededb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4a2a60be7efe872271b328a84bd0394ce67c2d59ca77082b5a4ff71b5b5f2707;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51a55a7f067596679dc3e69c0d0fe9c92b776f65ed24981709079891bb7d0edf;
reg         [ 0:0]                   I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4afb194348fb5347cbed837090c3d94bf4a27f44202d58ddde64915fbf8c7bf3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f468cc83b7f0da006d4b41ef40e5bc4e84e7ea6811d5d66b61690d80c82ffb4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I73fa2b0e761bf641629b61aa0508575039d5ce2efefb7dbb1d7b25da2b3553cb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I513c50e5893017204f1fd591753a0f5d29f4b4ffa8466c613a9d12d419ca8281;
reg         [ 0:0]                   I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib2deb611e086f8f21f132eae3b128b0b8dfa06caeab1cf2fe25f94801fc4e184;
reg         [MAX_SUM_WDTH_LONG-1:0]         I427ad9ada9b609bf66d313618975a2a4702011b7ef9e55e40d37db31cf075173;
reg         [MAX_SUM_WDTH_LONG-1:0]         I54c2c2be59b9e302a4527e1fe4136fa3c31561d04ac55f71fdc5bbf8b8488e39;
reg         [MAX_SUM_WDTH_LONG-1:0]         I40cd513b6eb8a99d78aecb88ba332afcdd021ecdb00ee89d894853f642077211;
reg         [ 0:0]                   I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218;
reg         [MAX_SUM_WDTH_LONG-1:0]         I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2de25ddd85167a3af17c87c103f1d19ce367d6e020475b5440aadb42896091ac;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icdeb4cc4b7cfd480c2fbeabb3f8e1ca72b7af731726a0ecde4c097dcf4d8f6a0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib6dc79711e470184d6cc3f360fbefc3c55c32f612d1743111dd6ca9b96c1a4e8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2be6b0805c51599f698f3997780a6f81119106f870a679c00221c9d173040d5b;
reg         [ 0:0]                   Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I09831b2bce6477d49a664abacd23b6be52c85544ebd549b0943f4218cc955bed;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ida6c7b0feb190489db3cdcd850ee5d64baa24ad7fc56b615ac1103f3c5311e06;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56189306e5774d3a224a89042fa23eaf4af107e2fd4fb1f6261943a46f8d8bfa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife7eb04d87c4840ec5a25b0b50ac641fa8ae6ff206065248ad8ac718cbfe5272;
reg         [ 0:0]                   I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ecbe2abd1b3ec06de80c5ba7b5f1ea7bc9484559a134199749c0eaefbc1f3c7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1120c79480e003c87e8160381c89f4a6baddfc6927ae56952a233f96662a8a47;
reg         [MAX_SUM_WDTH_LONG-1:0]         If0294554b2637dc70b079fff36543d68234f3f8e9d80ed67466ad3d8ab4e5f91;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4c82e07db2a69392d528b47296fc3ce9bd342a9ddd3720f059ec38ea10b98efd;
reg         [ 0:0]                   I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I03b3c7c34463d46735abd1392e5bd16a783f79adc25f3471eaede71318ac5799;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8cf7dd68cf30611d1b03b4205f1a8dae3c8f8f943c04773e335a2ea90c555b3c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic8dc799519d1df013b35ee5ba849490330504471458ece8164705be772acf907;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib44073e6dac33e4dc0f497a79d4bdba9dfa398c9e95af1cd3c5406449505fcca;
reg         [ 0:0]                   I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636;
reg         [MAX_SUM_WDTH_LONG-1:0]         I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210;
reg         [MAX_SUM_WDTH_LONG-1:0]         I59b6dcd7306c00a99dad76ca16c9dd989f5dc46e7358a8c0943fae147da7b884;
reg         [MAX_SUM_WDTH_LONG-1:0]         I385d65a11a7e793cb8b1cd9df81bb73d8ce3075e9eeb389c6b9665be6f3c5ce6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1ef957fc8b1559a10bf1f189ca736164c0e50b50786e31c70168fd2e0f65aaca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ce557a4098587fafd3adf55d2195fa2b5c7da844d59ee5c4fd14d11374b58be;
reg         [ 0:0]                   I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48;
reg         [MAX_SUM_WDTH_LONG-1:0]         I384bff3d8617787aa577ea8607bf3f4ce49eb412b603810e854e8ee59ef3114f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibcc6e1c0808d4a22bd66ca467b66a5d5fb1d60d5faef295c6abe67319e782ed5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I26faf05df42ea98f85655adde1199ac6e46b738ff8a2e0b218e2457bac1fc3ea;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id337fd09c4d42ecaedff4e08ddd14fa65c5646caa08bd75d6c274bb9a48033a5;
reg         [ 0:0]                   Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ieb6923956eb85d8a6c65882d8673b841dad39fe763732488f568784d7f5d746d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic1c0ecc66995dc98197e5e73789f8f644f15547d4b130262c526c636458d3712;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee6b04715421c83b0bd430ac4891dcf8a2df5f3fd80478d80de33d83f31d4fa5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6751fa1b7cb41d853b4affcbfbda7f7f959e4a7e4caad11f988e00eec5acbcb2;
reg         [ 0:0]                   I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic3c16686cf48a3d8cd9abf2ee2c917a5dd071e8573454b02340f6e847302b029;
reg         [MAX_SUM_WDTH_LONG-1:0]         I62722b1482f18c3ab03a94e845406bc30c1c47102fadc9b9642096ff3c504cf3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I968319c4ca969a6396cc16b20098933dd8669213ba401ebefcc50670c0fac5e4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibff476e387614c2089d64e400f457e70e4c8ff251bdaeb48e85c68f1756dadaa;
reg         [ 0:0]                   I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474;
reg         [MAX_SUM_WDTH_LONG-1:0]         I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I16a9ad58728f11ad740c8517c5b084638388bf79ef9e4b8e845eccfa31479069;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie73acb967f41ab47a4828279172548c8a36b7b67a4129138f12f9715172047aa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I769e3a9e63f6b86940c9136476d851dd2e123b17d42191d5fa078828c2ebbb6e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id8b5e6165cee66382652189754f7afb582423212885be9cda93c154f46942297;
reg         [ 0:0]                   If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I104e372ee724bc6151a4854bcf5896bd1c49ff41214b0a48b3ab13f1b06d3fe3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia841ffbb8205a284e28cfd445b7b459f11034a0244d777b7136fe0a6009b53bc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia4613fe4f54fd9c2b61f4524bbc42c67307f872c50b5af9e9a836e9cbf8adf22;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic6c4976cc23f404b5b1d328f991e6ff7385f3bb0d61392626bfa621147866147;
reg         [ 0:0]                   I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597;
reg         [MAX_SUM_WDTH_LONG-1:0]         I59b0c136216dcc5613e45a5a841bde1c8243d06cea7caaeaabe614e968228d6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I345aa1fe14f36a465f2bcb4de639be9f617e5d22257cf97f8eb35096383a8674;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1bea08777eb6009228b55fb534f502ea7deedeb705d33d4e56a7b5107a9a11e2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5d6f4230452aaeb0bd33f7b39b467450b11175685cde0958391f4e7f5ce44847;
reg         [ 0:0]                   I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I328d56833be24a38552b6110e2858dbbc3561a3783d9255efb5580d9f4071749;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id835c902546b418343c3e52de8260db4304844475cbc1532389305577624e4cb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8e604b3839cbca0e894ecdbb66a3c24f49a91c523f29e8984fff3e8bd1bb421c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I402b028195ed3aa64305d0cbc85fa79e1f172c79704f8fbd86b74770352a2908;
reg         [ 0:0]                   I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56ee0a1de27160410a2bc12cd4d550a3fcd4d560d81348cc36e94746f46f6341;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c0d3684d621cac560ca9866f49e30d1f66c34c35b2e1112f078ddd15b79d826;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6f62f4f2fc06f1cb30147da56b8fc88874f748262e4308b0d794c057267d9ac1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2054d562a308ba04e604931976e93c9c55bbbc95d01e5504ab55ca3d8394f40f;
reg         [ 0:0]                   I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3d365702f31c0b491b205449d36828e3fc8ca71d1e5b3ff872f9eda67fb06e39;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9cb1f43022cfd63f00fe801b2d938c16277eefc9dde55af7c332011f60180cb3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1deac6b91e43b89f481b4b593e33836db7cc46ab37edca0ff7eef8ad6b92789a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6896936df9cb439a07c80302e95b21023dc476bd78f678e93c7ecf5e3a159216;
reg         [ 0:0]                   Icf75206b75ca695f888c3d924d2f1822806f452b5d29a0d6084dbd1c00a15790;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8d320b2d799e480d78887d5a1483ff7fe5f1a986d75e808863a9085bfc3634fd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I363b3334e1423f125eae3636a561c36eaa744a2c8c62718fbc648dac5ac407d7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I05044427a4868a31ef17917e7795eeb32270ef20859f5d3d4699fdd408c210a2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iccd6dc287621f59bfd5a38c0a5f5a06e1195d0d5f465e7129b782ab12f8e01d2;
reg         [ 0:0]                   I4a1896458491f2613d2c7274b81fbb7a9d405272b871b504455b388a3695acae;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2de3b409715599c65489338e9218150f6c33cd987ece5fdd9c7b2ba5c06d3d60;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie388d32b93fe9ae25426208c96be3b8dc61e43e909c7d28facb3fae96dc366bb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I076abe19140e558596312bb8ed87bfb0490feda6f1ef7c0ac1df979cbfec7c06;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a738dfeb0fa39730802cd687a42613f8ca1967c0042bd54b092c2e36abd47f5;
reg         [ 0:0]                   If122210c8dc39e7ab2fecb27dac5c167b39ccd9e8e4cd076b2b3b92632357248;
reg         [MAX_SUM_WDTH_LONG-1:0]         I56c293e90676ea7b55934e3064087e3a4ea95a1c6ee3bd4d606afabce05357af;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3ab7d65dd9be4dc787c343b0e877e40ad8b5ce9299098e4f9cb86ed25fe1d1f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I20dcaab9d6a12d0b868ac37762ddbbf0199ab0aab46594b5775a27656ff61d80;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ice4daffb593d295aaae1b2165bc2dc9612bf70ee6005a4200f764c76c430dc32;
reg         [ 0:0]                   Iea6e52ee89805cbf2f2a65f695323d8dd7669c23df341897eff049fbcbd1db98;
reg         [MAX_SUM_WDTH_LONG-1:0]         If32e43e89968b9f008cb77759dc7047519d200c512cb11c105b74c404603fc79;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6740d7cf9a56e745fd86c9131b62b2dba6a7ae614338a59607a43f0b77d9bda0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I10ad038fb26d337df3013912d38403548cb5e12d6e175518ac7e924e583e1fab;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie103edeedef5ea626306fe0162187acb812025558381c8ff0ca8bb006a2caa17;
reg         [ 0:0]                   I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa;
reg         [MAX_SUM_WDTH_LONG-1:0]         I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I082f12331831c80bb11a3660e45ab9fa6c122af71c82374eb645f01f89b03a15;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie65f8e169c71198268320e9dea6a360718a61dfa0e33983344ab5070a97fe3c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia1df41c6fad9069c1aab753a907bce8625c2d114c156b2e2c0429d7df6c30f17;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2eb3b47e1f13607457b31a324a263038853d4c7bb85f4c9c00c26c16403dfa7f;
reg         [ 0:0]                   If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia556763bb9b39f7ecdea64ef734cbbbc108070aabd560d87872fb475201ee4b3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic0d0d1aa735e38d8af824759f30badc83db776ac7871d2f5d0c12594b25342f6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I33ceeaee9a8251525af0cb5b6c1b9968c58696493f1a3ac45cc5c0e3b44fd5a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7453e7476c16ded7f06fcc1f9c11a504545e00d1e15faf2f2d0cfb57b9f35c5c;
reg         [ 0:0]                   Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236;
reg         [MAX_SUM_WDTH_LONG-1:0]         I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibdd02bba3f13be2c6f23b969be65c45c5a1b1d42b06a5189c10b452af7b1e055;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic438ad9f1da18eb848fb486bdc7fef62f7a3ce12e948699f5aade5c2922e572c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7abea0145d10af48608127e2828ea265ca8883f1c43474ec82b2e24da693c566;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9aafd88945bf07d0d9b361fecf903a4c1b14db6dede3d95677ae0d01d0e36894;
reg         [ 0:0]                   I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7bfebc508c949b2dec0ac81a1029eac23947dd8b78872b238f1ff1bd0e19676;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibcfce28ff0415dd2da98a7ec1b48f013c33edb8b6224ee7637478da2889b6b16;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie2c653cb0d05e3e9f884f7e78efe071774cebd49008f86c8106fb180e8196fff;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia709de664b32e0acc613ab7448eac9837c7cb75de3469262a56bf32086894ab6;
reg         [ 0:0]                   I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3feefae60ec0eb2602217fb4db5cb7bb3d4af0e5d6656f09c286220f83c14e95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I588d1fefd4585f5eccaea213e11f8d74f1308c3bb15bd7e88dd5275ef62e236b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I211af75e159531ef945adcb8f51b79d5b1f27ee3835f2cc2f79124b235c10a72;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibd0e4e5d04591535c937a5389e0763279d4c267e0d0d7f1256a9271d49892307;
reg         [ 0:0]                   Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1857bbf85d1336737426b53588e78aa34ec0664ec1f3c4bc351040782a0c1719;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib5b72b3ca0b1aa00d12330c72c5435ad4ca90d598d05e7790f1da65af2f8c3c8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24f30205c1eac80e3a167d5b52d1328285db573a6671ad7e635e47f49646d05c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I26ce0fefb116238e66b72d526766ce8f9b9d1de0df15d835668d928384e44827;
reg         [ 0:0]                   Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibada8912d6b4053809b28c28b01acb109cd1c80309a62b9b5b8ae3b5a0ecc44d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I698dbb248637786ce7fde5591c80178aa213872056e5fbcb46cf7a23484143ed;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0d5b3b10a05b9ad2d2df1d67a669cf252f9dad522d241643ad3ed51b610a32eb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa2c9985b7daec8d06c292ca451d71e14a32aece2e26dd6d5ce3f102d70ed54f;
reg         [ 0:0]                   Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6f84b4bab9b97d15495d515da0fa036b9ebc5a7193c2544274b3121dc23b8ae3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I922ca03f57cae28107251c50af6bc0b96a46be661f758e93f2b80d0c23bcb02b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I60dfd53c9dda263ede70e2debced85d2e29fb7f897347d5fb6bbe068b5d42b6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4b915b467967001eb1ea2c496d782c2fa9506073cc4441ca6cc42f67e57ae822;
reg         [ 0:0]                   Idc77bba153be5873f87a4cf88c6ddc6a89bf8aa3ffcd29702126b01053f012f2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1ee241dd9ec346bf09b25ccd2f1669be719a1411914d367372a46c8d60cb0f44;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia556ece4fd10276fd9d7e0b3bd79ab15221b0891dfdcaa8a3d3f0988a356b78c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9dae8c584ed5197edc44374d711497fb81a91de44e3cc12d23de36f3269fdb65;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaab44235fea66a54e56d75bf5d2732a95042c033defaa2a906b2390bdafec03e;
reg         [ 0:0]                   I8674756fbdb78fab124727c8154adc4dcfd4674e3a4d9977d2fff619cbc42e5a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia34cf7cdac966a47b902c17ef799ca34f3c17e4f5a410b97d7f07933b977db3d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a2d4121a3aa27634d62a6eab291465d8c2ac688a263dfa0d3fa9e007d825aca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4643ca0b8bb8f9d58565dac92705b1e6ef755a8edd307a0105482001c06eea13;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib13dadfd1a4c8b6664863bff922da75c848e4e114e53ca32d4b93537cffe3fc6;
reg         [ 0:0]                   I4a3c7a36a82811aff327ec55776f5077aec859d5557df45568abcbcbb0fc5d5a;
reg         [MAX_SUM_WDTH_LONG-1:0]         If017b6342521fac4000803837465d5793375e9f4b8c2d9fda18843ec7b9e0752;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iba4a2105d76cbbbbba7cd474dff95136225ada8b4e62e607962200b0caddacef;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0a34efae03321f53acc6f183e7c3f22df19d0a0add67ceb5edcc38046ec33748;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3189d8c7911fc25a6079d7e30557a3b7721d0ac84c03b38366c1db55c1d3f95;
reg         [ 0:0]                   I931f943f5db8edf3580ebe67b3da2a0cc9a1b68ac6485930d6d9dc792bd36eb3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8bc9b50c83facba8db598d0c5c71cf811e181fd16038a08f5aa04f00ff2bed87;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98c91ea87b40d44f2e5830fa4e4b285baa5cfadd6d5419e88936592f664d8340;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic458bce5868967b65093883a779b50f1d51fd9fb924eb6bdb9933db186240445;
reg         [MAX_SUM_WDTH_LONG-1:0]         I20382630b2daac9cb982d267670777192b41ca7e729303eb524e38603f056031;
reg         [ 0:0]                   I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8663595964ca4eb094c6cb80c0eb4ad319673883a254ccc35cc4be73ea5bb00a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8192c0915a9b5e00cb68ec0dd1c26b26640f3f9c6e17e3de938b91fba44e3782;
reg         [MAX_SUM_WDTH_LONG-1:0]         I886c2494bdc82c917ee66135ce52c761c347c8fe42ccd63d769cf315b338f2da;
reg         [MAX_SUM_WDTH_LONG-1:0]         I24f0d7d25ccdb1594c03394c4cfccf9327de3684e2376c8f06e56077931820de;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibedce4b737f7d1af34a1abb100d92a4a680c939dfc6cc74ea55aaf139e0b9bf0;
reg         [ 0:0]                   Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6;
reg         [MAX_SUM_WDTH_LONG-1:0]         If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29;
reg         [MAX_SUM_WDTH_LONG-1:0]         I217ef743b51672b0333da788f3206b6ca50dd43195a27a9d1aa1b542b7f3c77b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8863222d9076063d0d2c673dfc8fa35d8fdb87a6b37ef7f98988e5c780d556e1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1a45983bc2d6c4bb8453ee08cc254497e08c85ca326de079180eda79e4a64b55;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6e02998651462a264077c956dce9fffe5b787e53970bb3c192ab8ca4041e7ad9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I72195f5a2c9e92ab9f5534742a45619c0c1840ca7e3955e24b7af70807d5a4b6;
reg         [ 0:0]                   Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70;
reg         [MAX_SUM_WDTH_LONG-1:0]         If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1cf05db080e64680bb79c5be7fb32bf5c038ff3ab7396d893b90914ad5472bf9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5249daa78d99d33112b5384478d38b33a088d48e042e4b0820c40fd027c0223f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f768fb70d35694f0691521b3989c85e7ce64041868b4f611ce7020ca3bbc1d4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0dcfa4dc673b57614cd3760b4c618e128809db705602e53f5bdc6f6030b54a50;
reg         [MAX_SUM_WDTH_LONG-1:0]         I64ae510b10cfc41dc62dc76faa1932a4f159c6e2f4b1aa5e618bec62a190315d;
reg         [ 0:0]                   Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48;
reg         [MAX_SUM_WDTH_LONG-1:0]         If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9cd6f2580a6f194817cbe4874192fab4f22fc58228a6deaafad44e14f2c27311;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie5f920e3e83787bd026f94181b522cf7f247cc0863da71e59f8291dcc4c43de6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8eed9a916e362776814cdab4ead58e68fca91b54a6648993b57e919c07e132f7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I859eda2ded7b867c15e420278c996c195f0217d795b6d53acbfc10d218279f02;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa68deabe5c470e4f9f865f60e32710252f5f104571ba859388fd37ff0ef320c;
reg         [ 0:0]                   I7b3ff601c78f414f5f48cde79235444d13872a0527c054356b3af150315b0949;
reg         [MAX_SUM_WDTH_LONG-1:0]         If15a6d2660b407d89dda6c113578519092d37491671c47feae8a7a68565a9184;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1848915027beaf897f1fede8fb30fe33c1f7e5a565022bcae733a9462c9c8447;
reg         [MAX_SUM_WDTH_LONG-1:0]         I318c86cd2c86410c5bb1decc6f5df2d544973c518750df70527d2c1fc0b2947a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id69048c2098191e826ad522a678bc79cf72544621a8d1d2ce28f0c5797251fbb;
reg         [ 0:0]                   I434491ac49be9939ffdcf469991bc3d23ef217b8414c677d78ec9a062e74ba07;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc0fdfece0d7aab4a85b2874a047e1bd390aa826df0d979166e8721339410c39;
reg         [MAX_SUM_WDTH_LONG-1:0]         I54fb2b89dce635f5e04010aa85747b0fc135cbc6f58f5b1a92414b2b82fa9e3b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifdde108a572ae924a2890624cb24fd7f4beb70c6c8942886fceac443de8633ae;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0af9db61e66fad28ef275cd396214b69dd646a4b79c44e1673c4ad61458d98b3;
reg         [ 0:0]                   Icd717b9b3dc725b8579e62b042051399a3b21cc10076de8e0bae480fcd24d607;
reg         [MAX_SUM_WDTH_LONG-1:0]         I09301323ed69c3f202b9693f2db743880d6e7618dd91405aaef90c34e61d1caf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib6c59e6ecf314597ab396dbceb18037c0d32f40a9022055628288855ec99fe95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1eea8e0dc933632ff46ad76cc672689ea6fb253ee0c6168d915353d14fef838b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6bd5ddd44f3524fc7691c1957820f067009d145a484faf5edd0d2e527836e12a;
reg         [ 0:0]                   I0c556fb5fa4a1297825cab8dc64089faa86f1cbe67bf106748d927849e16e007;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icb4397b9bafcf2461e592a0050cf42f2832d3497c940f82fbe98e855a1153129;
reg         [MAX_SUM_WDTH_LONG-1:0]         I193b91d093965a3b2d7ce6cf215348724929cc0c1a3851f9885f822cbcf9ccc6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib31c2929d1523de377924c1f54c6a251313afcbd3c1958aa3e9c0e097c391485;
reg         [MAX_SUM_WDTH_LONG-1:0]         I60d9fc72ce19f1ab5a6385844f0660250ee06d76e80845945bb345754280418a;
reg         [ 0:0]                   I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia5a27c8c5d46b95fc3ca75cf9e499c6cf406d7320e97b8e0daffe069322e6466;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9bb7b61602527be7313761f2a4d22ca145be6a35d06702f60aa9c6c05e9e951e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic3229f0918087445c3b245f3b6a66fcf9d241cf8c9b7a22ff7cc3f127bea4dad;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac6d1591feda87bfe1caec1ba6e2a272327d77aff99c6f47f8907caad520100f;
reg         [ 0:0]                   I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I389c3b8f8caab2e397e5f1368db3c31b6c9d81578e1c6ff3c77614bb3fa283af;
reg         [MAX_SUM_WDTH_LONG-1:0]         I261d8c9755317b6e7d448fed52871b8996ee8b2966c2cd1c0d9c8c4fff09c1ed;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8802f7a26c9a45d00b3c92f9d62988533adc832b43fc024798ead3130d41af9c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2955c07f64b9d8ca9a7a1ea0ff4fcc472588cf5046e22d529a9a674e264bec1f;
reg         [ 0:0]                   I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8e2591213eddf0e31054520ebf62ecfa31656b0b4d8cc948e2f0ad6705f72967;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ee55f4d76c10bda1e1ff4074e72e0c0e51486a3659df6c99998dd58f48ac2cf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaf6b2159a554a3e4e02eed8fac29e769a0ed0b4023fc888e72167c90055b82bc;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia11f0a7c148064962721b3b128e05210fab5edf48970dd483ba21c75d7076ae0;
reg         [ 0:0]                   Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibcd8c95e386f314abf1373ef45a9e95ce079f6eeaea2beeed3118823f184bfe7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8cde7e5629b3ca36c06d61c7836e7944e7fe1f12ee5bb6722ba97f125eaa5d54;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9f8966a82409d3b30ee1cd52c7e0b4976cd317c1ec6bfd7c6c23e4157a556d9f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id1cb12cdb0a13b705c9450d25160d92c2ce8624a1fdd447cc4db14c29512be59;
reg         [ 0:0]                   Id3bfe7fc5e0a1ea258f912127a3c77f7cc5ad791dc6166266f64c574b8ed0e81;
reg         [MAX_SUM_WDTH_LONG-1:0]         If999edef9d50e83e5c53e4715e8f0ae2699c9ad1960e7e16ec5049a8ce0068e8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I281aff7f22feb2745825babc1e61ce1ee1bcafbbe54bb01b19ff94ac6ad162c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0834faba181b93b43416922703257ebf7f2d35bcd63746ca52c83e57dd801731;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia61ae97a6d0793a9e542fbebdea72393e93d4e1cd4bd260432bec83e5503116c;
reg         [ 0:0]                   I370bb7df3320249e804ee9d3d371b1e82809433e4f7e00f74ea0ab59252f4176;
reg         [MAX_SUM_WDTH_LONG-1:0]         I17d1cca0614280eb976be22c9779a9238712e3fd3d27b84bc092911227433180;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icede982a125cdcc6a88aab18ffc06e98ca57e02601729b20fdafef5236a03ca4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I365aeac8393552a9c42403a734816538b26d9c1429d9dcee2ac6d312fbcd917b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic7aa7756d5779803ef1deba260ec7a2dfbd59071f84e0e73118751dbd57b2737;
reg         [ 0:0]                   I3d17552542ca2452e4f458fbd0aacb1a5b62ebee4be942ac561b87376658c9d8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I20665258f942651538aba58d63ca7f531a375ce0ad65c83a1aad4cda0815b334;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia771e5a1a22d051469c95101abb12e406a5aa0518905b1c475fd4fa0b7fa520a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9af1d3493b4b64704551be835abaf50ac8b247571a802846076fcca1f5f8fc6b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc0a08bd18253bf9fad9b320fb7462c70107db49b1c8f67126a9bcf2734f54c2;
reg         [ 0:0]                   I5ae887c145ca6af35eef2229e55c297f4b6ffe0a2cc47e55e6dbf09e1f11a9e7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5337e70d66d8fb81df05813fd3a172c8337b5d2ca39976efd9dcaeda77844be7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I75bb712b6207e8af8c090db486b02880a7c3f82ca47a48929c52e898e36967fc;
reg         [MAX_SUM_WDTH_LONG-1:0]         I05e3db1dd36c0de58cd3d6d5c692cadb9ac76c905af96474615ac491db900051;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7a6454c2bea6d09f07fe94c2c000ebf70ae11e4552e7e6e2e1d53e09bc529e5e;
reg         [ 0:0]                   I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238;
reg         [MAX_SUM_WDTH_LONG-1:0]         I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc7f54032db8aeb207641aefc8926732096c74282c740ed04545ea01d1375d62;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaa2a9a1fce1a32dd04ceb055eabc32fe90fc765c2246d2a29f0e847a8ab49f1d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3bb50ccd25f72ca813c999533e808c0dfbe3747a6dbe023a303d64e0cd571423;
reg         [MAX_SUM_WDTH_LONG-1:0]         I32f852a9a6c5c496bfbecddda78b07f0cff10e6f360c3938827fbe389bbb1d64;
reg         [MAX_SUM_WDTH_LONG-1:0]         I79162ac11cabd67e684b36c8633d4a001a7f794c60468829974f8ad972e9b6d2;
reg         [ 0:0]                   I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I44868fdadaf261c99a76756dbc2feb061aa5795b84be4aaaaf2b2f14580d85cb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0e0b35e726d873d7a4d436a763ba90d981031d080d8030d7d1e11907bb246f06;
reg         [MAX_SUM_WDTH_LONG-1:0]         I35bb67b450432187151294ded11a662620636aed3ca3ce1396869fa2b60ed816;
reg         [MAX_SUM_WDTH_LONG-1:0]         I90bb979f2ef58854b3b2a7d6b0a574774403e9766c60b1888f1ac97ccf4b9889;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ieace5fcde163f3e9bc1be0f05b04d00432343111a05c7195e0999a3cbb3d95d9;
reg         [ 0:0]                   I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8dffb8fb698239dca36a5371fe756164e127a33e709084a74d3d2f548edbe1b0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d8b7acb9dfc4a40ecb4156435977770c6a8f6713d612777664eb4c545208943;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icac43b0373871bc847869a8c5a86a423b2bf8378da0d3f1753a42ac604f5785c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I309283aa468ebadbc72fb7bdb48e76697f5222c1e527837ada3ba12084ceda60;
reg         [MAX_SUM_WDTH_LONG-1:0]         I055caf108b4457e691ec20569b48a56478f8b0cbb9211271c3a7cb2836605749;
reg         [ 0:0]                   Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0bf924bbc09ce9d0e83a26d569bca939f3bd410a63fa3b1ad631798a9171102;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3896b59b701e291956a090ff59ca6867a6267fb825629de82c88309ade2dc8a8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1112f35be1ed8725b875aec8350b0843ebff9231fd3d3a49914003c23192822b;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic953289eb284e6e85659eff600c7b373dfd72773441baab0ae1ac4585370d79d;
reg         [MAX_SUM_WDTH_LONG-1:0]         If07db5ea1a4431d5d3e3040559bf352e46983992fe80c37e84468e7f798caacf;
reg         [ 0:0]                   I00fca56df853315156adf3a6a5cdecaf6256b108f16f65b1e93272f0c7796e9c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7214b0ea3f1135ee6e703c8e873696254a514ff1e88c32d42757c8ed40a5b907;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id66a032ba386ed0856ac30d1393b9bcbdd32f34a514b18903c95fc66b287c7e0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I41dadde0137c88dc8b0e9d86734803a46461074a08c6f61e73c8cce898ce64c3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I55543ecec7c46f5fae535eca894545a441edeebb10f1b2bfef7c7fae234cedd9;
reg         [ 0:0]                   Ia6934e7e07061fec0575e9ceb1910150463d7c530d30091ee48fcc50bc2d0cf8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib9f05dc23ded7e25eec5344da5ea617060c2cb525c22aff7dfc41f86026b864c;
reg         [MAX_SUM_WDTH_LONG-1:0]         If7778495e794f7ec0ace1408db22f95ed302e9f124858dd6e119eb3c91520821;
reg         [MAX_SUM_WDTH_LONG-1:0]         I047343beda3ba4373e81c19c51ea3ccd5320a6ba2a595860f87ea9e041afbece;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9138132d9e54b759171955a69beb971d2b73d6cef41137e9219277fd7627d6da;
reg         [ 0:0]                   Ic8358c4f85a5a177702d111cdd3e705172bedf92a6d01f2c5d25b5e33c75538d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4d36f91f636848b5418807d5da024cbeb73a4b63a9b55c2b9bf48f22f2196857;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5a11b582e017795d316b18512d5f7809300e13a89ee878deccdc3e4ee9556e3d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0f690c5588c55c55f7e38c94b4b0678f65ea3214eb2b3923e6888f15ad2e632a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I36e15452cc41552f83da26036b7b94a2ad425d1441a3de1d4e226851a8bcb3fa;
reg         [ 0:0]                   I2e37b13b583174f0ca14a3fff3bbdd50d584c2a917a020de586b559bb7df4c45;
reg         [MAX_SUM_WDTH_LONG-1:0]         I55699a1c81182c259ac531c5587702742eb60c998c424e33a62849441a5a94fe;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac99102c92e103b1b841f87f7c024aead79f11f036aff50058281258beecf469;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib74288457c278f35939cc8e326fa0db500d368d628b4e60af7921c79991a45d5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icca50300b717929fbd20809910f35bd0b6fdeb04585be02a41a9aeb2b23e0041;
reg         [ 0:0]                   If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0f6953fe9ab3a2018fcdf430ea420ccae2fd35b2acd637cb083370cc86155cc8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0ed51fa81db29c53a4033d2a60ceccacaba9e1abdc340f1226e4951b8af1d49a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I15f92f05ad628c0f786341269ec6b7aa37408eecb1415a026b776fe4b1ea167d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id182102124b3765c410c79e6b7560532537d8ce5d243f64cab3c4a73ac894292;
reg         [ 0:0]                   Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601;
reg         [MAX_SUM_WDTH_LONG-1:0]         I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I92c3d579813e542874bc16d04e9aa52c9f79b1b55fab5f166c74f6ab61bb195d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I552bcbb774b1f6cbc437d0e597e9f85a058a1c86dc9327c0ac420c6cd272adfa;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc1b7731fd55becb0c39c2ad581762a4053fa931b7944cfbf14ee41929363b6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib2ff21fa69dd26a3b35833b51981a6b4e03be26d774d933dd860357d347282e0;
reg         [ 0:0]                   Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icf03aca159cc538c2d6f4b1b616e5c6c8dc4f66dfc24b50408e54d746671a222;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id934d373281e6054a71d367d79cddd1549b8048fc9fe481b15c8b8f6099e9468;
reg         [MAX_SUM_WDTH_LONG-1:0]         I381168c5956c61f426a711cb5861a659681cc9f9772accf6ecffd355ce8db307;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic7195dd57a1287cdadc40d619ee55d7a59d4a02e624c74267ab5a631dc66a6c9;
reg         [ 0:0]                   I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b;
reg         [MAX_SUM_WDTH_LONG-1:0]         If27abe3474af746eb5d14fbe518daf8012c4ae8f65e9972aced680995387a413;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc36ad96928d2d8544d21273b9764c7dc17dcf79447e8ad92b689f9c33debb62;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia3a1160cab48ed755a51597f93348a5ff2a29df29582523f0f1051175dcfd3a1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4b4f2557be01daf1e3a86e3900f7220915b80fb490425d6bfd0e6f2ac3d758d9;
reg         [ 0:0]                   Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I59d501073967763b8f11f100cc0aa90180a85e7396d40479244bd2a74e1bbb81;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51dd1d6d9f1dcdab1e85e392e5fffbbb22555f9bc89aaafd686ee55bd8dcd14d;
reg         [MAX_SUM_WDTH_LONG-1:0]         If117910f998c5992518fd3258d34731a1dd45db76e7af467934d5c0b8b455c0c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6414021c1267477ff6a5b8899ac081a7f3c840f899c3a08b1b42ca91d37f945d;
reg         [ 0:0]                   Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952;
reg         [MAX_SUM_WDTH_LONG-1:0]         I5375e515cadcd87ad137d29768eabc89cb773c65f1838f17762632fe6915b805;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1366c2561d741ee41e937b32668f5b2dae17f38f7ab9192ed8d4670e570096bf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4ed1e2ce8c1861ad771d926c40a92a3335c27ed9c927da2c4b4c8d246f888cd8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I34dbafcdf27f8460fdfd7a329a955300c42889d6f99e9396df4fcf0a80d7e84a;
reg         [ 0:0]                   I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9fbba72f6f8a1120c18220196387259e4e2ef9be67b89f4c4d941bd2716c16b1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iaf9bb39df39518f42c265087053d0e659319b41a5ce82aad117fb21646fc5811;
reg         [MAX_SUM_WDTH_LONG-1:0]         I23a214695af25c30f017977039b6522a79e1ede0b71df88555b1a36a613ea32a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7d3dd2b2f1be7541867d824bf4cdda33f1e8e6acb187e6f78ee354a9030dcde4;
reg         [ 0:0]                   Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab;
reg         [MAX_SUM_WDTH_LONG-1:0]         I242b12e2ea6f2cabed454cdd179b9a0b2ea51a43ac2c450f84ed2c650a2cf789;
reg         [MAX_SUM_WDTH_LONG-1:0]         I66e51d57d162e80e54fc2e9bfa91dd74805a0cd6604ef63a5645f50242e2397d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I610a848a26543d03e396503018f1541e8a2647f8c97ebefcddab43e6cd91ad88;
reg         [MAX_SUM_WDTH_LONG-1:0]         I16852d5801d3a353a9d084a0b9dd4fcc537eeb8277037f64f84d1fd1b1b42102;
reg         [ 0:0]                   I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iefb3d17f1de1e179afcfcf9f8d209375b9cffd7efc7f3ae88ca55d6c58b0d7d6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1abfb953ea909659ae25d197a2ecbefc307fa6580318bf8dfd723883f2cb242d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I388e7ed193084e1a629828ccb5e027b54dff58603c1e644f81fa233d8c397511;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icd26d5b89d292b0466a08a131e8d00b1da2a54043a429e61b02f38a292c980fd;
reg         [ 0:0]                   If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1932bcf87fcb5256afa2f82da25621ca1cc06f6e256ab9b05d1b3589613bbe02;
reg         [MAX_SUM_WDTH_LONG-1:0]         I807bb4f93cb4990ea3d0b5f5bb5ee1c9e281eadf997a92a32fac10d917439ac6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ce261f7e73a1bc919627efb495dbeb739b6b9ef526e0d575ab46524d6f50092;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic7138f5e1ef57f1e0d904946b13c6e16a293b6fba7db6266a9c40079e40c8e2c;
reg         [ 0:0]                   Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7baf74b530afc8aa64e5a9f2b7879a0a6573eca1818262c1ac817c5940b0fd75;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ide134ae79fa666de582a416826cc2d4a579d888b98b3b820f3c5e445767d002f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I76566fde1f58392124d201e9b66f3a221ea658b9be074b36c54773b34997faa9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie8db353155b2c11a919ec581a22860b11997a2ec74cc8be6c36b04716c9fa558;
reg         [ 0:0]                   I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I54f9f4218a4fc5202873aa8c9e0fe7564af5e7c244d438f8c662117204056632;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e64afd49b1b6224dd6a8f10660ef803524895019ee93a630209c21f66fdfb26;
reg         [MAX_SUM_WDTH_LONG-1:0]         I813a94c07943df9b170773639811bb908b1dafdb2a89be0d53e81e2b98faecfb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3a3f389915c4e6367d45081282db8a902b0acbee573fbb0da4c5d935043bc2ff;
reg         [ 0:0]                   Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8a0fa39f59af823fa6b73d097b287483857fcaeb20ec459e4fb5812c8774a796;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id0ab6ebd5d082a3d961cb6b58b59350db5bd2c3d85c08a14901f6573b80fa446;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iccaddd2cbff52541bba9854cb236957b9ff6e50e07f2be5f60b08fb247e44962;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a6d992471765834fab17a42d3d419bedec8e1fa9eeb10617930e06d2aa2e5b8;
reg         [ 0:0]                   Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02;
reg         [MAX_SUM_WDTH_LONG-1:0]         If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib78e3653ad432d8c12b68d0085fb8deeb5405ec0571e9153bf204f598fa23baf;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idb9e9500623a940d82d7b77b7c613132875cd4287eec27e495a5d2a1fdb16f6d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icc42075b4ed713ad08010e19baf3a6ca84a9dd07cdfa71d60c1b6d05634320db;
reg         [MAX_SUM_WDTH_LONG-1:0]         I611cde8f0d43b4ca69572460c144fab6ea9088b62f7ee7ca6b2618893e002359;
reg         [ 0:0]                   Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I41e79867cf93976d9e1db38f48b70e6fc09fe4ec448856483d064ed9ed2f5055;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iad7a7d92a71ec5a2a4ecfae6f78716866da577038b41a649d32a5c4db56257ca;
reg         [MAX_SUM_WDTH_LONG-1:0]         I73866569df6c4e95ef7273a1370e9da252db2d74b0df1884bbf87a80a05a8fc7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I90c36434a94834ebe700c144c2feb5f0b2a543bc43692f5a23b5b5495d417c64;
reg         [ 0:0]                   Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436;
reg         [MAX_SUM_WDTH_LONG-1:0]         If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd;
reg         [MAX_SUM_WDTH_LONG-1:0]         If3ae39f173044773979d138817d4e808bd30278aafc2968e47e95c79c1bdd88e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I417c9ec039c09269659f1426df4443750e00755cf0694b0fe5e508c563e114a5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3351df654db39d7ca929147d06b79348195c4dcac3d4f398ef2d7d4491a151bd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I76e78b4f2c67b24b90b5ec2d4ad5f189296fdd4f21eb6eb8600fdfc9dead405d;
reg         [ 0:0]                   I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2;
reg         [MAX_SUM_WDTH_LONG-1:0]         I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9a7c4404df96e54123d0a04369056ed0844a3683e09535b029ff8896fd7bd60e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iddb4bf2e6f1f1c5a0c910c4939447f53a9794ded6793cf9fd33eb927ff22833b;
reg         [MAX_SUM_WDTH_LONG-1:0]         If0c7c112ee1274d779fe816a1d31c0f6c98d88491fb96633839a9ee0277d1a88;
reg         [MAX_SUM_WDTH_LONG-1:0]         I107b0aecdac212418e4f0054f31ea2a9e89dd7d4620ec8fff0725e7d29414853;
reg         [ 0:0]                   I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id2edbcc00e89016e0bd07ccb9dfab560cc91bf111ce3b460700435370e90e2fd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I35e88d9a4df07df57aa080c63822b5e79435d28c2f9655a449bd68dcc6aa7709;
reg         [MAX_SUM_WDTH_LONG-1:0]         I93523e2e245808a8657c66a68778e78a2b7d90f2d076f0be05a4ce53d5803d17;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0e18a6aa6a4f5814b2c895163df2b575a04229c654840b386f7654e0765ca631;
reg         [ 0:0]                   Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0911515aa6dcfc8293b4c33ec6d3d7a6227c26e3de3ad8fb3aceca8473c37bc1;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iebc32b1def039cd8820e6149458d4008738f72a7ab9f73448bd352b362c0c852;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iec3e7529badea1bdcf7d907613c7e25860e379167f064645f36c73bd50d9bb7a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iff7936d861e3a88db1b8e9c2041b7f61a956e483c47f8f16d721acdb81f69c3e;
reg         [ 0:0]                   I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idcb6f68f9742159aa2fe6947a2f9784ccd2b9d36bd3864ac8b6b38c842f5c5f4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I925b92518cdbfa9b8934753a60adb3c96413a57c111ab4beade1b677548443a9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7352b278443169fe5c6f9133c12c026cbc017f6a07531cd9c93b8d58344123c;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia8379750d4b5cb8da49adad32a77ec592f600fa74c5e099458eeeeb93ad133f0;
reg         [ 0:0]                   I99fb6dd2fc4414a231a70d23f26ed6b852ea4a563b41d3d8aa364e16d953eeb3;
reg         [MAX_SUM_WDTH_LONG-1:0]         Id6e462224a7c7f18670d48e3a7c6d35465875f9638395e7dd87b3c494985d418;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d2b275c4f7f134ee6a3999c3f0223d6b626df4441f891a9427d3d8f1f725fb7;
reg         [MAX_SUM_WDTH_LONG-1:0]         I60ea282a4be819088dc3a40aad4a3031c831802d89e57d4c365a1a4d4ac86c3f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ieadb5d27e6ce4c37e58646b5eacd57fb1a249461f9d16576dcc8bdf46bf4f3d8;
reg         [ 0:0]                   If0e6db2779536df3835ac1e3c316bb7d9cf2e88aa7cb70f5b05563886cb4f3bb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c0782e7324e49c90f18114dc327f50948f9bf80b906f202a50b101832a88baf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I1eedc611ca90fc435e769af408fd45a0299a28c0ad26468af7e870bb5fa26608;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4872d474646c996a00b01718661c079771beab1291ba697119f4a0163b5b061d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I521983a9bbafb4754207a50436a99446235ae7c9cf0070958e99082cc336cc38;
reg         [ 0:0]                   I32eb2fcd88eff04a6295199db748b576fc1d585c2ae058acbf3150711574dd5d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3d8ccc88024eed4b5d118a6c3b8c06553fcfc8645a8569278e7e7e8d3b41597a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib0e28df62d3f3d60795ace1cb4975098004b434da3773f09b2f829c6ef7a8b21;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2a58a1a6247cd23a2e2d4ec408d68ca9f77d6331a8a67f975dfe0a1db72f2bcd;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d712b4bb4e09ff4a0ff934bbaca37083bfe3fdd143d20c9f85ec220700af40b;
reg         [ 0:0]                   I244e0f2c03df982bd121a8a0240f862b4e0212ab54dbec0984f987577faebeb2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ice2f6ae40746fa0bd1c5b2db1aa0bac608899f3ec311d6e8459e126e446f7947;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia36b5d24ca414ff96899820bbe3f5fc319b1e82dc558c2ec8af7559b6c45992e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ideabf29ace18ebaa3db078d782fa2d3b2db1422ddc35c86dbb12c94f172ac364;
reg         [MAX_SUM_WDTH_LONG-1:0]         I82214920f75f46eb33a8b5e21ea60398b1c58a185ecc19b1ada4e7cb441e8773;
reg         [ 0:0]                   If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec;
reg         [MAX_SUM_WDTH_LONG-1:0]         I193ddc6f5bac9d6f9e6599d78ec2c22aabe3032583f3dff87a62b3dca9074fa1;
reg         [MAX_SUM_WDTH_LONG-1:0]         I27be9ab07b6db7a211f0f2fc97fae8866b139ac8b76fb72d5b207866ef5dc538;
reg         [MAX_SUM_WDTH_LONG-1:0]         I9c74de21b57f62df69930fb5dba0c0a81dcd57ea06cbcdd3e1dcbc9077a7396e;
reg         [MAX_SUM_WDTH_LONG-1:0]         I6a231da6c84868f89279c52b472159f3f28b097d98b55fa959cf8b65bd7357b7;
reg         [ 0:0]                   I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f;
reg         [MAX_SUM_WDTH_LONG-1:0]         I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d28f08decf784d91ab2c0bb92cb9b95d798ec46ff319335f399bf55f24ca0c9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2ce9a3e0eb6568348a715f3d26e23ff836ca88d2a48d62beb9b06f46ec986df3;
reg         [MAX_SUM_WDTH_LONG-1:0]         If13322a1bb24c2938298fda568b15f72bd6258fa12017507e5c8c34aa31969d9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifb7752c1ee4d32c33015b0978e0bbc378b26a7467ea1c4983c2700f2372de3af;
reg         [ 0:0]                   I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421;
reg         [MAX_SUM_WDTH_LONG-1:0]         I29cab53a69f72bbcf1812b364c9d4aca2dd9ca2159114ba63770ba7bf154c032;
reg         [MAX_SUM_WDTH_LONG-1:0]         I98b2432228e13880d555f5f32794fec8e0c4b85eb066e597f61dfae883cada43;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51bb519f0f46144969987729901cfa4e19f29f9703a5c2129ced5c6bf9c4531c;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3865ea29a692b3a2567934ed101bc0dc34c941c7fa7c6fa6bd04a0670fea64c9;
reg         [ 0:0]                   I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifc0ce7736e9c48c2d5e0e39ccf90c85218bd13a7e93695a158971e86e560a9b5;
reg         [MAX_SUM_WDTH_LONG-1:0]         If5eeb2eea320a2012569a69de41e3e45dbf74bd9e8330a3c0a1b6fefc8994f01;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iacf07c5d8bc2563c377f66311c807d18c4cae1b4af253c3c55cb940c9d49257b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0c2168302de09a1bb09056d8e2f6cf9a4191a5151b99efe57fe8fec69e2c349c;
reg         [ 0:0]                   I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7aa29eeabf60e0de8e049cc83631713eecc92a33b00ab66889601b65a8584021;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib7cd9e5a80b095f4c71eb6005d588f15ea498ecbf90748e128e42c0feee08dbe;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ia9f187fb62e136eb42c8ab963813a504fbd8ed5f7390f608f923c3d5f8853a05;
reg         [MAX_SUM_WDTH_LONG-1:0]         I482ab667b97b8e90796abc13f93d317377f279dcbd4c9699b5bf776cca58e12d;
reg         [ 0:0]                   Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic59104908c4c5eb1da72d1f877270cc3a75512d885653de8de2aaa5bc050ae87;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2e28e3dc68c6c9d929ff4706e92b74d5b52de590d44dc846007d24a929cb60c9;
reg         [MAX_SUM_WDTH_LONG-1:0]         I29c2a83008b667730e3fa038ef10d5c8c989348c36320071fe5a93d15a608d65;
reg         [MAX_SUM_WDTH_LONG-1:0]         I7e9eb2043321328a9ced3e4d319e6963e60ba7928bec6115527f55f70cbb8db1;
reg         [ 0:0]                   I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987;
reg         [MAX_SUM_WDTH_LONG-1:0]         If70d53608aa2878766b77726f3e0f650f572b7e89ea4df1a4504306868cc44be;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifb7ec2a54d000887851d37b4b0f1be483d3caef91a4d07b19edbc19995fc77c4;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib24004e855a53de1330e5ec4126e220205ba20169ae9ee4ec34135db389763bc;
reg         [MAX_SUM_WDTH_LONG-1:0]         If81c09fd3901cbccd2410864fc3e2d7087c400fab7cb319f6de0e030d706dc1b;
reg         [ 0:0]                   I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3ec9f20d41034d8e73b2a9210188b70e7b2c68e62b25fcb5f140598043681a6a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I21d1d0816fb6a0c22f2e850ac9a2d9d1f582c218de0eae741d1c9916ad2bc5f9;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iedde649e1098e7cafbda605e624786ca97ff3b6e68c7ee8be00b813d8ba5521a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iee58ae84679865c9bfa421865961b359874636d1a9a6a85bda680627cf00cd2f;
reg         [ 0:0]                   I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96;
reg         [MAX_SUM_WDTH_LONG-1:0]         I00a07c03491a1f197d8ff004b3a7816850d0cd272e4ab9dd574ed104f730500a;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0fa68b59aa1d936947137ecb31171e019a59aeadc82044e25faf04536b89d301;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4e3ea3d10bfb18320ffcdf21e5b7f279ab94cada35ceb624c8bbb1f5fed062ae;
reg         [MAX_SUM_WDTH_LONG-1:0]         I37b48c08b0e188a8ae4c35cbe94bedbc2be0d8ccfe5dc8199fab4bf3a5c2b4c2;
reg         [ 0:0]                   I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d;
reg         [MAX_SUM_WDTH_LONG-1:0]         I311137155e974b61171f0b9f85b3380cf230186a137daeece322108026a54fb4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I86d7cfde239760ee206e636d19402cb5decc9d170670b47874bb6e51950e797a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Icce39cddc9b07a5408d7b7cc73a0aee0ba96dd9b59ccb5f9da245a8115636e81;
reg         [MAX_SUM_WDTH_LONG-1:0]         If0c116c5bb5aa35db83ca1f71a49e32a260c13ce39a02cf3b683d3cebcdd412e;
reg         [ 0:0]                   I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5;
reg         [MAX_SUM_WDTH_LONG-1:0]         I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc1d7004fdb14267759bb0b179acbaf24853d6b0efe051dfd48de07495940dca;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib01b562cc42dd79d910091cbfd3ecb8cd0b386f396893baaee60076b8c04f906;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ib1b3ee65ad4ddc6d66bedc912f129d315715913cb1517e24bfec0669f2b3ea04;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic2d2abe362d0a76e22e5bf3d902cf55d1091dce5ff18a17ec2b51dac09d2601d;
reg         [ 0:0]                   I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18;
reg         [MAX_SUM_WDTH_LONG-1:0]         I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic667337f6e8f713aef676104d2c4af6a634660e47835d615bb7b74af34c3e979;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic0a75ab618b9081cfdcd40620ad47ce4da348de800f33a88cae7bcee7ec46f3a;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie6e50cae460faffae965f9ee7bcde9b12d5efb54a7d8f03d45a34cd1cf6e36d7;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iac4ccc031aca350afe26f7ca6b09c8d4c124dbec5e0e705ba473f4c2834952f9;
reg         [ 0:0]                   I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481;
reg         [MAX_SUM_WDTH_LONG-1:0]         Iedc1f868c50438002a4d97e96e0dac521014321ddc6d61e49b5eab223b997086;
reg         [MAX_SUM_WDTH_LONG-1:0]         I18cd7259e4f753e93903dc1031fc51c25f000a37959e858574b79394f1dff508;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ie9395076cd1821b1a6cd391c4ce616cdbb0bc759a2a9f3a7ba32ec60b9c6015e;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic30aa34e60dfa155b665def463cf115fe22112f358895a836b4179f33160134d;
reg         [ 0:0]                   Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I577e72330edc830f5735c0ed269566f49c7fb3c4d196d3742fd1cf3c66cfcc95;
reg         [MAX_SUM_WDTH_LONG-1:0]         I08b93985c2d4ce016468d10b7f0187ec3cd8a803308f2333bd361255e00977b6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Idf041d85612e43dacf84491d005b30e93873e31c1b6e56df2e0ca7f0babdc5a6;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic9eb7815de9b84b1a3763dbf218de5d7d844ca252937b7685b20015bad378659;
reg         [ 0:0]                   I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205;
reg         [MAX_SUM_WDTH_LONG-1:0]         I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ifa413778a53ec09ef3948f1ff255ab5b73d9243508614c057c59a153ad5289ea;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibc8a3b5a652d7343e1696747ac66770452a464ae8bbdd112799540acd80824d8;
reg         [MAX_SUM_WDTH_LONG-1:0]         I3e50387897ad4d501a045ec8c1ed398fd84ff960cca94f41bd41fcd6462783bb;
reg         [MAX_SUM_WDTH_LONG-1:0]         I25ddd61dbf2b3f1b4024d769f62e690493ca0fdd01b3550226c9661ed9230fe1;
reg         [ 0:0]                   Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884;
reg         [MAX_SUM_WDTH_LONG-1:0]         I4dee2f1c5fecf86cc83b723fe96caccffdc564334698e43f9c04db5a25afc978;
reg         [MAX_SUM_WDTH_LONG-1:0]         Ibdf4b745b03013632bc0ac5142c9dfb98f197c78e95b71ce1074f84a5b5c96b4;
reg         [MAX_SUM_WDTH_LONG-1:0]         I0adfd7bea27acb0ef24fc07bb0649de5bc0ce7dca6226beef48e27cea9aa4df0;
reg         [MAX_SUM_WDTH_LONG-1:0]         I870372f2d3e9fcc2db983123cb83c7a6f1b5e9f022d915d5534425322e8957a8;

reg  [SUM_LEN-1:0]                         I93c1856af28a13c1890271dc68b7b6cae884657bece4e0d452fce3ef922a9c12;
reg  [SUM_LEN-1:0]                         Id76ecc370ac753fefd8cbdfb525a5868396234d646214915a49d70ad4cf925a7;
reg  [SUM_LEN-1:0]                         Idd909220a9540c998e23f1b06cfca187d9d83bc0673aeafbd0ed6c20c9d39f4d;
reg  [SUM_LEN-1:0]                         Iba7e42dfe0894a09d968f0190d344d90387e96a8048a01fbb5d05c15452f6ce3;

localparam I7c47889d7eda9026cce141952f929eab96cdb46806801c429c11b094be47b7b4 = 50;

reg [MAX_SUM_WDTH_LONG-1:0]    I7bd679f7d7da9dc0742c725247978f1c14611083c7de896c4c2de108c6766fb9;
reg [MAX_SUM_WDTH_LONG-1:0]    I11abd59187e2db0058526cb1ea58af9061d439139fa151aaa74184499fcfd24d;
reg [MAX_SUM_WDTH_LONG-1:0]    I950415762b14dbc0817ccfb0d09d95d700be57ecc9f8011c6163f84336da6e43;
reg [MAX_SUM_WDTH_LONG-1:0]    I9841a5dd86a1b359b25fb293e74cfbd88b34e11f22bb61170ecc921048620dc9;
reg [MAX_SUM_WDTH_LONG-1:0]    I4c8a0d23fea7158b5e99eea187df1d25395edf7df1db8482b41dab7a8bc25030;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia6f33a5c8baa6ea053642148b8e414d0b9d17a66f4e71f6e44e1f6c6e3e535ba;
reg [MAX_SUM_WDTH_LONG-1:0]    Id7d51984757deb5794eccbf50647e7535041a18dc506aa16b4ba0ad36bc66b0c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib8b4f3fbd26b51974ecee1565c3d0c8fa7abd94e467a7369a62ceafa7ea5ddaf;
reg [MAX_SUM_WDTH_LONG-1:0]    If787a878ae1cab622e44a13190d301d15d0c7ed9271dc50e997c926071f1cd02;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifb337611e63cb9cee9828aa75fcb6d978249e65bcc8770d51fb4dd1644c96a86;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic3ea8409cfacf50e41b97c65b0440348d06b8f196001ba1fda6348071b47dd23;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia49277306313784711d5d8ff63e6a0a77d3fbae050dc1089c734c826be497dcc;
reg [MAX_SUM_WDTH_LONG-1:0]    I13f5f01dccbdf3df23c5bf603a9657e161c1e2368cb5cb48b212231d2fba7794;
reg [MAX_SUM_WDTH_LONG-1:0]    I7c6ea337917ea8eb0696c514db7ffb66719763162bdd0b7e0ac764c1ae63d24b;
reg [MAX_SUM_WDTH_LONG-1:0]    I8fe688adfc161cafc0777f3c3ac9ae27372603ec55cb3865f90f38f9dbb59439;
reg [MAX_SUM_WDTH_LONG-1:0]    If7c696b260799e0ccd86bb377086dd1be59c9d94754dc52605d659391439d3d5;
reg [MAX_SUM_WDTH_LONG-1:0]    I16ef3abe43350c9096f6c7e597c48fc86ed26a073055b7bcd696c34676529372;
reg [MAX_SUM_WDTH_LONG-1:0]    I2f4a0e474435a97fa5d2d056d9de566288c0624cb094d71685934475b58572f1;
reg [MAX_SUM_WDTH_LONG-1:0]    I554ab27e696a028f48da8ad39e2db6668b57ff692603a9562cd7e8780bfa491d;
reg [MAX_SUM_WDTH_LONG-1:0]    I78d7fbedde9ab5751194c52134dec1b83ea8d48c4ad77c0b3eb952143612ab71;
reg [MAX_SUM_WDTH_LONG-1:0]    I9b494d3414d329e4419da30566795e7b36627870c521c463cefbeb7b48196d3c;
reg [MAX_SUM_WDTH_LONG-1:0]    I8060bc4cf825f705f2218152b6a7a8600692076ba01123cae35feec231f128dc;
reg [MAX_SUM_WDTH_LONG-1:0]    I435bc44b4b8aac5fe9ba3c30a74d51a42250154c16d5750e075057d1743ffd69;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc131936849b96a3bcc7bed4c38ebe94d51c56feb4e96d25dfbbcc3670568a16;
reg [MAX_SUM_WDTH_LONG-1:0]    I6d0d8fc19811812bc80267dd50fc4742e9efceded7a9428707fac605fac90368;
reg [MAX_SUM_WDTH_LONG-1:0]    I15e7d6b702e93b31ac4e46f9ba4cf63da33641629eb9cd414d1e2c8cf54b750f;
reg [MAX_SUM_WDTH_LONG-1:0]    I26e6175466ec922073d5092cb4168f87cd1289008e4b99400c5b6c2fec3eaf5b;
reg [MAX_SUM_WDTH_LONG-1:0]    I97449b979933d41c6555a04ba5ba6cae73e44b040387a504f6f7e2ecb763ad08;
reg [MAX_SUM_WDTH_LONG-1:0]    I272bc7cf289752b36b9811d4ec63f5c17cb40399f39607b00ba51817fad59e1b;
reg [MAX_SUM_WDTH_LONG-1:0]    Iff259e6b8d77d06a8354c4d1662328284ede633f1ca4ec4731dcdae94e869f66;
reg [MAX_SUM_WDTH_LONG-1:0]    If4cdb00eb64cb9e80d78f3dedd797796f44f471b76f5ea3ddbc6f8521257e4c9;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac435cdd22e5425837ad24bd6141cb357c302af7ee7637e1cc2ac25474cf7506;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic9e13fe7c29048953ae3698eb5d214d6b71367a78bf1042dd6b58064a6cc596d;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf9f5e717c65afd1b3bbc3d6c1bd960155773ec7790543f56c86637a891decd9;
reg [MAX_SUM_WDTH_LONG-1:0]    Ife767fdd58724398b336a58803ca328013f3a8228ede0cf108dcae054001de56;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic55bde9a87033c380a5cfe5736d205c15099a2f2cf440f88472d7f6e65d360e1;
reg [MAX_SUM_WDTH_LONG-1:0]    I3af3a7e6138910d118e49b29a6de8bb8e6fbd1cfe13549eb0feea6cd07e6865c;
reg [MAX_SUM_WDTH_LONG-1:0]    I55e293b2d9539b16ee0f135097b8ec02fc9af54fc96ec3a3058af417b0d04e48;
reg [MAX_SUM_WDTH_LONG-1:0]    I3088ff7517eebe83fe5804308d22b8c6190077f576f2e680848092e21116b94a;
reg [MAX_SUM_WDTH_LONG-1:0]    I8de3f6aec12696eef7d069510ff25e6e620fc4fdde5f92923a707116da636284;
reg [MAX_SUM_WDTH_LONG-1:0]    I6996b52f42eb9075a634fcdb07fafaf45c5aa99193446869751c4859e7c1f963;
reg [MAX_SUM_WDTH_LONG-1:0]    I3fe543ea18333fd169c6d6e692a5b42232e8abd2b14072a4daba9bacbe921d2f;
reg [MAX_SUM_WDTH_LONG-1:0]    I29d04420073229582b38d6b3f7d9d638351e92073269d5528b09b080e5fd5670;
reg [MAX_SUM_WDTH_LONG-1:0]    I8090d844610f0d62cc25a9c72c2d76d9d6783a067de9c9ea9d5a1f5c48744c70;
reg [MAX_SUM_WDTH_LONG-1:0]    Id60b432b19836d2e0919dc2e0201d162d7446434080aff7165fb949aba097f7b;
reg [MAX_SUM_WDTH_LONG-1:0]    I96248ed668211f13555b4a086e7534b958b901242794b9978d673726d56286e0;
reg [MAX_SUM_WDTH_LONG-1:0]    I78023336da442165a8be56b4ebf7b41f4bb48bbc2b05c308dcd344c8f36c476a;
reg [MAX_SUM_WDTH_LONG-1:0]    I05a7291b0f3122dd9941bdd5ce72362b3b0b1803abb126606c82744979184be8;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia2952eb350b07a9cd76752e1a5f76814ed095eb0ee2a284f221b1c74e38d822e;
reg [MAX_SUM_WDTH_LONG-1:0]    I9f0d592f1a57b1d3e2c206ffe5a79185253205dfe7b20be53091145aa16f9719;
reg [MAX_SUM_WDTH_LONG-1:0]    I62d2fe36d10e598efb7f38f4f57e4511d08c366d7df7f51bfbc63eaaf216035c;
reg [MAX_SUM_WDTH_LONG-1:0]    Iec33764f14e5b0a736fa76a2313325240a520c065b59c6cdd0f2fc5dc36a975b;
reg [MAX_SUM_WDTH_LONG-1:0]    I9e89eff507c5a2386876f56afb505a22f00d8c0f8a32635a00501ef8d56ecc6d;
reg [MAX_SUM_WDTH_LONG-1:0]    I0d6546f557347e1d72c176a40dcb077c9c4c78ed89975154f5bbb3875eb1131d;
reg [MAX_SUM_WDTH_LONG-1:0]    Idc5ae39b0c3c764ed6d9b7859b7627b97e24c2b4df7d97229a88cfc0c22ccd87;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibf4bbd894f269bd6e6eaf9511141b91ac61b5dd3e77b4ffd07aa88474f251ddc;
reg [MAX_SUM_WDTH_LONG-1:0]    I26ad8ce808bb26201de4f63afd861583af9abc55c7623bf15bd1808c0b0c2be4;
reg [MAX_SUM_WDTH_LONG-1:0]    Icbbddd7f07e1deff7aacc0e96a33556b62ba127dce877dea351b421ac8d00313;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib87cc4d1070a195aa8118b92d29d7c836685de2e44ba1b21388677c8e8a5fb25;
reg [MAX_SUM_WDTH_LONG-1:0]    I8dc734304648fe3fba1dc7108e8697cb88b61a2ffa704491b2b9df8cc8354825;
reg [MAX_SUM_WDTH_LONG-1:0]    I830406b0cd2e64515811ab932e9ce01d413f0a68ab7939a2fa14e4eee7d04a5b;
reg [MAX_SUM_WDTH_LONG-1:0]    I113d1ff61779dda7e1209787ba652b8b332fc5811cdc0aae65a304aa89d56766;
reg [MAX_SUM_WDTH_LONG-1:0]    If50a43f14a383995b16d784cc119d01749fd30928019bea1b7aba0039c4c350c;
reg [MAX_SUM_WDTH_LONG-1:0]    I7dd3baf838ce22ecec10d3c1a3d0dd16582497f9e447038aa46bfd49571fcb4b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia55512c30a26e336794d389f3700b9153cea83619467b731571ba72a3a9374bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I799968e729d7842ce09a838203458d89b96fe9d2d7a5de0cbac32eefbf834898;
reg [MAX_SUM_WDTH_LONG-1:0]    I2e17b8ef0d25ba5beb474e7007ce1fe5f99f6f7cbf24e5241761880a551f3c12;
reg [MAX_SUM_WDTH_LONG-1:0]    I7cc2cdc76a638cf4fabcdbd60142d7e4fa11f11486c85b7add7d4f9ba16042c5;
reg [MAX_SUM_WDTH_LONG-1:0]    I03527e99f5c488d7864664f339e2094fced797e4b46101f3c2bbe0b892c2d299;
reg [MAX_SUM_WDTH_LONG-1:0]    I9c110ac43d6a359d54082ce347cfc9885dba985b743aeb66bf25962b4539a6e9;
reg [MAX_SUM_WDTH_LONG-1:0]    I44089ced0a31e79af650baaa02274890b1f60ac7398745a0e4da4b2242f849c7;
reg [MAX_SUM_WDTH_LONG-1:0]    I1308b215c5082a0407de73f2273fc035460ca21b553479402290c244cdedad76;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic0561c97824b9d5b0d84c33cd05cd4f95b9cacab06eeb5e022b0cecd043c6a75;
reg [MAX_SUM_WDTH_LONG-1:0]    I533b2cd0b272eac7c3f9005cc355cf85ce73803134a0fe0ec194628c3af0ed91;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie282d05ceadb0d075cca024b7311a5e477e903295d7928735a3c338287734846;
reg [MAX_SUM_WDTH_LONG-1:0]    Id8832e8e711bb3e7fe9136084b9832a2677803cabec7f2469144eb3b6d4ee3ae;
reg [MAX_SUM_WDTH_LONG-1:0]    Icefdcbf9ca1f8e02b93f295ed8dbc43258b29cbc0cdf9c9ed5fa60117263d502;
reg [MAX_SUM_WDTH_LONG-1:0]    Iba1a21e329197ff5e399aca440cec6d6bd3d9593c332cfcba84d52d541ff1ae0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5a93c88521f26a686316f032821a4e9540fdd8e93570ff35437df7522d34ab7;
reg [MAX_SUM_WDTH_LONG-1:0]    I91c159ee16a42dcacaebf8cdac4c59d45d2e93735cffd86620ffaf2b859c8795;
reg [MAX_SUM_WDTH_LONG-1:0]    If7fb04f8e3e8eaef8fcc0486d12d1e37a887bcdecb366c1e8b53a3e1cce0637f;
reg [MAX_SUM_WDTH_LONG-1:0]    I6dd215113f113a81bfa59464b587ae7c95f02c1461664fdb818ce751c240b96e;
reg [MAX_SUM_WDTH_LONG-1:0]    I08384d6ff32b692ca710ac4170d45cb5d2e2df509bbc473af140dc50f51fe46f;
reg [MAX_SUM_WDTH_LONG-1:0]    I6159ddc580c73acd6e2391f4c6cd9989ebaa8947db61972e4fb97f1e12efd17b;
reg [MAX_SUM_WDTH_LONG-1:0]    I88f1c4536adedb4ffea1b595f5fa753329c4aa2187a3245269734a18a122e189;
reg [MAX_SUM_WDTH_LONG-1:0]    I6f52a21dd933b23b7565abd508c69070b8cf652dc313689f62c7f04d7acb934b;
reg [MAX_SUM_WDTH_LONG-1:0]    I0421a9a7aa72d6f574071ffb4c65878f997e6dc2b605f0d8b351358b08c47ce3;
reg [MAX_SUM_WDTH_LONG-1:0]    I60b41ade4579462091cc59f1faf9f78f236a3bef12f893facebdf8e6b00096e7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5d526172ae46c2a06c11e15361cb13141d0ba754320f60ce6bcd97a9e495221;
reg [MAX_SUM_WDTH_LONG-1:0]    I7def9ddb7ba2e414a44523f17bbff45806f0100ef624a52e91b03022877a7771;
reg [MAX_SUM_WDTH_LONG-1:0]    I305dec30cf8323b9af4b0a6d285a31b3f5afb2e79c1a2ea77ce70a4409a7c765;
reg [MAX_SUM_WDTH_LONG-1:0]    I8ae4ec097c879009d8316e76b0a2ff9f4228310728d8b4dc196543a3976d26e3;
reg [MAX_SUM_WDTH_LONG-1:0]    I123e1ea1b1588abf2d5d4ede7027783bfb20d60ce3fdf365b86c9f5c84956a72;
reg [MAX_SUM_WDTH_LONG-1:0]    Id9d184571e769ba27b0a5a10807ba8da3e6ba57ed7d66aad1cd984ddf5cbcbd0;
reg [MAX_SUM_WDTH_LONG-1:0]    I05782c612bec6ce9c2707bd6cb6efd55e1da4d234be502ac88cd02453c61ca60;
reg [MAX_SUM_WDTH_LONG-1:0]    I0549cd0fd3abf1658d503a09b0baa63d09b1411eaa524e56fd30b12f8498e549;
reg [MAX_SUM_WDTH_LONG-1:0]    I19123fb30bb6e02a13f39e3e96af227e63abb1351e53cbb91b8d9a79be96053f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5d22b614e704f01c688034adcd70603b8e69658cb66c96fe3ea76bdb323c222;
reg [MAX_SUM_WDTH_LONG-1:0]    I886fbef883afc3146952de2fc934131aeb38bc2134c096497981d303594f1f37;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib897fb3696e7d68b81ff3c1573f5cc234d32e10d066864ec203487a8e56f4ece;
reg [MAX_SUM_WDTH_LONG-1:0]    I5bb2c70350634acbcf64debae260225ea2ef5b67ce5d03f38d56d3db9de687f5;
reg [MAX_SUM_WDTH_LONG-1:0]    If81604260c143a45d248461563d4d94edd94bb71d791a637dcd30c5c0cbbb965;
reg [MAX_SUM_WDTH_LONG-1:0]    I0806d1e2ea1771b325ea80b71fe9223f495a3831a560f579401b4e94b6ed172a;
reg [MAX_SUM_WDTH_LONG-1:0]    I9075819cc111daeabcc2ddedb4a4297b1a42ceac8b93213f7f76d0fe87c8c275;
reg [MAX_SUM_WDTH_LONG-1:0]    I317bde7e15c3a4d1456e9653a45d4d574509cca539be5c064af2ea89db634f45;
reg [MAX_SUM_WDTH_LONG-1:0]    Ice9dcc5d9ccd6caf90dda22be9ce113c53c7eb492cfd5e0b237da4f92aac2d7f;
reg [MAX_SUM_WDTH_LONG-1:0]    I54b0290e037c2111cfef49e6b33d9a3fbe3e85f8fa8a5c707832cb5477f5c0f1;
reg [MAX_SUM_WDTH_LONG-1:0]    I7925970ac367f8374fe02f6e4c8c339c58808928696f0acaf85d96fb3f202f00;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib398240cd12e68fb5b3ad4842123a4a16f27cfcae3db8bf1f38de24b82e272aa;
reg [MAX_SUM_WDTH_LONG-1:0]    I9df56fb9c7b812f3ca5949962100efeb5889d69ff60754cb4eb3e0dd18376d45;
reg [MAX_SUM_WDTH_LONG-1:0]    I93f4f945a6dfc45c0a002e0bd9251f56c68570c71e862e222a853f8855fb1165;
reg [MAX_SUM_WDTH_LONG-1:0]    Idf3bd173aa5e956e898d5800f3317a1ef71e334901db42b94f9c6aa41c87c2b8;
reg [MAX_SUM_WDTH_LONG-1:0]    I7b25bf7d9020a7dacab3d15cd039a86780e41ed33520f5272ee788252efd1b9c;
reg [MAX_SUM_WDTH_LONG-1:0]    Idde70a085816497aa92518899b882b67eb7989897509c445847e24204f5e978d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ied43949ed7bc9c0c92af912b9e283a3e674d42242e0fe8e3d9132738d512fd23;
reg [MAX_SUM_WDTH_LONG-1:0]    I18e4b7dc3295cc6f5968878bde7abe5447cebc77dce83fce47db55be2237efc9;
reg [MAX_SUM_WDTH_LONG-1:0]    I4a91f2655f96c11b03fce33601bc8f71a0fef4dc1782f7158126cd8cc5a1d690;
reg [MAX_SUM_WDTH_LONG-1:0]    I343c495ca033301298c16cbb81a11a7f9d50dfa8b93ea9226caa182c6fae8737;
reg [MAX_SUM_WDTH_LONG-1:0]    I451de528c384521cbb78ae32b3d4640b0cb8d507c10e11ff59a74a9caadd2117;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieca82bcdc6bd68dc2a28a3b203d8adaa09f89fbf0df6cacd8656b54b141d758a;
reg [MAX_SUM_WDTH_LONG-1:0]    I876c143c75e838720b2a1ee393f5da5ba08822ea13fa1ff459d68d7b0c0e5cd6;
reg [MAX_SUM_WDTH_LONG-1:0]    I88e5fe043e16a274d915245b02d2094d05fb7710f6078dd6b33c2a21676200c1;
reg [MAX_SUM_WDTH_LONG-1:0]    I101eb18f34badddefbdefe0c2448e2a8a243e4803ef3244b25365881bf227145;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia249a4e7b5c5f1f4458d969c346e560a28969f33c9b0371c6bb21776d319afcf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifd8d2fce7b2a1f0fa487e5be6c007a21b5af1d79da5447d461cd37c189e43561;
reg [MAX_SUM_WDTH_LONG-1:0]    I840289556d82218416d7f8652d40586181f7b4ecedd132450594aac1bc47a081;
reg [MAX_SUM_WDTH_LONG-1:0]    I98ee0d4994c76a87aaef2967ab6cb88af05ab0a7972d2dedbf115ec19c426fa0;
reg [MAX_SUM_WDTH_LONG-1:0]    I953a4a4cbd4e6c0ccf4880cec5c947f86d6542f9a7f125d7c8cd71f8665b9ddb;
reg [MAX_SUM_WDTH_LONG-1:0]    I908d977677aa9b15536027b54cf497ddb8741b339748986180944418fd848448;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic0fd25473d5639721dddea090dc037e39e4a0c08776c0a343408dfcfc402fa99;
reg [MAX_SUM_WDTH_LONG-1:0]    I46777db6f6f68d76ef34c4a9c585ac04e8a978663fecf72d2dbaea3287dfea2d;
reg [MAX_SUM_WDTH_LONG-1:0]    I4a4338f7d9bbbf60ef4dc6e821d22619911e41300b49e83d57a0a959218a05ae;
reg [MAX_SUM_WDTH_LONG-1:0]    I5cbb1dce1049c737c8e052dd6b84121d353e3ee02202bcb8e5fa27261029c96d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib4d2bee91a2ab56208d3d1f484e63f085a162ab9d482690dd3c5891a2a34d808;
reg [MAX_SUM_WDTH_LONG-1:0]    Icb9b19c9fb878af708bd3b433b656104d0f1ae64cb5d5a3f8dfbac08da1fdec6;
reg [MAX_SUM_WDTH_LONG-1:0]    I9989d555a1c808f108dd152608d93b00d7a396de9492733ffd5165700c869840;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibc813c005ecf7c077ea48779116cce31bffebb300fab262a78d166c4e270e3b0;
reg [MAX_SUM_WDTH_LONG-1:0]    I58ea58692cbfa8283ab19d6e609fe472aeb9da51d3f3616a9069eacfb18b0bf7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib2fff9999fc00e81b173cdaa0737f3e4f711ccd0034a6611e0e9111acff3893f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia441ac067e28123cc7cd9d005d0f5a1628da5628d4473db60d61b85c61e8d9b1;
reg [MAX_SUM_WDTH_LONG-1:0]    I58aad5a5682b85bf58d67b9b00883f015e4093979fae9138f7dcd813618e26dd;
reg [MAX_SUM_WDTH_LONG-1:0]    I511b38f7ea620301cc3bfa759ab56a2dac9061fc83fb1281673a6cf276abcabf;
reg [MAX_SUM_WDTH_LONG-1:0]    I0b2c4982c217189306b4f5d3bace84daaa25f2bcd089f5de092f9a7900106c6c;
reg [MAX_SUM_WDTH_LONG-1:0]    I3dacdb67f2492ed12375b671dc593349c75562e936401def91b4391c153fa572;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibba131ee71ced96650ce76aa4695641a089046f8b8345ba312d6868dfbfb2787;
reg [MAX_SUM_WDTH_LONG-1:0]    I82a2a0149ccdf627e13b7d422945e626fa268c22b3c30bbaadd0a8de14ddcf32;
reg [MAX_SUM_WDTH_LONG-1:0]    I7efedd1a063df95cac921f7cea9ceea1ddd1afd3a70289c50ea2a4807310518b;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib91519b86b75cae1ba5b32dc531cae021a01350f4e184d39373bf5553f89a7f8;
reg [MAX_SUM_WDTH_LONG-1:0]    I58cee4a472b2fa2f17266cd6ab55d475f304bbee835aac31ac7879d77b8a23eb;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic4e32c1234be0a530c66106794dc1114e4c88611be106ffde42a7ae486560ae5;
reg [MAX_SUM_WDTH_LONG-1:0]    Id32cba1cfd5a10024378db5089213ad668054033f8614d1ae09b83fd483a25de;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib0978aef78ec9b21853831a81aac1d87a2410594c7839432302eb5fa99a4c0ca;
reg [MAX_SUM_WDTH_LONG-1:0]    I257c396883faa57c509e7257bed0829f9ca51f30a1004ce730d48e1e5b40c0ff;
reg [MAX_SUM_WDTH_LONG-1:0]    Idaa2e762bb01a89e36234967b22cc76cf290937df9295939bb4c4ad08cb8413f;
reg [MAX_SUM_WDTH_LONG-1:0]    I9d7b0f41f5cd73f907351990b23117fcaae4302a36d194e6953b54d40361f8fe;
reg [MAX_SUM_WDTH_LONG-1:0]    I8d463b693ea969ef3023c411c0c9a1fbc49f81d348282c031b963bd8ce0527a3;
reg [MAX_SUM_WDTH_LONG-1:0]    I6822ca486e86051ea654b41b63bfefc12a2218ec87a88d8b5acc3e3c8a604c94;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie515c89eac4b602d36f70f52a3fd62fee155da2eafac9c1b14bf1917b62bab44;
reg [MAX_SUM_WDTH_LONG-1:0]    I3464299c3a5abaf050c7176e4c0e17ade3cd5d6d86e82addf3e12d662def2b86;
reg [MAX_SUM_WDTH_LONG-1:0]    Iefd5db28023cae3483fe3f0f1dcd5e302d642a0b5750cfa9940a9a8d6326cdb8;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic98b2baa4c4b3d4541ae5e7f9ae0b032d4dee98ebd73901690f561438ecfe5ce;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie6d2cd42fa78c1cbf17c7f18dfb4c0cc5f79f1fb0bda02dc92192252f99dd047;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibbcaf468c4ded9be4d2d82d059bfad5174f330444c98aadb71831769a32f70c2;
reg [MAX_SUM_WDTH_LONG-1:0]    I17e36eac60eec64de05cb738d1e6055086891ee6fd7d8fb300df4f98a3405276;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib8956dcf80473ed75d04e9fcc74400f54ee0b840fce7500bcd68ea6dac6d4473;
reg [MAX_SUM_WDTH_LONG-1:0]    I873ab672a8d92c69b75cd8e627aaec129f1cd371c9f863a6bf88e3965909a6d6;
reg [MAX_SUM_WDTH_LONG-1:0]    I206a4b82a444ed76c846a17eccf6c9ad62c42263b472949cc97f838f6a416073;
reg [MAX_SUM_WDTH_LONG-1:0]    I428333658d20f4417e24a58fe364d5a647332ef76ecb7f15d83dcccf1aeb3d11;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc4886636576352e5307fb1fefefded0d693fd059a3fcdd6b4c9dbab1b908114;
reg [MAX_SUM_WDTH_LONG-1:0]    I18886d5e45fe8011ebcf9a20aebf875a01f1b793a54ccefdbe44a896e92cb0db;
reg [MAX_SUM_WDTH_LONG-1:0]    Iecd27d9347b5f52e83b7d0fbf7e51de4a3711cbece5ee265b12663b77b58914b;
reg [MAX_SUM_WDTH_LONG-1:0]    I5246ce1dc41e20a5e4e3312a997e8c5be2d733f0cc95f74caa7e668f9ad2f1d6;
reg [MAX_SUM_WDTH_LONG-1:0]    I668775bd016b2384bb3d1cb0a1e89a76d2af15b2307cc6a5d2e0d6c699b02544;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaad1ab5e7603d5441b228c5e899eea7781b6f486b836a7b662f38ea832c1b8fa;
reg [MAX_SUM_WDTH_LONG-1:0]    I9d56c14b3465733b5c5fbff528a7a7d85c918a857257ba8e302ae84a0f4734de;
reg [MAX_SUM_WDTH_LONG-1:0]    I7ac4d72123feb2b9af1a6c3da5adba445042363194ef471c8761e289178d0253;
reg [MAX_SUM_WDTH_LONG-1:0]    I7addf7487638274202ddfd183ba052556f89f82da9e873224c5dddf27d2d5a66;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib0de9295b071389ca7b6bd34f7c9371614337b0be04ccd9ab9819a8e39ade463;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf6cba7551eee2b4d2b53263af6fc190558f5b29af52c060adf5bc9116d56341;
reg [MAX_SUM_WDTH_LONG-1:0]    I01a734e70411ca4d260541915dfb0aa0eccbb88be6043a4a46e412d3b9f1e778;
reg [MAX_SUM_WDTH_LONG-1:0]    I04257aade4809f3b60c5cd618c5a29008d1b3d7041330bd5c8db7df720da3694;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib33ee0ec338d1389ec9010793383d24de32231284e86a9b03fd2902743dc8a00;
reg [MAX_SUM_WDTH_LONG-1:0]    Iecf3e0156bbf76dff96948ab7bf67772773b6bd62bd0e0fbc86a6eea8b05d4e1;
reg [MAX_SUM_WDTH_LONG-1:0]    I80c4eccc6e6be84f8936ed3e9a9457a862eca015298ba2db70745f25a65a6571;
reg [MAX_SUM_WDTH_LONG-1:0]    I7355df30b826dd16e0f1fe3be878df80c2ca672dfd1392e2a81ac34fa3df69ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I8f671fbd5e9e240cc2f3a9c60c1340fb4bea46c25cda7ea5e42c7ca0c2360bb5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie3806d0fc4177d813aade41ad46537a9a335516135161cb2ef18ce822cb301aa;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e8e17839b8f0cf30290c33a60662c784f062950716903854e36856a58f909b7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic46278073f42d4eba79499cd6293cfcb33a74310e7b2ed4bff06f5cc63dc9ebd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib1101385e86160606eeb12ff49ee86ca465f227b19c9bcad4811c6a0183c0ddc;
reg [MAX_SUM_WDTH_LONG-1:0]    I4bfb42a957ed14280a129921d4d635017b23dab77b121f51abcc5e738114e446;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie11729721562e4a52a189a242aba934be636847d35de867cf00d26690c69abd0;
reg [MAX_SUM_WDTH_LONG-1:0]    I84cdf374f692a63dab22cd91edd4f71e1aff29b51b06f0bca914f92407bea09d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia2aece9bdb39e997b99e491171667091adbee475ea9b1c372ebbec109f9f714f;
reg [MAX_SUM_WDTH_LONG-1:0]    Iabfa5de761b3413904b919f913ed73bf27f5249b7dc6bf8471a23f06a30431e1;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf6fe11d7e6948c0bdb9cd50a0135c3b0fac213aef728b8a6555b7601c51cb7e;
reg [MAX_SUM_WDTH_LONG-1:0]    Idf57b2bf209c68bfc70fe2759595334fabe3d50dcfc4fef8637586c6623c9c29;
reg [MAX_SUM_WDTH_LONG-1:0]    I31ea69d26acd05d303178076eb123a7b2bbfeca82c2690c54323889753261f1d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia84ec437292f1ad3e702b4fa896a4f545cab7253574d294243af0c1e7de47155;
reg [MAX_SUM_WDTH_LONG-1:0]    I52cf6523f0dd5f666334b2646768fe4499c699c8f6b27ec32ae325cc0981a515;
reg [MAX_SUM_WDTH_LONG-1:0]    I7da5ecb7bb8a413a5c6c51f0aff1921be97bb5df5d56f6648c27ee4196fa93db;
reg [MAX_SUM_WDTH_LONG-1:0]    I81c612bc8b32254693a4a0c89fb21865b161dd1673f5610732b31dd5663f160a;
reg [MAX_SUM_WDTH_LONG-1:0]    I5b143cf694d99dabce0cb40d2d689fd7232531ab3a30888f811171b6aa2e024f;
reg [MAX_SUM_WDTH_LONG-1:0]    I050437a5474ba60337593b28d17e2bec5c76d26ea8afeac61be93e8ba0ada42a;
reg [MAX_SUM_WDTH_LONG-1:0]    I0442e99f7519b58fb576a898b41563a174beef69bb6a525712224f5d767a5867;
reg [MAX_SUM_WDTH_LONG-1:0]    I4bed271962970c26ab72de275bea4b2fb0565d7e44f15b2a1df631bba9e5d4e2;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaf95e616f53a061a7bf59bf1128d2cf6a5ef64d24b292671a3124a6e010d964c;
reg [MAX_SUM_WDTH_LONG-1:0]    I41b85a49eea9c0d773ecce66f0023338d3ee5a94e14a87c867a74960d30211cb;
reg [MAX_SUM_WDTH_LONG-1:0]    I3390b463514e772ff0afe74698bc4850014fbe363d105ce3d0e8810706977682;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e5c11a25b8726c787dd0ffc08e93b671baf84832d9413eb7031a6fc17e8ad76;
reg [MAX_SUM_WDTH_LONG-1:0]    I6b499c648458a2ed0cf0b27d81aeb706a260c5615a8def0ae89a1a44693061c5;
reg [MAX_SUM_WDTH_LONG-1:0]    Id3bae057e39f6549ce13910da61dbb41693ff87efebfd241bd1410d3da7195ef;
reg [MAX_SUM_WDTH_LONG-1:0]    Iecf240e8fe5f620bf43121455ba23a715b23f53e049d2a36f4bf52e2a061a8dc;
reg [MAX_SUM_WDTH_LONG-1:0]    I7958c747e1ef37e2995c52178d143af6a5f3acdf7c6d1cae518c82653ec18716;
reg [MAX_SUM_WDTH_LONG-1:0]    I697a55c4cb2dd56ce91465bb6750d05200607607d7eaa0b27accbf7f20ba97c4;
reg [MAX_SUM_WDTH_LONG-1:0]    I2785beda1166504e0b7ea979dbf6c2c5574159cfe36c60fced2dc64ebd05a9bb;
reg [MAX_SUM_WDTH_LONG-1:0]    I0b60295163435ae3d3b31e9613d753e7e41fd66c11fdf2e7248d7864e11d9d84;
reg [MAX_SUM_WDTH_LONG-1:0]    Iccacefad631e33ec8e54f8261759ca110fefaa6fd9fad08940205708a7180eb1;
reg [MAX_SUM_WDTH_LONG-1:0]    If07308cb71758beb15e4a33e3770aba8021bd5572128b9bbc1c8db48e7f807b4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic2bb8293812351030940ea0e0a882994714d60a4963e82e2291f6f2d386fce8e;
reg [MAX_SUM_WDTH_LONG-1:0]    I83ded8cd9258de3ae8deb907ae3b813cc228b189df92f42c55a4b0eaf411c106;
reg [MAX_SUM_WDTH_LONG-1:0]    I89ca3ef99e4b84441ed3cd9f386109125b6da2d23485fc22513b1d8ded87f894;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibf9f290605da4b6295c786c6ebc135cffc80a3352b42e1d841ba5f6fbbf06cc8;
reg [MAX_SUM_WDTH_LONG-1:0]    I0b2f8e7646b38057090faea20bf55e51f17d23baa4daf0c16d00e75e4c5f0ebb;
reg [MAX_SUM_WDTH_LONG-1:0]    Id2dbd07db2080c14fd0026396339e31183fb5bb6a476999102300cf81f34b93a;
reg [MAX_SUM_WDTH_LONG-1:0]    Iba5fd100311e883873db0c3474169654308059bc4c43d52479a4515fa85e8900;
reg [MAX_SUM_WDTH_LONG-1:0]    Ied8c84dd66ab8e8fdeb83c6156b8a6f8cbcbee27c41ccdd8c4d199f70ea67e8a;
reg [MAX_SUM_WDTH_LONG-1:0]    I1ae7d02f524c03ca060c3dbc879653486c099ecee485690ce40a355fc1ed843a;
reg [MAX_SUM_WDTH_LONG-1:0]    I43bd10e4f520ec08b30e8474404cf62a6ad869cdd1d280a2d221e0d76f228091;
reg [MAX_SUM_WDTH_LONG-1:0]    I7e12dde03af7a5ae0d05cdc9b29f31ef726c7bc51a7f07e374bfbc0846a24f0b;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e7725af7e163a3f4ee8bf63bcb825b6d62f4b9260a7c68d0beeabf35eea9391;
reg [MAX_SUM_WDTH_LONG-1:0]    I9a798d59823ac9a032d0daa203a7bb153e483bbe4fc47083c1d7e4a65e400156;
reg [MAX_SUM_WDTH_LONG-1:0]    I453d1e19585e0fb4fa66d684f0e6b37f56990cf101cc3942d5d4fc7e2313710a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibdfea3d72843376261dc3e06e3f19be4556508098d1b4d37c1c4cf6928860719;
reg [MAX_SUM_WDTH_LONG-1:0]    I39249b7f0d22c6116a7dfd0c0748123ebb6a9b7f931a492a534702157ab28c3c;
reg [MAX_SUM_WDTH_LONG-1:0]    I1ee3ce036ac0c878003d846cdc3fa9f6b5854855789ea575f0005a9c9937c58a;
reg [MAX_SUM_WDTH_LONG-1:0]    I91c40ee5121cd738ba7213df9bda6130b101385a28d8a5fef6544c86f6bd1e3d;
reg [MAX_SUM_WDTH_LONG-1:0]    I465489f86885351586de73a0aed556821e0ce34d1c2cebb67227004b4503eb3b;
reg [MAX_SUM_WDTH_LONG-1:0]    I37646f9ba79338e88c3d793a27911c88d573dc5c1cceaeaf565606c5b61495b6;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e95ffa3fdf70dc76c935f7d4dde6f39dfba8eb795f7ccc55510ab3caf678410;
reg [MAX_SUM_WDTH_LONG-1:0]    I592170f431e8a8e15769fe2e5f3bc43a7c514290149bf9b93a8f3d3a748094a3;
reg [MAX_SUM_WDTH_LONG-1:0]    I2fef37935343317384b1d29a04765327533fd87d4fe82a74f24b8196b3dffc92;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie57f94a45eba4db3826b22e3eb6acfcfa04b6d0669e22e5b78dfae4e7659b205;
reg [MAX_SUM_WDTH_LONG-1:0]    Id5eaf1d953b17df3896f9a30f37363d1a69fe3a956b97d307c895065ff32674e;
reg [MAX_SUM_WDTH_LONG-1:0]    Idcb8d71f1ea9d314ae8f26e9f4b9e25ed245bad319b9af2f71b035aca6d8fa6a;
reg [MAX_SUM_WDTH_LONG-1:0]    If307a1ee8e5164bac03971d07c03c3c0440857c7cc29df11a751b3bef9bb1516;
reg [MAX_SUM_WDTH_LONG-1:0]    I3efcac0fab0af81582237cdcd612c8d22eef1a6534816484190db28f3e7f3a96;
reg [MAX_SUM_WDTH_LONG-1:0]    I3f5dc950ac82420b73e1bc98c8c412f7e91958fbf455413c6a0ea5b2569e078f;
reg [MAX_SUM_WDTH_LONG-1:0]    I42ba6c66d951bbe03a57fa7a4926d6323f30784fe87de73cce065cccaa9814b1;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac102173e8323a836c8f86d266f551fc24ccd14aaf39c7d9ef26c465d38706ac;
reg [MAX_SUM_WDTH_LONG-1:0]    I2976810df2af0dd2879fac8afe975126944b2e40a51dc7dd169051bb5086b3de;
reg [MAX_SUM_WDTH_LONG-1:0]    I9c3d0fe7d767050217425eadb8e780e5eeeb31239f2f517ae5d122bee4157180;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia7d01a6ab6c0646f75030a0bd04a711a9c50dc4674c921680034012e67a0c3ea;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic8108e830a58b12b8e3ef4897cee70758d1539ae6609d73b5455b94b0eee5510;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic96ea379edce04b88c524fd17a2b6fb2283e45735640aa3d8ffc7f1bca77c78c;
reg [MAX_SUM_WDTH_LONG-1:0]    I4c871d8c6a677ef8fa6c955524def78e8df6f9f3fdafb141d43db76d4569104d;
reg [MAX_SUM_WDTH_LONG-1:0]    I6f7a9d597443df1a96370dbd5e1c1f9cb563fdc4db1d00fa66e8a287fca9bea1;
reg [MAX_SUM_WDTH_LONG-1:0]    I6ffb18ff0417e140b26d84cece8d23ea507516ebb60dbee4438e9433713c9f81;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia187792bad45afcf25df25b18a076d255536e94db8d7bac4df79761df5f16050;
reg [MAX_SUM_WDTH_LONG-1:0]    I9c0a341c77ecbc1b3c44afee03ccc5a8f34b1275db9c439eedca9ff61a1a1eac;
reg [MAX_SUM_WDTH_LONG-1:0]    Id8cd2e026867692af509cd433fda0fe6a8b5ccb8ed91bad6530d14172dbf7375;
reg [MAX_SUM_WDTH_LONG-1:0]    I2ad4afbffd2865f5c89feff965381fdaf73ac9ba4bc6e802a39014fe554b09ea;
reg [MAX_SUM_WDTH_LONG-1:0]    I31adf91b5f31b4232ee24f82af27e02a7ed1f8535c552409f353690340b64b2c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib96bae85b07ff95f5a6716cad97c765010937888a28ad63b16eef3b6ae93b3d2;
reg [MAX_SUM_WDTH_LONG-1:0]    I91cff501b877ec0153cf2d85abd12870d65d1aa997a6bea7d653bf387813998b;
reg [MAX_SUM_WDTH_LONG-1:0]    I42295332275fc6fcb94c042fbe6b48d3d03038fc27c535c7e63674f58da60bf0;
reg [MAX_SUM_WDTH_LONG-1:0]    I445cf6fbf071cc76e6fc981d7f2f201d0e09d3f47c1227feaac47fb57a14e85d;
reg [MAX_SUM_WDTH_LONG-1:0]    I96ace764b2f8db5049595445104a408a641999152f2a6c63d22bc6946c27322b;
reg [MAX_SUM_WDTH_LONG-1:0]    I8741cd8af2f9c3a548c5c39709d7a186f0953de5af6d09d88901e0083a539096;
reg [MAX_SUM_WDTH_LONG-1:0]    I97a73864c1c919943cec586befbb524fa6d6da6a60e1503bcef8116c646b71a0;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e4ad715cc833c775ed97e88f28c4196d28bcee4370205307f4266e1fc572cb1;
reg [MAX_SUM_WDTH_LONG-1:0]    Id1fb56c160d418b26fe2b51dbe78addbbd2743e7a342e0b6bebd2e8d3cb1ce99;
reg [MAX_SUM_WDTH_LONG-1:0]    I20a501f960ccd425135a3fcb8e667d68940a5950d939bca37d107d479984c038;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie28b77da5cb0eae41811ec7dbc5f86111d64b794121eda9f2f0515324579f844;
reg [MAX_SUM_WDTH_LONG-1:0]    Iefca48dd9d0f3c717b0a3b081894e93ac451ed275f3cfa7aed675f58327a2d02;
reg [MAX_SUM_WDTH_LONG-1:0]    If6592aef798f1b26c5c6593d99137d00bab8e8631070e89dbc6a3e11c89b3e92;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie14918150ed723163714038f6ffd2c64b07d62079dc03ac8fdeacde45633def9;
reg [MAX_SUM_WDTH_LONG-1:0]    I5a03d267642091bb2d177a6689d91b995983fde126d703c6474d730b455ab56e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib6dfa3959980c5d348630e2edd81fdee8429a3003b0a21369b99343bda03e2a0;
reg [MAX_SUM_WDTH_LONG-1:0]    I97f8487b89684c5c6952770b0468738f72682d6230be6a5a31a92fe50bfb239d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibca42a442c971d363e4f848d203d2782af05ddbaad93e8cbf334328d94a8a499;
reg [MAX_SUM_WDTH_LONG-1:0]    I84744085fa951f13f4fef6c44fb0180e543fa6793e89f4dcb14c3da6b27105b0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibc54f1c4736e5a4608208441ce8d81831a0b6c7448083d6e6976981f8a38d1c9;
reg [MAX_SUM_WDTH_LONG-1:0]    I211a150dd66153a3c2c72be4c24145e4c9f0b2f9a3032fee9233985ca9d2c4ae;
reg [MAX_SUM_WDTH_LONG-1:0]    Id9a38b1906060dc5739f9446bb2dd1a6b6603924d4b7889c931988fb52cfafff;
reg [MAX_SUM_WDTH_LONG-1:0]    I8beede7aeefea570e5c65a76dbc5ce1f4eb114e444ea9b4636258bcefd9d5f34;
reg [MAX_SUM_WDTH_LONG-1:0]    Iabd5561747d288862c0b289a28572fb5b0159a3fff7f79c59bf60f1612ec1e3f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia4205a1d01cb014ebf8e1d539dbe1c7270bf9bfa8eb7920b136417bdfb9f498e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic45f0213074aad63c68cf3fe879ad5b0e70a5977f282822ab582ab88ae7236bb;
reg [MAX_SUM_WDTH_LONG-1:0]    I123d4c26243478ad4cff3406be39503c6b378cdefa50bf60249ec03d3a44270f;
reg [MAX_SUM_WDTH_LONG-1:0]    I0f75d5771cfa314d28e188de297b4bb53c2cb732724a630e10580ee5fe87cb23;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib6f695414c34a124de17de5cee8798a33f0968f7eca5143f21f88c228ffa6345;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib43a705a217dd9f2321c3e61ee116d257d8ad59bff5b4f80435f9dd96a8d04fb;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e014fe75658214d8ffa60f966549b131bff6a16020d7858523ac829b0126838;
reg [MAX_SUM_WDTH_LONG-1:0]    I31734ccacbfeb8a5c0c30cfc84934f8d1636ce4ecae14fe7809d6aa8df35a9e8;
reg [MAX_SUM_WDTH_LONG-1:0]    I701aa61e04d2787a36f529185ddcc94c832834d38ff92b37456b64ce46c69b2e;
reg [MAX_SUM_WDTH_LONG-1:0]    I4b9dd5299690e88d870ceb4939b7f8fdffc8419431458851a3691de4f78f9f15;
reg [MAX_SUM_WDTH_LONG-1:0]    I81b8212f2e15845be4d129b192895f659d31a061a3a033bc3ac9ebecc75f73fe;
reg [MAX_SUM_WDTH_LONG-1:0]    I1f070cf569961de917cbd287e7b14a2ad6e04a4474edfb92c095f6e9cea1efdc;
reg [MAX_SUM_WDTH_LONG-1:0]    Iae16b002804d17ac9e2c9655dda031f3f0ac10d703bc42079ee2a5fd3ede604f;
reg [MAX_SUM_WDTH_LONG-1:0]    I5aff0a6c62deaff6e9d15280ae8c3cc326ae7f9ea6959dfa41a92c770b592cce;
reg [MAX_SUM_WDTH_LONG-1:0]    If6fe8b42d897a8c92c628edac7869deee179622fa52fa779f2d9a0279791afc0;
reg [MAX_SUM_WDTH_LONG-1:0]    I10a223d797492c10ad8f6aac1cbdae83833e701ae6314ed988ac117debc98c33;
reg [MAX_SUM_WDTH_LONG-1:0]    I8cf1c2115398eb404050fcfc654b198694d3c54eaa592d0d725b15e7937d8cd5;
reg [MAX_SUM_WDTH_LONG-1:0]    I6ec1c8ffb963fef21e978fcfd0268bc24dd283819081437974fa5a06caa64c25;
reg [MAX_SUM_WDTH_LONG-1:0]    I781bae0d109036c417f71e00a3df3440df3cecd691fe1f67c147c4d2de217f7e;
reg [MAX_SUM_WDTH_LONG-1:0]    I10ecf0f58ee2fd15e2b4135dc03cb4053c364660c6d2e2bd03cfc37aa6d6621d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibe646b6da0465c3fb411afc4e03d45f553cf91e67cbcd46674a0051ac1092e30;
reg [MAX_SUM_WDTH_LONG-1:0]    I8a61ed94b6198131fccf4feb6be7327f59408e9de4def9c4a155167192c5f065;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia57f6e4dd9ce4389f90c78df4fca73a681df346f58a85f61a74e842427848347;
reg [MAX_SUM_WDTH_LONG-1:0]    I3d284d86f6c46162d3e0f913a5a6b0e1f2e34fc7ced6a0c226d5e78da81a0633;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib07af5e0c881985b1aa0698382702f78d3ec7ac69cd0deae7496bc63e519a738;
reg [MAX_SUM_WDTH_LONG-1:0]    I332737561309225f302f64e49e8b3e4aa4dc35344858059b21e146e8cb84a466;
reg [MAX_SUM_WDTH_LONG-1:0]    I7e3620302652666ddabcd16531a36e7af51722c39bffc4224f256a34ca33109c;
reg [MAX_SUM_WDTH_LONG-1:0]    I6c8cd97a5a950e00f0b9892a96d99ad1e5bae6c2db215bbb532060b753233aff;
reg [MAX_SUM_WDTH_LONG-1:0]    Ice95c4df972e8e6a31901269a2d291a70fe4e8dd1d86ea5ded5a16cb1c169890;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibdb4937356d2b1cd2091a695635cc7c69b694f775f4c4e8680ea49df1ea6722d;
reg [MAX_SUM_WDTH_LONG-1:0]    I95e467521db517b858e59156f95992ddc522a7d038ac6bbe691a91b567cd35af;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia9160306dcccf07d591c6c85cf86175408905d5e1bdfb36206d9c4bb5b917dc4;
reg [MAX_SUM_WDTH_LONG-1:0]    I207af234897ed272d784f4a9f8850eaaa2fbf47f583ed1f0564201e33dccfb66;
reg [MAX_SUM_WDTH_LONG-1:0]    I0738f605ff9ccae9ae63f8e6fe7a9b537d97e13bf3f23c7b0daa4fc414eb7eb4;
reg [MAX_SUM_WDTH_LONG-1:0]    I7c10e2245efc27a4e2a96467eb4e3fd9c28be5f26f65c560653ff4742fa5143a;
reg [MAX_SUM_WDTH_LONG-1:0]    I00e08c73bb2036cde2d53598b9977dd2504934b9ba8b58bfccdd21adc2fd223f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia718f1fe0157bb564650d817f5ea7960bd0698409dd04d9b31d54c95a3f90318;
reg [MAX_SUM_WDTH_LONG-1:0]    I95b908a4845eb4b14e8f933057bab27e44c6a867e4bb02d87417740e3150e018;
reg [MAX_SUM_WDTH_LONG-1:0]    I600d6bfc6bdecb80f4f9d6020bdba9b4c04bcb359e66e793a3bd6732173d0b17;
reg [MAX_SUM_WDTH_LONG-1:0]    Icc13ce9fe63ee1c11fd5dddbf0a294cf6ab7ae703f742a92150b7a77868a5a16;
reg [MAX_SUM_WDTH_LONG-1:0]    I2fbaaffcceb2dc6a4f6d9d34140997b18356dc3803bb0a6c6d5f1b3f980e18da;
reg [MAX_SUM_WDTH_LONG-1:0]    I3c91639fa462a2a7e65410080b46408b692ca4639ed17637b1d465f38631734d;
reg [MAX_SUM_WDTH_LONG-1:0]    I3adad3708bb709ccb06c77ab54c92b6c6629853f740147fd958e6200aeee81bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I706a44814e015449aad217d9bd9e0056813b075d8e622aaec4dc08a3518cc0e5;
reg [MAX_SUM_WDTH_LONG-1:0]    I18e5d7f94022748f9a5645c2b0e385407e0f00d6f9ab28a55982fd36330ce524;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0090ea9b75c69dfca34ac43abee88b20734f7afb9c1d88f95eda3df6aab27db;
reg [MAX_SUM_WDTH_LONG-1:0]    I062483fac022c2d74cc4bb84d57c636a3bbb67d68dacf0da453e3b5f71ff8846;
reg [MAX_SUM_WDTH_LONG-1:0]    I15ba9fcccc2e3aaba7bb5967d35eeecfc3bfa7ce27f82435be6dee9d0a4af829;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic1034fe189ea09f2aa3b69428828a2b7dbfe9389dcf48dbdbe0f15b9157f7c49;
reg [MAX_SUM_WDTH_LONG-1:0]    I8a3c94278b7c901702cf1b70e89c1832afee395077555d27badd4e2b6fde0b7a;
reg [MAX_SUM_WDTH_LONG-1:0]    I23d075a3ac353b3deca0a572e9cbec9b1ae24ffc7f134b36c6f938d949bdcb1e;
reg [MAX_SUM_WDTH_LONG-1:0]    I3599299f7f89ed3c6b11b31caa26e6b30553b9dcc1d5968283085959f822a4c6;
reg [MAX_SUM_WDTH_LONG-1:0]    I8954b3335e6848eaec70a960b632233aff75de56bd0bb895e2b4ae49095fe19b;
reg [MAX_SUM_WDTH_LONG-1:0]    Icb88d7eda8505d92744b075a1c229e3c0f6a9ff062bf5cd35f6f84467b451e9c;
reg [MAX_SUM_WDTH_LONG-1:0]    I20ac47b3e52f25ce7858fb7952654107faed4cb5cf3abe1ba915710d1af4c933;
reg [MAX_SUM_WDTH_LONG-1:0]    I53a66c670d7345059cea712c026fe8c524e74b030af0de054cf6e053bb304248;
reg [MAX_SUM_WDTH_LONG-1:0]    I034d52d03f918c91bfc6236c72b0d40b688e2bd353f9ca1f03f4c61449bf128d;
reg [MAX_SUM_WDTH_LONG-1:0]    I727007bc323c90e0c264e5b8688898c0df1bb72c976fbc3513439c14f15b5733;
reg [MAX_SUM_WDTH_LONG-1:0]    I0011eafd50b7df59be2a4f143443c0ca8ea87f9a93586d07292ba02fdc2b9b4e;
reg [MAX_SUM_WDTH_LONG-1:0]    I7f3447e248449854eb030c79bc32b602d376441a193e25bfcf9b8a0eda83b57a;
reg [MAX_SUM_WDTH_LONG-1:0]    I288ddea916663f74bb339e7a94ac9c86412f39671ca69dc7ec1da05a1800092b;
reg [MAX_SUM_WDTH_LONG-1:0]    If023ae056e9b4b370bc83a2d5604602f45a01a005bc19a769c874536faf4abbb;
reg [MAX_SUM_WDTH_LONG-1:0]    I48ffe541268d63545fa48263d8df3c288af7b2646b4dca546a4dc521aa247651;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia81ab6d41925460c11303075dea72c7fb3fe533d88450c32414823fc5b10bfaa;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia7a158b91a24000cb6211d129d65e781a4e28b8333f897bb401042fbe17c37a1;
reg [MAX_SUM_WDTH_LONG-1:0]    I698aa30e42ad4f250363d29dfc5117677b19f2da0afa75a013718ac5b9731d6e;
reg [MAX_SUM_WDTH_LONG-1:0]    I144fae9c9898630fa027b3237ed3434c76965eef2eb015effa7c8677b19c91a3;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic595c984782ebc89b61fa2a64e994aa66eb4979ab1e30e890886355dc247a67f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ife11a6b34a661bffcf9f0147459d2f5a23d6c5460c59142668ee0f0506755225;
reg [MAX_SUM_WDTH_LONG-1:0]    Id73bbd3c91f1e5fe13f11e8849f77aad2ddaa35d1399140ceb5e133da8e11227;
reg [MAX_SUM_WDTH_LONG-1:0]    I2d89506b7ec0311db709c4aba53b749ec1b531bf4bc7867f3866c39a73aada38;
reg [MAX_SUM_WDTH_LONG-1:0]    I390750ab5fb20d9be34ce0e294c95ca61ab6e511578b636301037a34f9bd9c07;
reg [MAX_SUM_WDTH_LONG-1:0]    Ief01c27ce040b3f50c19615a8f5d9bc8b467c0f88a778888fe186887b19fd580;
reg [MAX_SUM_WDTH_LONG-1:0]    Icd850fa1e932d19313713c2d376413e7b81faea883442278fbc700a2238f6779;
reg [MAX_SUM_WDTH_LONG-1:0]    I5fa215eca11a15c7ad85760cc87a0f8e883d02472c7af460b13cbe214a596c62;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic336cf50b44edc74db080d1127ba09a4313c0972702200ac5207aae8ce6b1062;
reg [MAX_SUM_WDTH_LONG-1:0]    I19b5f6ad3c2f2551b49883fbab077c8e3d76392fa42a5030b1f832917bc2641b;
reg [MAX_SUM_WDTH_LONG-1:0]    Iee901b35683b34719c33d63d90b8ae11fbc338a170164aac943fb0b495c92b97;
reg [MAX_SUM_WDTH_LONG-1:0]    I4d316d60bd6537dcf09dd9b7eecd93c86af11ddecc1ee65e4b9d65c136527e0d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ica10d27b8c94c1e740a2287ef28e5d3fedab4221b391b0a3a1da3a472f094039;
reg [MAX_SUM_WDTH_LONG-1:0]    Iac3e25273f8b972112775f3aa57274eabadbc2da5eea147328f85a941b959bfd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifc38f7d8250994e5e62716048122eabe81722a32478caab729cfb06aacfc09c2;
reg [MAX_SUM_WDTH_LONG-1:0]    I47b18bf83ed7f7e8a2c69814aafa41a66b6838a5a997d036c634f488f1c584f1;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia9f80db3bd889aa11f43f6aa371715d6aadc7d3aeac0e9519f79b787da6e545c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic4c53101c741f07c928018af5696d83f45a29d0e5a9f766bd2f1f1404f3eb59e;
reg [MAX_SUM_WDTH_LONG-1:0]    I4b15e4ecd6a6f2139463d94eb4061a410569136410e469abc38dbf8cc03948a2;
reg [MAX_SUM_WDTH_LONG-1:0]    If377629f88304a78a44bdac612907792b54c49caf9dbaf85b3061be5baa2f5e6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibb72bc519d54383d213250311085f6368ead1c943881ccc23f944e652f934063;
reg [MAX_SUM_WDTH_LONG-1:0]    I91e90d84eae561663a2e9e59f79782a78095807b98187add5501500b8c1cb126;
reg [MAX_SUM_WDTH_LONG-1:0]    I7af411084739689195bff036e9d5e9a950a7691f7d771d4d406aba4c32d95116;
reg [MAX_SUM_WDTH_LONG-1:0]    I06414f803df7c8e59f01524020e09627cb11f3809c3456a9a64655062b110885;
reg [MAX_SUM_WDTH_LONG-1:0]    I4eb359966514f007fea3e135207ab27fc596987f985b8a3ec6bf51dde2ff9e38;
reg [MAX_SUM_WDTH_LONG-1:0]    I60f3a2c7d8e3935c04abc8aa09b0a2ef540f13bc98beefc600fd70aa25421191;
reg [MAX_SUM_WDTH_LONG-1:0]    I698accb14122caa36f489e7fc522e39188ee03651ef0c6670eecd60162cf2f0d;
reg [MAX_SUM_WDTH_LONG-1:0]    I49a96e94f51c41ba36bb7a8d466771682602e2dbd6f65e13d7e858a60b554f3b;
reg [MAX_SUM_WDTH_LONG-1:0]    I79d13cc47977ecb1fb0ca304be8c225a427063b4328cea4c4a227521a1f26018;
reg [MAX_SUM_WDTH_LONG-1:0]    Idcc1ce57eae666070b5b9984cf69d5d2409ea92b36718906218185325b5611b2;
reg [MAX_SUM_WDTH_LONG-1:0]    I54feba5563ca84d4a04e3ff7ff5ecf689d26961daf0ce27f0be8988087296fc6;
reg [MAX_SUM_WDTH_LONG-1:0]    Id60b48bbf346bf95a242f425de7f456aaba5b3ed35cf16a07ac541ca8f480319;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e89f3937a947ff09fef0df8085edc1dc09a36d7bbb39027d358384d54088060;
reg [MAX_SUM_WDTH_LONG-1:0]    I800a86b8eeb247f39df85aba37dbaa93060858c235c6ac6b0912fca85af95477;
reg [MAX_SUM_WDTH_LONG-1:0]    If4b0b6bcc29aecf6816eab93edb0cb358730913253ae72d15db63ae06b19c52a;
reg [MAX_SUM_WDTH_LONG-1:0]    I63132df742cc353a39f27a7a5a00e0990e9e9e023f5c2a8bd571fcd6dd2d760a;
reg [MAX_SUM_WDTH_LONG-1:0]    I0734166e34887037bf713bdf1df0f7219241551cec455ed45881734727f90032;
reg [MAX_SUM_WDTH_LONG-1:0]    I9f08c1a4053ac65909c96d240c83e15017c81fa41f351b0a707fb7882e49f4c7;
reg [MAX_SUM_WDTH_LONG-1:0]    I3af491b2352720f2bd378052706f4ce571453d59b0fc78b3cb0bce2d51ce5700;
reg [MAX_SUM_WDTH_LONG-1:0]    Idb883f1d90a389f89c3e04f54dac20f205951bba3fd0a00e9432498c4def1131;
reg [MAX_SUM_WDTH_LONG-1:0]    I4e556f27c558f3d1f76d2ed4a3f0b1a68d74e5c0ce6370b9eec599e7f76f8bbf;
reg [MAX_SUM_WDTH_LONG-1:0]    I02962ee90b42f9b95262049bd2dcb7da2f43333787a578d5f5721681773db287;
reg [MAX_SUM_WDTH_LONG-1:0]    I739fb2ce1dc1a27f40af1c53d575108539718f9d60f83de60531d7bb201685ff;
reg [MAX_SUM_WDTH_LONG-1:0]    I1a6ae2cf67f356fae1ec533488e09c6696277823378b06751db7ec97115d9c00;
reg [MAX_SUM_WDTH_LONG-1:0]    I931537d878467c473ac81aec8f9a7d79f286024e62ada1e5f363b93d6887070a;
reg [MAX_SUM_WDTH_LONG-1:0]    I61e7244c25e176443b24d592ff4299482d572c1705c3e0a6b44698b5366ea3ff;
reg [MAX_SUM_WDTH_LONG-1:0]    I3b3f53fca961a376010d1a5b0c49f91d58b351d0306b8433ac22a70f5a1f1673;
reg [MAX_SUM_WDTH_LONG-1:0]    Ica809c2eeaf6926552d9f811bf16c30146853674185c2315876fb5b2ea6d0769;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie3e85438dc476813cea40910227c7d63eb275948fbd481f56cc51656c1bc8b34;
reg [MAX_SUM_WDTH_LONG-1:0]    I877734e2edefa267510037759c9490dae213d2e046beccfe87e16c1aeb5583c4;
reg [MAX_SUM_WDTH_LONG-1:0]    I8b5d8146640c84b84d0d6bcb2362fd5bc7e7462e1905b32b998b1f00f2da3645;
reg [MAX_SUM_WDTH_LONG-1:0]    I57ae0fac4bc1fada55e48ef9952dd7b81a55414196fc22fb27a20b723832aa84;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia2343365eee39c9305def2bd744d3e44bf20b5bab8a48c6a2d95908f74f3cd18;
reg [MAX_SUM_WDTH_LONG-1:0]    Iadaa0bd11c77d7ea8c8cfc4b0c805c5afe6b75f597b03729ef2cb704dfe48286;
reg [MAX_SUM_WDTH_LONG-1:0]    I0543957798ccd8923b2a5b736175c6888eb71c1466a1e9cc7d7635701e103823;
reg [MAX_SUM_WDTH_LONG-1:0]    I87c64e9e81da569414617b07e39a7f67b0b76c71643cf7257b7374feb6fc9750;
reg [MAX_SUM_WDTH_LONG-1:0]    I481cb000cdc7a32db6aa5a6b0da57b76f53f5bec6ef93d4ee25557e1b12064f8;
reg [MAX_SUM_WDTH_LONG-1:0]    I23f5e95dbae4b1223d603061df9b75b9a9ae8409c6bc4ad1fe23d3f5c7a68bb1;
reg [MAX_SUM_WDTH_LONG-1:0]    I16778a093510ae433495baf9d2b7a74ad4c5315403d0e8aa39eb09cf508dc201;
reg [MAX_SUM_WDTH_LONG-1:0]    If2cfdc638b3cfc13d31615533cea59a4bf8123299239956479d3f1d702ef54d7;
reg [MAX_SUM_WDTH_LONG-1:0]    I114dd7172ac111bca494cc4230447a2dc167f12f198288d34cb5311c279a73b8;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie72b5524b212840dd1e69f4fa41b4955ca028c1ea7fd2f3440843cc2ef6d4be2;
reg [MAX_SUM_WDTH_LONG-1:0]    I8b151ef6b3125cf983140726d775d948a253c13f020d3d1e75b585afb979bc8a;
reg [MAX_SUM_WDTH_LONG-1:0]    I72329ad9fd98258074b92a7e88a88c68f8db57e7d6460e9c29ec7f3cc251de29;
reg [MAX_SUM_WDTH_LONG-1:0]    Icdad18f8878b4e9645b4f2d2434f913a6e0f732a20a6a750e25c2398a086ac2d;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaf14e804e3bb7cda8e67e39af906be2c966fbab4a6e73b8d60ee7ac5733669e4;
reg [MAX_SUM_WDTH_LONG-1:0]    I238b01744b520f8759a7e466290a15b15b96fc95b4b8a14afacbedb1657f7069;
reg [MAX_SUM_WDTH_LONG-1:0]    Id29a54af13b6045a8a43f741c229ff88d4aeeffef29065cb29cffbd861479f7d;
reg [MAX_SUM_WDTH_LONG-1:0]    I9ccd1f3aa9f849bfe7dd9ff5f9de6fff64a444bc5286321a1f0e73e990d6a996;
reg [MAX_SUM_WDTH_LONG-1:0]    I02ff320cae73fe5cc67804e552bffba75496861f085869eabab140094a18fe90;
reg [MAX_SUM_WDTH_LONG-1:0]    I6eba99f7e39a1779ace2db8cd1806d099e7cf0678ec385baba570209f784b5eb;
reg [MAX_SUM_WDTH_LONG-1:0]    Id4182b8f05992677e12502bcc058d967481d0dc2c9c4731b657f04696a5b5bbb;
reg [MAX_SUM_WDTH_LONG-1:0]    If4927b8f31777ef2940c413336113e906e0e3556c31b9b3233107b88b1d71999;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibf57f9e63049a49e05739966f1ec2fe4520b2959db6fee3a18ead9ca03aac230;
reg [MAX_SUM_WDTH_LONG-1:0]    If0025a7dfd37802d1a1fb43d82ff871c2867504735093f0ffaa8b0d85fcd4d1e;
reg [MAX_SUM_WDTH_LONG-1:0]    I24dbfd322139e6a1964e587f89b06274c35617e961a5f61f90c67ee3b20ff208;
reg [MAX_SUM_WDTH_LONG-1:0]    I8bddc257a28da31b71dac60701bade264fbf14f8377b1f504ef874c72e0d45a1;
reg [MAX_SUM_WDTH_LONG-1:0]    I225da3a8a67ccba14e13c78ca2ffd83b37ac9a961371f1aa617f5752b1bb337e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib9855ec95d5c99f93ad4c5565e622dc1c2d1c4a3b5d0937219172d97ac290756;
reg [MAX_SUM_WDTH_LONG-1:0]    I598f53ba5c7ffa41f21af94375843b0b7a911670719edc80705508ae32ac0ddc;
reg [MAX_SUM_WDTH_LONG-1:0]    I18eefcf5075eee79120ffa0e5875cbe7632d1db84b1c498107413f14b72820f1;
reg [MAX_SUM_WDTH_LONG-1:0]    I7cd31013bf73ff7f7aafbf06eba3fe8110dc5490a280c2d79ce53c77896f564f;
reg [MAX_SUM_WDTH_LONG-1:0]    I804112f16593c6ce81f6459599203b07642485939c898d78e113353659a62a68;
reg [MAX_SUM_WDTH_LONG-1:0]    Id8a5ef9ce42d57c3feb442ca091604f1fc51e648a89794ea3fbe4b30537fd286;
reg [MAX_SUM_WDTH_LONG-1:0]    I6ec3df474c20bfab5d99aca971523dec8454a5ad4536765f4f9bcb0c31978cd4;
reg [MAX_SUM_WDTH_LONG-1:0]    I862b7b7769e1ce1579c40d6363e23230c9253630d97fe8abe72b80e8a8b5440e;
reg [MAX_SUM_WDTH_LONG-1:0]    I1ca12951f309a25752defa88fa366a90a13ce83b7fb40610c01a8c11a3c2e59d;
reg [MAX_SUM_WDTH_LONG-1:0]    I786cf639910ac9a90b1abf55f9e3b66d87c4bb98a2c8e38142969ee5aefcf6d4;
reg [MAX_SUM_WDTH_LONG-1:0]    Id059fc689baea934a9f278b1066a92d6aff850608c0797dd7257693cbfa40102;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic6d228f83da7a1c9a71d8fe70d5adbbab8856e5fd3640d805c4076f5f7d53553;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia61e8ceb90369d4ed8ed86b9cdf7d4e89056cf4fca5c7e223bdd7b2c5656ac9d;
reg [MAX_SUM_WDTH_LONG-1:0]    I30a86fd347fff855a807034e13d6e751b35d4330df8436470af7bb42af947668;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic3d44900d87d02e6912d962514abecacc6e1f20fb71c052d58a896c5524e1703;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibdb62dc1ed705231a9d0a9e819d824f81e62746fd6d9877557622a8293c7cc3e;
reg [MAX_SUM_WDTH_LONG-1:0]    I1fd78c97c2a03a51b8d2a3dce2a553514aaeffdc051bfd3820d409da4b8189a0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide94701dd8ad54a630c6eadc44221ee5786180f247fcaec8a7787f25c4070968;
reg [MAX_SUM_WDTH_LONG-1:0]    I4c5882b979d1f315e20e4a8fc06c794c0217b97de2613e193cb7a213c2119c97;
reg [MAX_SUM_WDTH_LONG-1:0]    I5b480e9176a1bb70ebc65f73af78889d266a8efa7414cb97cc5255a5ca5f01ec;
reg [MAX_SUM_WDTH_LONG-1:0]    I35ddc6b67ba559d53bf4b297c2cfd82bcc814a88095ccdf7d6f22fb59113ae98;
reg [MAX_SUM_WDTH_LONG-1:0]    I9fc15e538a85dde7207e48d484f796d96ac712463c802b6995b216e71fb74d93;
reg [MAX_SUM_WDTH_LONG-1:0]    I8029c5b828acc50a3a785cab42ada7d51c82647934a9dac7f4a738920f1a332c;
reg [MAX_SUM_WDTH_LONG-1:0]    I1d5563063ac8386b450a3a36bb3d0a3586cfd6d11471071685e3f7f897d8eff2;
reg [MAX_SUM_WDTH_LONG-1:0]    I99c4a78ad7af699907cae52326915f18ac1a2a6f9d99b2aa71c34d10fa78fbce;
reg [MAX_SUM_WDTH_LONG-1:0]    I1de9fe186e9fdadc6c62a9c6645dccfd3709778f3243d2a4155bdfa20d27a544;
reg [MAX_SUM_WDTH_LONG-1:0]    I4b18b20124a63f85e812047188401b685693ae009c87ae337b840a7a3e03f140;
reg [MAX_SUM_WDTH_LONG-1:0]    I73c8c2e52e23d992ea9758a361fb9550f0ac7f08bb93b6b26c6fab3b234720a6;
reg [MAX_SUM_WDTH_LONG-1:0]    I289b4317d3472843dd49dc75a39395f8c39b9fc0c70000205510d08404d824a3;
reg [MAX_SUM_WDTH_LONG-1:0]    I95b68240d25deb08902e18ba5fc3ed7af68c0a6ae8e629edcf59930ed55c22ce;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie6ccfd08b7627ae7cdfd608c7054781099d7df5a0f133672db189134161f76bb;
reg [MAX_SUM_WDTH_LONG-1:0]    I96ba46d5aa5ea6b2cc6a43df70554584d43f49a6bb171722373d28a2b0f1caa8;
reg [MAX_SUM_WDTH_LONG-1:0]    I1a54a485e54cb6d528feed952641c7e5350f3d386ceb62ddd2778ad179aef345;
reg [MAX_SUM_WDTH_LONG-1:0]    I072f20811fc3b3515b7794a416e5ba39cca6a9579de36442fb39771729dffa8a;
reg [MAX_SUM_WDTH_LONG-1:0]    I7f1329fd762cf679c07aced91992aea071fe128bc24f06ce88bf49e876578a9c;
reg [MAX_SUM_WDTH_LONG-1:0]    I26c556de81da143a85c36f6ba98648e110114ab97302046b7aec581a62689a3d;
reg [MAX_SUM_WDTH_LONG-1:0]    Iedb10f981e08498950a50589d8c2fd5dbff191f233da39d5819ddf2dc5172651;
reg [MAX_SUM_WDTH_LONG-1:0]    I2e063205340c315025edf32a4ba91e5f7cd39f37fc5800906a3862780cdf7d9a;
reg [MAX_SUM_WDTH_LONG-1:0]    I7bbabd42e7ee42c653f61b4bbd72ed2b076dec2c89baaec2b4589bd55b92fa6a;
reg [MAX_SUM_WDTH_LONG-1:0]    I90a0e50a5730714abafa98a7ad70e64903062bfe6f8deeb528bdd7008958bd11;
reg [MAX_SUM_WDTH_LONG-1:0]    Iff82ae02f527d0eff3c9f8bb9d8fc818cf9bb7e3fac1a127849eea6ba27a62d6;
reg [MAX_SUM_WDTH_LONG-1:0]    I4df045f8dab91c2eee20a03bcbea586a003659b77d8a6e941bd2b2ead3006d04;
reg [MAX_SUM_WDTH_LONG-1:0]    I9e8877d4beab63d4bf103c07e1cd9330daccde2cdd266b2942f56b2a8e8a926c;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaf763109fb82e88c7ec019f7b9b668f88f84a5d4f760592d2dc9172c75be0aab;
reg [MAX_SUM_WDTH_LONG-1:0]    I5059641c5d09a0369f6237643b75899865bff068e9aa8779d0befdbd53a6b754;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic24e91afb654a0ee04d27daccc66b42d5e001a5962acd08aa73c3e962e1f2c88;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide8930fe855e6fb7dd5b689395a121a16f491421d448454c9c021f62753732c0;
reg [MAX_SUM_WDTH_LONG-1:0]    I4909110fd7213171cbddcd3545ba2a0d3a135e723189edadc7c64599fd2f1f53;
reg [MAX_SUM_WDTH_LONG-1:0]    Iea55b5544c098ecff239cee665c2642cce17d3b546df6ea3d0c832a118c535bd;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide09a550a1cc61dd543f2dd7a6e38af908474f7c815ab70318871dece429d0bd;
reg [MAX_SUM_WDTH_LONG-1:0]    I1edf83d193e0825c58f470cb0d4ccd85e3df4652ab68fe3a701a6ee0e8a0658a;
reg [MAX_SUM_WDTH_LONG-1:0]    I3f3cf1014fe01e02bb46b2e8a19716cfaecfec0e44fcc344107589dc409044b1;
reg [MAX_SUM_WDTH_LONG-1:0]    I3724769b2a595469f910cfcf1f002009d9fc27808df7e59ce728af9a923726d5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibfb48072643b2cdc460b7a667940129aa243be78b6d57abbd483d5551fa36eba;
reg [MAX_SUM_WDTH_LONG-1:0]    I6efd033a5e005d772ae427cab43bfeacb72354d6905822aaf8d484125615d0f5;
reg [MAX_SUM_WDTH_LONG-1:0]    I44445d003eed631dd6933d4ade176469fe9a4ef0b21b0ee20067b5aae73704d8;
reg [MAX_SUM_WDTH_LONG-1:0]    I8be8cfdcda8c42fc83b767d9cdd6af256d434d307b8e324bd533b5b016383bfc;
reg [MAX_SUM_WDTH_LONG-1:0]    I31ef992f17daed0e1947c4d26611e7377d8b3049bb8ae2ffb3d56f3db5f85916;
reg [MAX_SUM_WDTH_LONG-1:0]    I6483bb2ee2f7c35aa35adc7fcb6cf8cd426e048f4aff95cb9f4f732f97adaabb;
reg [MAX_SUM_WDTH_LONG-1:0]    If550dcd8751a8725d597ff3b723c6b5cff949b2e3087c71d36782ea291f7bd3e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia810fbec78dcd5215c217347900257a8f892a4805dc2365ea79eaff74af7e64b;
reg [MAX_SUM_WDTH_LONG-1:0]    I5e14fc93aa39853d74e7844854278275828d0f5428f2af96c00c8b0ab141c868;
reg [MAX_SUM_WDTH_LONG-1:0]    I8a5d6a4832abe68ab6e9ae33b1b6026805c5db0d186df37fe623a2d9931b2534;
reg [MAX_SUM_WDTH_LONG-1:0]    I00c96393d166280a0d866d1999d4306a650507c7bc407202924f6684f61e219e;
reg [MAX_SUM_WDTH_LONG-1:0]    I2cd11587dc2659cd92fb2c4f894bbd9d252affb93f75c3c691dbb02225b4e887;
reg [MAX_SUM_WDTH_LONG-1:0]    I6aaddd1a59b6e96dd8cdd4a57d8fc03132dde1c5b0bd06dd6f0a240c2a04f947;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibee0b890887202cb33c8fb07639c7bc536951ce8e661d561d7e7a7355db5f9e1;
reg [MAX_SUM_WDTH_LONG-1:0]    I0a22f1dc32c83db6603459232e78078eac21f865aabe0b9a03923e63cea874ff;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5e2defed9b5fe67a6a551e253cf68006aca5e13092f7e9b53f8186c76a156dc;
reg [MAX_SUM_WDTH_LONG-1:0]    I102751a9d577151cf6f780ced3299363623ab308737d8483ccbe02118244d2bf;
reg [MAX_SUM_WDTH_LONG-1:0]    I5c29250eb53f0eefc2332419b6c8e82f97741659657c08af97f8443954a5385f;
reg [MAX_SUM_WDTH_LONG-1:0]    I4a55baee8cbea583890824bd3ab4c4391b9d44203332575c030077c6e0e9f862;
reg [MAX_SUM_WDTH_LONG-1:0]    Iaae1f131bd6bb3b2fd8e363e97f6f9e680c7ed035a086cdf2bef5cb7e023c6d5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic1711dd767cbb72abed2584c5bc27d5422882cb4299da3914c684696eded290d;
reg [MAX_SUM_WDTH_LONG-1:0]    I1f749b245e6db4722494bb36009a7da73ca94f408d8a0ca7829b6d5258f78e4d;
reg [MAX_SUM_WDTH_LONG-1:0]    I4dcd8811ecf9d39f66ab4cf1e07e739c7972e9cf2ef9ff6c0a948336e22dcc90;
reg [MAX_SUM_WDTH_LONG-1:0]    I48c76be33e4d7a127ef1f7eb5f4952f81439eced5be914ff90aac6d963267659;
reg [MAX_SUM_WDTH_LONG-1:0]    I1a1149d160ca76d7b9db443f5095737e563a7b75de7375f9c148f4f4dbe7e7f0;
reg [MAX_SUM_WDTH_LONG-1:0]    I67e66b155579d855e0c14e91d2ce1fc6fe1d2f869e4f56b37de5f700d84073fe;
reg [MAX_SUM_WDTH_LONG-1:0]    I67a45b7ce414632252362c1556be0e627757c871c136d8570d4300fa316205d3;
reg [MAX_SUM_WDTH_LONG-1:0]    I51abe903b403df434eba534a1102cabe0a0e976c047fc5cc97a6c8e73263c531;
reg [MAX_SUM_WDTH_LONG-1:0]    I0c851ecaa50ea3e1769828a7f51da7a8c3b0c0a11eb9002b108693f09e60667f;
reg [MAX_SUM_WDTH_LONG-1:0]    I31d4c202b8434aacebdaf5a60c34d7bf3864a5a7c4707efbd1cc3dd82a9ba59e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia28734d68fd59a227094e3d5643b87d918753610e867c1d047d8878bd9a46be3;
reg [MAX_SUM_WDTH_LONG-1:0]    I735ec7a402f471520335d15ee3415e874f56381a2c0cab5c3a5b21f7d6f71474;
reg [MAX_SUM_WDTH_LONG-1:0]    Id9db55519cb1208a2555678410c950b6fb31e5fb04a0ae12d6b0a9de4d750b43;
reg [MAX_SUM_WDTH_LONG-1:0]    I4e6e6be5d9a7a85cc07a42c3a252e38fad4229a40bd68bec6728e7efa85984be;
reg [MAX_SUM_WDTH_LONG-1:0]    Iab63efeaac16bfc91c71a1a0819747c4576111221b2e355300a6e02adddb1aad;
reg [MAX_SUM_WDTH_LONG-1:0]    I0e9e95de14abaad3f4dee2c74242d09121b496fc60f22dd3513b90860e7d03ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I67874ca15a0723ab01392f527151dd5a60a71a0dd16cbbd572fc50a343c684de;
reg [MAX_SUM_WDTH_LONG-1:0]    If434186e818b5a899ad4add63d67ba1dbed823165df4559ee78b39d8c758c727;
reg [MAX_SUM_WDTH_LONG-1:0]    I843cc48bafe9c4d2e4647f2909064999da8c2f4d8dcfeaf533fcd12c32c37ce0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia6ddd4cda9a70e95a6ff1a9369bb2851b90588337f2cdad6ab43fdd6c6e32fdb;
reg [MAX_SUM_WDTH_LONG-1:0]    I0cc63aa921326ebb19427e9e06862cc0a42b375a328061bc7f6580bf3f1d3b12;
reg [MAX_SUM_WDTH_LONG-1:0]    I0c92cee9eb9e3c8300210834a106174a25005d9a468a481e0f594a960b5995ab;
reg [MAX_SUM_WDTH_LONG-1:0]    I3e73f999bb1a0c087c2d4023920d56b1525bcb43f9d1bbc1b49b57d6c9c55127;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibfb1cfcf89fe21ebca17ed6bd834fb8567cef4ccfb8f03fd5edaf59000ba0cae;
reg [MAX_SUM_WDTH_LONG-1:0]    I4878199f761be0332cf7d653cf1e73cd52f938bf9ca0f32724d499765f313d46;
reg [MAX_SUM_WDTH_LONG-1:0]    I9dd21c6b63d36e7dde6f3133ab04263a47559b648e8717de7065e7f140911d3d;
reg [MAX_SUM_WDTH_LONG-1:0]    I3db60bf522be36d36bdcc35d1d5da9cff2db6e8f89b179726fabca1a7c67b255;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic5921b5017385aa779a2016014d381a982c32c64d1643e79631a8ac842d5b584;
reg [MAX_SUM_WDTH_LONG-1:0]    I29e9674dcb3b06489c5f9017b95878c6a75503e1dc4e2ba4c9c6a7a7cd74d885;
reg [MAX_SUM_WDTH_LONG-1:0]    I6853348c8635a69100a45e6b2b255d6111daca84f2eb28629edd64f8c36f014c;
reg [MAX_SUM_WDTH_LONG-1:0]    I0bafe9c7cb10e6696f6b6dafb74a2113145f7ef1cb70496d068a61ba1de1bea1;
reg [MAX_SUM_WDTH_LONG-1:0]    I929870fcfce11dff715cf2210ad4a4c30db9af500a8d380153f38f0ea2b7c2b3;
reg [MAX_SUM_WDTH_LONG-1:0]    Id56cc1c8a7f6213208fea3ab1298a107ea854d908609dbe2358ba954989e1784;
reg [MAX_SUM_WDTH_LONG-1:0]    If7454cbad692d8d1ed806663944dde3d846b241d1f69736da66374c5e54b8de5;
reg [MAX_SUM_WDTH_LONG-1:0]    I9d23867d2eb5d9dbcc21e9242aa71e141a2ecad61f5ad2bb69d798b2fdd1873c;
reg [MAX_SUM_WDTH_LONG-1:0]    Id4f16cdf2e148fb2732fdbe215ff0edd44d29c41dff8c5b307ffcb8305832972;
reg [MAX_SUM_WDTH_LONG-1:0]    I32a7df875889c28b6d8f86a42071ad142efd5a66d6328669bcdf1901a225079f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ideafcce97c26d412480370ab40d8261f37e8bf0ba68bf7d04f4099a517195dfa;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie3cada5731ce9e6c51353952cfb87527bca19aa77436766bdcc843dd92f1cc60;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic56053af1a36bedb5e1670282ac0a93d782faf76d25a25edab3dadb09a302de1;
reg [MAX_SUM_WDTH_LONG-1:0]    If4f8191d57bfd0311981d36c3836f8da526830c6fe2dae5933650b290075ef17;
reg [MAX_SUM_WDTH_LONG-1:0]    Icc14287e817338eea415b9f8dae2527d6e71853a49869ea829d1b51aa7013dab;
reg [MAX_SUM_WDTH_LONG-1:0]    I42336bb9a452e51859fbc836c4294468aced58a32a221057096f5119d459edc9;
reg [MAX_SUM_WDTH_LONG-1:0]    I424c57a79fc220d56d1e499af6318dd2a2f4a4ebab1c83cc7762658b8c34479e;
reg [MAX_SUM_WDTH_LONG-1:0]    I89b44baf278e7cf024304d7bc6cfa759a735e5da0cf25a96a83e29fa83d12bd8;
reg [MAX_SUM_WDTH_LONG-1:0]    Idd51d2eb571b7a35413e786a8a9437a5ef34a13b84d269e29c3319a4bb7531de;
reg [MAX_SUM_WDTH_LONG-1:0]    I5b2b2323ba78f198e4c86b284772fed82ae708af1da14bfdf215a7b34f811204;
reg [MAX_SUM_WDTH_LONG-1:0]    If51ca9faad7b057d5a086daeaf1118808bbaf90b484e38571530cc3bb497dee9;
reg [MAX_SUM_WDTH_LONG-1:0]    I3c03db46b6474bbd284be2e345d2fae9939f0925a62da2ff9b1e2f3632740b0c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibc35679e4c52c119bb0ab5c5a485b11a4bd43ceba90f9998d9704d08ca3285f9;
reg [MAX_SUM_WDTH_LONG-1:0]    I9244711e562e8ea7e5e0de1921bdbbc5b64363d51d121922f441d8f36e949c69;
reg [MAX_SUM_WDTH_LONG-1:0]    Idfb0ecafd00955b66bbc43f1585659b2fd82fa239ab0274450da985354bc4c14;
reg [MAX_SUM_WDTH_LONG-1:0]    I6a5f07e66bbd7e05ab9c5adc7bdc99f269386519a6212431d5793e766239e862;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib423f5e14b109a601cf9e9d403a7b5c0ca0de8d665d065d8f317760c5705071d;
reg [MAX_SUM_WDTH_LONG-1:0]    I0dfd7663ac138a56ce3fe38c03c10675da9e417e38f56ea0fa4f9f1902d725b3;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic3f066b6b8dc09e89e9796c2b739b37e64af709758029ee21800f9fdf02c533d;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e6aa1d0b76cee0ce4862aa5d01ee91caa123335ab19a2150e8c4315c7d958c6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia261f7672256403997417633102f8c1332ae17195bc38faf0fb85c4e4dd14da7;
reg [MAX_SUM_WDTH_LONG-1:0]    I4d6d60296569a9b2a811f8064057743f13fdc60379669472d28df97061ccedb0;
reg [MAX_SUM_WDTH_LONG-1:0]    I81c33c11a5d878aea61749e54e68c024fda21f27f7f4fcf45e5b042e8ca4c3fa;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia50c90193d9c7ee51018451884df0da92f138710bf95fc32e439b39bea3f3b01;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie81fcb1c1ed576d911918860ec73a2b7823bb2d435a0477ef407393052729326;
reg [MAX_SUM_WDTH_LONG-1:0]    I2d2817ad47b56d0a7ff72c326eabc6e2ffb1819a2748ffe3a4a42d3794cf2fc2;
reg [MAX_SUM_WDTH_LONG-1:0]    I80c7df909269b691013f9d178bc3e8c896d4d06ef4cc4b0ac42858888ae8b92a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib36374f40465c181d1b8d65f23001a10ffaa250f0fd89077848e6a49a19c56dd;
reg [MAX_SUM_WDTH_LONG-1:0]    I2a9f642cd74521fb661e381a3f57eaf539ca18ff62ee2130aa94da51cd13d4c0;
reg [MAX_SUM_WDTH_LONG-1:0]    I2edaebf9e3781f53167708c4854b01219957ff020915c8d2fa7b68e50ede1d66;
reg [MAX_SUM_WDTH_LONG-1:0]    I2f928325d150ab718f3b764d3fc4e15d88af5567b4554ef8bbd02f4c3984f544;
reg [MAX_SUM_WDTH_LONG-1:0]    Ibf0c6b2fd7ba6e86f7cea34ea8434ec5353399651fae6f00cae29cfd32174563;
reg [MAX_SUM_WDTH_LONG-1:0]    I157157e9b85b39f2f22c57c4beae22472512ec83319dd9ac30075b4266761031;
reg [MAX_SUM_WDTH_LONG-1:0]    I0162ff342347e70b1361d5f3ea70c6f872d9b95ede7f80a0a18a69c84b5ebc8a;
reg [MAX_SUM_WDTH_LONG-1:0]    I1f9214a0b2b730fd678664ec457d15dcc243ba1d68ea198ef2792ac2440608ee;
reg [MAX_SUM_WDTH_LONG-1:0]    I581a3a40f892233a7bd0dda3bb84e2e46095c27e45d53ed32ef5226f9d25ce43;
reg [MAX_SUM_WDTH_LONG-1:0]    I8a3b07f660ad94b304ffecabf47d3378d3ea73b1deccd771fd1982cec9f23e39;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib1e8234d991235274c74ac026c33d868403b3d03a18a0c674e07dc4f94d614ff;
reg [MAX_SUM_WDTH_LONG-1:0]    I730afd6404f505477b32f86185baccd692e9e64865f66f048a93e33d1cac8df6;
reg [MAX_SUM_WDTH_LONG-1:0]    I30b6c3fe760f221d2861a5b6061034f6dee7320a04cbd7de2a3c728427f927fa;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia7c03e6396e5145d0027d0963c1f8b7068636ee262fe31aa442a5512e0d4e99d;
reg [MAX_SUM_WDTH_LONG-1:0]    I7fed914efeb5727bba8c1dd0a5cab385a750a2cd9215923b596d1ae914639761;
reg [MAX_SUM_WDTH_LONG-1:0]    I0cdb70836bdb3237ff43b23b1676a274cc0dfcffb214799b78ea02c2b59049fd;
reg [MAX_SUM_WDTH_LONG-1:0]    I5502a12455fae3619e0c2297d5e4a8062415aa3ddd8f0bbf67a73233bb6df733;
reg [MAX_SUM_WDTH_LONG-1:0]    I7a52610226b8a85bdc6a0b49cd74cc644d2fad0e8f98ee24c46ccd3664d0af24;
reg [MAX_SUM_WDTH_LONG-1:0]    I55d6bfb606269d9d01dc348f732caf9cfdc7042c845744b7a25c0a74d0afefbe;
reg [MAX_SUM_WDTH_LONG-1:0]    I7ba56fb0b187c50e86b74d8dfa7d7b3a1e2bc341cfb56a6343de1e7bb60742ac;
reg [MAX_SUM_WDTH_LONG-1:0]    I95d408de4742f651f694ccc8f61d215af1e9b9be2b3860dca46c143e03b3ffec;
reg [MAX_SUM_WDTH_LONG-1:0]    I446e1574b1d7bd427fed19be1920c5c29a3276d9ec816ebe1e4465cbb762b1fb;
reg [MAX_SUM_WDTH_LONG-1:0]    If2f521cf64a5e19b1f744d41d929a37a37689534d0e564224b128866d853b043;
reg [MAX_SUM_WDTH_LONG-1:0]    I58d3b6391c1720bf6ac7458ce499fe3b0573e8f7f324db1a796d1126e42e57a6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia3690db3bb1809f3df1fcc3a2dd5f807a0ef26c4cf61810b0f9bb590951f8e36;
reg [MAX_SUM_WDTH_LONG-1:0]    I0583863d43273e6464e5e65a8714be627f867a0320302382d94ef661b21f73d0;
reg [MAX_SUM_WDTH_LONG-1:0]    I47d2361b09dd6690b6b0a7827348e9e420d8b97c4b620a4e4928c8cbd84c321b;
reg [MAX_SUM_WDTH_LONG-1:0]    I6f71faa84bc155810576a85be759d7c06d84dd53b5e2dbc74ab0175e5d64d3fa;
reg [MAX_SUM_WDTH_LONG-1:0]    I403d7b440509677065b38ca8634080a8edc4c8eae54a9923c50885861866a7d8;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a8f6218aa06df768133a9b95140db0cdd600a5d1a04a2004479693cecd87571;
reg [MAX_SUM_WDTH_LONG-1:0]    I7c843a280d8a673e3c59a22f8bfbd5860c3284b189ffa281759aa44233eee225;
reg [MAX_SUM_WDTH_LONG-1:0]    I7f31f363b408908ca5cc070f150594db404279b7c5326f5da9abe8f60138bd51;
reg [MAX_SUM_WDTH_LONG-1:0]    Iff8bdf9ea44924628e777925357dcbe728f0ef4be0a3574965c811485fb57689;
reg [MAX_SUM_WDTH_LONG-1:0]    I0d58818dc0f3ed67f1e3a10ddc7cd0592bfcb8cb3db1c329edea24dfb0ffde5d;
reg [MAX_SUM_WDTH_LONG-1:0]    I16863fd89fef9bef09bbfec8d23ba6d42f4de7902a5928e9b43546b4078fbb0c;
reg [MAX_SUM_WDTH_LONG-1:0]    I1d5510ca99815d74f26804206bac7f1e7eec3727fa89d91b014becb49a815abc;
reg [MAX_SUM_WDTH_LONG-1:0]    I241e6ca6efe96759bbb20d710c448c9c322aa3345fcdbedf625e297070af52e4;
reg [MAX_SUM_WDTH_LONG-1:0]    If8ea1abf5aef298950b84058c5e76029f717309fa685556f09c32b72959f648a;
reg [MAX_SUM_WDTH_LONG-1:0]    I4eb03f5790e18ea72980b8c37b602469d6dba5f850ca3721f49279b4e14cb7c1;
reg [MAX_SUM_WDTH_LONG-1:0]    If4c7abf17850a5fcd64bb4ebaef1dc806938542a3bb2b9eee643fdfcfeec23b8;
reg [MAX_SUM_WDTH_LONG-1:0]    If15171a1904299c55ffc5b4c9059900188c1c87caca3f4807c4498abe038becb;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf3a16773d04781aa96eb511825cc59c609fc887b464a86c7839c57ddbba37db;
reg [MAX_SUM_WDTH_LONG-1:0]    I5eef24c8de2049e0e8bdd49346b6be22708a135d56c096907e50ecfbf3affdea;
reg [MAX_SUM_WDTH_LONG-1:0]    If0d87a6c6a4dd34bcb5411a845e6e7bc7fbeb0e6a34933f64283c880ca5d3d8e;
reg [MAX_SUM_WDTH_LONG-1:0]    If8c51307ae2c537425caa18b7c3dbbf0530e94ada2a2a600262f57f93bf60d24;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifdcd4016757d0cef222265289850476e0e2a6547732f999ca0cd8449f7134bbd;
reg [MAX_SUM_WDTH_LONG-1:0]    I27737e1ab6f67dba3964412127cf6c91c7a58f6ba77e5b6a9808e2775069ad4f;
reg [MAX_SUM_WDTH_LONG-1:0]    I72e85032ae85773b79f3a3dab895c9667cd32c6aeb44c000096ddcbc0f7be0d5;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic7abe3b0fe121e025ad7f7802b7800f4097111a1108ad088e869e81e5374c42c;
reg [MAX_SUM_WDTH_LONG-1:0]    Iccb7ca5c2ab8a9a4e3776ef42997d1d645c5542c25ed35b161702ce450f90fd7;
reg [MAX_SUM_WDTH_LONG-1:0]    Icd7ce463860bc6f62da8d62b71970658ed2c5d5872a56b8429d9223197ef0ad5;
reg [MAX_SUM_WDTH_LONG-1:0]    I8952c026089661f4ddd0720f6ab16e46334fc934e6775e7163aad8cf5dec6b68;
reg [MAX_SUM_WDTH_LONG-1:0]    I9efd4f4bd4d8dfa270cb1c5a2e3f5c6cbfc3c5b672540ca268e0765170e6c748;
reg [MAX_SUM_WDTH_LONG-1:0]    I4408d142165f7f5bcee86e820e4ce79b4ecfe2134d8e50809080e0c27e4e2df9;
reg [MAX_SUM_WDTH_LONG-1:0]    I29141cb56b9f52d74c42d689b180cfcfe7daf23ce573c1f4eaf21525370e5376;
reg [MAX_SUM_WDTH_LONG-1:0]    I567366a85ce4a20ac4125a297426463bc2f2c71511a97bfe2f4a01f6e8da6403;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia71d81a2779b6eb5f39fad80ee4e7bbcf394b97657cb094aec163180224939e3;
reg [MAX_SUM_WDTH_LONG-1:0]    I9beeb3f92470748db1e059cd6c5a929d1eee2a3ecd0ac097032c74f4134a22be;
reg [MAX_SUM_WDTH_LONG-1:0]    I387ea75c114fd752ced502cc147dc9ad385dbf69607c04edf81ab74b6867f2bb;
reg [MAX_SUM_WDTH_LONG-1:0]    I8d10cf5dcbbd1a765ece13156db0ad4651b41cc5ee286720226649a707accd16;
reg [MAX_SUM_WDTH_LONG-1:0]    I55d5daa0c4cb89aac08ecbaaaec1d6afa2379b277051281d3c15abaa6af05edc;
reg [MAX_SUM_WDTH_LONG-1:0]    I5460bdaa1d2a7c1cb2e75baa2c211593afac76ce5160a620b385393217b4185a;
reg [MAX_SUM_WDTH_LONG-1:0]    Iba39b0599ed448a7fdb07f6042ef972612b54c7251b256373b30788f64f616e6;
reg [MAX_SUM_WDTH_LONG-1:0]    I58db55229ca30218227b598184e85d57a0e3a8b61308f8114cd709232573e566;
reg [MAX_SUM_WDTH_LONG-1:0]    I94ba926e07e8b3cbc5429ff6bf73020e95dda7b7c0059dc10ef646b2980bd80a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia6058d7a3749f21a827ae6a0f4e792d6cd62ab37d668d607861bdf3985489d97;
reg [MAX_SUM_WDTH_LONG-1:0]    I405b2f517ad52ec3c94eb9d1d695f6fb9700fbd32fb49fca23588911b5dd0ef5;
reg [MAX_SUM_WDTH_LONG-1:0]    I0217d8dc004467c4c431dbe27dc564c042c33d06a5be72a29ceab927708c4de5;
reg [MAX_SUM_WDTH_LONG-1:0]    I14102f52e9c6fa58677dbf1260a5049a6c2807b245f123cecfc3f1a413badded;
reg [MAX_SUM_WDTH_LONG-1:0]    Id71b753d1cf473f4f4bb7718f412471692e08afc0ae9d25e617c2360df79ceda;
reg [MAX_SUM_WDTH_LONG-1:0]    I443558f78c6ebb16bcd49ca586ea62d2ba12ed3bade0e54ae9bb60f83d2598de;
reg [MAX_SUM_WDTH_LONG-1:0]    If5c2310896ae5dfd3f83de1affe79fad0f0b6b2b673efbceb7d296b33a6900e7;
reg [MAX_SUM_WDTH_LONG-1:0]    I7d078740e07b48774c64f6dfd7bb0f56821dd685e014f0b9d4e3b7da45383e34;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib3562b77830a64f31728e11cc54a6d19b55344891eb82355e3fb4491086e8808;
reg [MAX_SUM_WDTH_LONG-1:0]    If7d42431922752de30d5506e1d501f65453a4754d7cab03976695cdee9c0c9a4;
reg [MAX_SUM_WDTH_LONG-1:0]    I269a90aa42086a30a9b03141bf37e3abea46a1f1c06710baf2d052a5bb404248;
reg [MAX_SUM_WDTH_LONG-1:0]    Id88de8b0cefd527c486f8239ff6f61d6ff86085e420d2be56ce58f4d82d78a7a;
reg [MAX_SUM_WDTH_LONG-1:0]    I107db18dddc718b9fe7354d0f352f72df94ad4653ab0712d5765a495ec29242d;
reg [MAX_SUM_WDTH_LONG-1:0]    I642c0e5f0768f835a6ca3ee6f65875346121b502770acb1ce833e9aed46d4ddc;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib699efc076bd227e0138482c43c5fc8cf0d0d87078e063262fc4b537f554697f;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e0d77d4d38cb3b1e5ece19e010043e9a4f0802819f3e70f0ecc9440f65eff4b;
reg [MAX_SUM_WDTH_LONG-1:0]    I3eaa094e28f19bdbec184b0ba0f3792f90e67c77bd8dff9af6042c5002735505;
reg [MAX_SUM_WDTH_LONG-1:0]    I62b9322a1d5ff38480981e00d8469983588d084289f2f927f3339250b5c35985;
reg [MAX_SUM_WDTH_LONG-1:0]    I2af0f38cbf134ae07c76f06d4aafee537bcdfe91b1c4aff1ae27898e18da5113;
reg [MAX_SUM_WDTH_LONG-1:0]    Iec6be5ba578c849ae0e4fee9c059ff88c36cfa7c14cfe218cad7f7f1d6744024;
reg [MAX_SUM_WDTH_LONG-1:0]    Id18c335cef6d5d988e55f6fda5a09a24ee80f4d4755f797a11ee94141b69b97d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie85ad3f88a177d67b69eb3a03e4a9d92f7431af9de9ccd06f2caa01f9d144f33;
reg [MAX_SUM_WDTH_LONG-1:0]    I53e788aafc97015db67a8363c91d81d369d80c4d24542fa45faf7833fa4189c1;
reg [MAX_SUM_WDTH_LONG-1:0]    I8f74cd611f5df70ef183e9d4a86b5ac23349be8cb99cd470c596fcaa6ec95248;
reg [MAX_SUM_WDTH_LONG-1:0]    Ief3910aa326e0d9782566c81ab1cbd09faf46d3552f78d7ef5fc9de1d9c245d6;
reg [MAX_SUM_WDTH_LONG-1:0]    Idddd98e139a087c7aef3922ea2542dd364c9d30f70665754f751ed88dfbd3701;
reg [MAX_SUM_WDTH_LONG-1:0]    I474f7c67e6159d041be6d6f4f96fe58f9b7086757936ebbc86340bcd9cd9962c;
reg [MAX_SUM_WDTH_LONG-1:0]    I2a1c16f7d4c3261619c325f4b5cfe98993d5957a2ff466bae11c9cec6006cac6;
reg [MAX_SUM_WDTH_LONG-1:0]    I881a2d7025d422202455bdff165dd982c2f4953b361f29688e75ccdf9e04d476;
reg [MAX_SUM_WDTH_LONG-1:0]    I8245c1ad016aa3d7290e1097eb966b09c8a38fa5bf62bcb7ef179f448104f47d;
reg [MAX_SUM_WDTH_LONG-1:0]    I10206e80304f6e623a256b6042ceca13c691a34ef5b6d67667ab4bb11f0b0087;
reg [MAX_SUM_WDTH_LONG-1:0]    I50f15058dc2e50a994089de4a0487158352c882d4639449d9db322a05ddcba3f;
reg [MAX_SUM_WDTH_LONG-1:0]    I0604d25b233f4206fb580d729452e9694d4b795553a4a788f993c992bc433b0b;
reg [MAX_SUM_WDTH_LONG-1:0]    I5b2860f88d7cbdbc92264ca1bd0f97c610e7b1cf340e2b65832553a1762fc865;
reg [MAX_SUM_WDTH_LONG-1:0]    I62f27f0dc53be101d8fc7f026a673fd33a5397534153859f45c113e6820e9c26;
reg [MAX_SUM_WDTH_LONG-1:0]    I92cfa50424ddf1ada795366ac6c7b31cbb1b1330486911824b881a1fda443c25;
reg [MAX_SUM_WDTH_LONG-1:0]    I1d996fec699e93fc4ce63060990c6347d998a81f0b3aefd88339d5d620fd152d;
reg [MAX_SUM_WDTH_LONG-1:0]    I33546fedf41dca9168afd7d6916823e8c24aa3c4a855b93820215c68c807a56e;
reg [MAX_SUM_WDTH_LONG-1:0]    I8617f958a4de5cf233240840c770360befaafe599fbec1e351b24baf301ecdbb;
reg [MAX_SUM_WDTH_LONG-1:0]    Id824ed4e68ef3624b9a4d6c5924b08a7b727df62fc9135c973c5f79768c627fb;
reg [MAX_SUM_WDTH_LONG-1:0]    I3d71ea5bb4c4be8ea80abe59367519a071132c913eaa5c6538baa8c3faf243d4;
reg [MAX_SUM_WDTH_LONG-1:0]    I6adbf5489cbaa65213fe0804e7494a2b8be9db9132a6ab7058764a1a53480999;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib4e392b7b8f87358dd5cdefe7c272531bc6bb1f27bf1411c1a2f4331809a83c5;
reg [MAX_SUM_WDTH_LONG-1:0]    I6b528ad76bac25170636a86ebaf7efd14ee7159ea2c83500021e39e968786428;
reg [MAX_SUM_WDTH_LONG-1:0]    I294be7c0765f0d4209d4442136d706edb2080883d5c78a3c71d66b5946116bef;
reg [MAX_SUM_WDTH_LONG-1:0]    Id834a34ad825df7c595e3754b5a5638badf560cfb68ec8de2903e73e88b1a113;
reg [MAX_SUM_WDTH_LONG-1:0]    I09e3897931014e7bd9540023eb8fe1097e36eb5c51db24357b492a132c3a8805;
reg [MAX_SUM_WDTH_LONG-1:0]    I674ac3fcd5872491a3c412a02e367a9c29e4dac14a8ffe8b6382c60a29fde8aa;
reg [MAX_SUM_WDTH_LONG-1:0]    I9ac796f1901c19aeab344ea2c785af3ce41bd23dffe88b1b5216f8f8c0b16e40;
reg [MAX_SUM_WDTH_LONG-1:0]    I0d186e0127f200b704a4585b2fc43ff1a9ab19833a90ac881abde94b2da89376;
reg [MAX_SUM_WDTH_LONG-1:0]    Iae8191d31be3785db5d8e5d328fb2d96b0b5d5ecc7f9d14f0bdd3f61a9bb6781;
reg [MAX_SUM_WDTH_LONG-1:0]    I4694c593512d9d84542af4ca5b0f3022f9b1433d7d6435ffd4b1e53093bf4a58;
reg [MAX_SUM_WDTH_LONG-1:0]    I78c5059e528b7671e27f847d6042b3fa707258c664749d857004679c6ff96a73;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic83ed3610853814d7c9d6932b644f9c924fec7d67e303160a3c5b99c625634c0;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie33f8884c8fca47e2055b28f4398f3207f7ea20f8d0858d2a0699ef2da5a8f03;
reg [MAX_SUM_WDTH_LONG-1:0]    Id140833a04f0b4b903ad4e99046b17f76d4c405703fba227d36342b6f1fdbd08;
reg [MAX_SUM_WDTH_LONG-1:0]    I90d7a3c4ac0a18444eceec2569cae3d5dcb3d33d2e46c329068b0d35ad063971;
reg [MAX_SUM_WDTH_LONG-1:0]    I5c7c7df860c87ada06c17210746ef84d27aabaa26e9cad20397822629716d4a6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieef9e0d39f2e213f365af4a6a34d0d2c7d50155e8052e9b1944473641922e9eb;
reg [MAX_SUM_WDTH_LONG-1:0]    I4771e59053fbd3e261c49e0be7e742e7cf9c5bdad030b67f1b955e13e9bcf083;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic8c13812ba09457021ec6f39406b1106dc025551c62da4259930c361f19c3a2d;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic7aae8edebf83f3971440fd0e86e7700ac4cc0c087c9996d55cfecea8c489fa5;
reg [MAX_SUM_WDTH_LONG-1:0]    I091bf548253a3b22f92aca6479b70ccb74a5f9eda8bd80e6bc1e059021f04b9f;
reg [MAX_SUM_WDTH_LONG-1:0]    I5c1c30033bd61b271c765ba00b033a58c6389d4bd353ce68d1b193bc7138baf4;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia4370635785f2b904fb6ab3b8cdb86fba5445230a9d3d02cd908e04d92726f3c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie73ab4d16ef614a27522cdfd47f670a38ab58f89bc10c74975cf0b30400e198f;
reg [MAX_SUM_WDTH_LONG-1:0]    I76b8cfe5d3985f3c0f249680ed81aa3b21cd7af725925846e8875ef9e98a550e;
reg [MAX_SUM_WDTH_LONG-1:0]    I58919d58783467b7ad0108f86d6260f3c551692d00e6639260a68a7a512d8689;
reg [MAX_SUM_WDTH_LONG-1:0]    I0d276f9604ec2b8621a86706ad1772058a29e94902e8eece60e3d07948e24cee;
reg [MAX_SUM_WDTH_LONG-1:0]    I5463c05b1b55c142012470d627accadd8e34924e77ef6d139b3fbe1db1cb91e8;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifca2987d8c7f1ca30013ddfcdb82a888ebbd7bc3dc421f7e3d6806f5f3a9aa2d;
reg [MAX_SUM_WDTH_LONG-1:0]    I5ff269ab544d2b74059a73d0ffe0492473b214d392d8c2ee760847e6c07a361a;
reg [MAX_SUM_WDTH_LONG-1:0]    I26a6366fb57427f6a0d87d4cff8a293a0752887e71b829e747c27980a1a3dbbf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieb5560e3a4f6a9c4543d941ac57bd3805afa7fa17624e5739e8e639e8d0d0c5f;
reg [MAX_SUM_WDTH_LONG-1:0]    Id1b9b5118024dfae0e058f5418c9e988e0a5a598ef7553947de6f92cd7399201;
reg [MAX_SUM_WDTH_LONG-1:0]    I50e1a6fdaffcdf8fa99074f4480dcc21971ba8f5747b24a33232f9152b07af1f;
reg [MAX_SUM_WDTH_LONG-1:0]    Ieb31a59d63544ea160d3934f0e38e6333f8571e77352bdbfd338d68c437f02b5;
reg [MAX_SUM_WDTH_LONG-1:0]    I81e45b654bee6c74edb5e034c89bed7151c60a69b554a35710d1b173fe45ea22;
reg [MAX_SUM_WDTH_LONG-1:0]    I5144a2cef7d82b7a91f9d83ff8fdea356bb01db215bc167f0c498d55d1faa622;
reg [MAX_SUM_WDTH_LONG-1:0]    I67484837f2e585fbb85de404cad8f08ba58bd1faa81b9931f88473d7f4a9a06e;
reg [MAX_SUM_WDTH_LONG-1:0]    I4404bf7e923ee1bc0230835c00684d298572238aa8b9602dc48e177464224a53;
reg [MAX_SUM_WDTH_LONG-1:0]    Ied796eff44d61681c5d5de05933e785d387a97b2430fee26d96b0b24a1a54c12;
reg [MAX_SUM_WDTH_LONG-1:0]    Icd8838ebb43dad19fa96e741b32851dbaf5c469e0591a1231898a7aeb6ecc788;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic6d60bc06b0eb51b5ff4b8cc0d0ccf55fd8e5c53aab23b3994ca8d094920d619;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0feb2870e46760bd3c58e5af56a40a73fcc6c9611766c77c4784f88c35f440e;
reg [MAX_SUM_WDTH_LONG-1:0]    I60b4f2cd3f513ded6891a6506d0ec74357660440c94e62f4f7e2f886c1233204;
reg [MAX_SUM_WDTH_LONG-1:0]    I90b9d06240e2a49693ac4ebe37203439a157a38d068e630c45341d7d677b816a;
reg [MAX_SUM_WDTH_LONG-1:0]    Icc84144f0fef09379e456de5410487e7882d373874a686f1b61db92511a91e2a;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib5ba52b9ecafcedb064e66c38273f7833d0b6d0239a7fff9ef3a0e30d0f77dc8;
reg [MAX_SUM_WDTH_LONG-1:0]    I38a6e64d23e0dc1a449445bf10e786777e978aeab68b3a99dc5335b93c67da45;
reg [MAX_SUM_WDTH_LONG-1:0]    I83b2a186b150fb7290623bd1cbab9d044e9b5c760ed36ae218fb775354e46fd2;
reg [MAX_SUM_WDTH_LONG-1:0]    I507512179a289ecb7d9ddf5e853bb42798df8129655c06e568e0a4a1d880ef71;
reg [MAX_SUM_WDTH_LONG-1:0]    I6182a01d42a30ec5e8883e7d4f5d8f1d657f78052fa4c8ca2c160aecffda456c;
reg [MAX_SUM_WDTH_LONG-1:0]    Id645d98c8a2ba63ba9060280b1810d0ab7120f007f3f174e1a501a1f487190a0;
reg [MAX_SUM_WDTH_LONG-1:0]    I6822880688515ff8108fe78fadc5d22b953ce5face9928836f824aad9355a713;
reg [MAX_SUM_WDTH_LONG-1:0]    I694ec7b5bec025b308c4cb56eefedc2be0842202dfb047b5a94dc749c757bdde;
reg [MAX_SUM_WDTH_LONG-1:0]    I99a4bc7f129030d12eeef0507cf52503af3df70717d1ba9c38b5dd3a5ffcb616;
reg [MAX_SUM_WDTH_LONG-1:0]    I668aff5da6360f719a2467c5189f3e53e8eeb310f4c4e26f55f8c39e9dcc4be7;
reg [MAX_SUM_WDTH_LONG-1:0]    I4583579034ed3bcee2ef0ea2b32a4adf0467f78a2770a84da9948e8d366c1f4f;
reg [MAX_SUM_WDTH_LONG-1:0]    I86729a880fe730068d538da490087a1ab6789327f964722c9c14bd9b1c2af35b;
reg [MAX_SUM_WDTH_LONG-1:0]    I0f8046b4f96acee2bfb4719bbff91b4b1b81c78ac36ec6e95008a3d9cb5ea6ff;
reg [MAX_SUM_WDTH_LONG-1:0]    If08c85e70828c39162bc16d65747d3d3d0a6176e8db106b262bbadd651f745b7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia0ee127b17b441cc11d664edf15d370368494e31b52c4865c97a065ef8bc43b8;
reg [MAX_SUM_WDTH_LONG-1:0]    I8c494bcba3ff73ff29d9d388708fa34caa73b883730349aef6c2648a2f5a1409;
reg [MAX_SUM_WDTH_LONG-1:0]    I7ea6f607967e7d251d71b4c4b3dd545a4a9ae8298c3ee2356bbc16ebef06cb2e;
reg [MAX_SUM_WDTH_LONG-1:0]    I215148c89dc37a59b3eaf2f38679554281379dc6c8e57718e1c22c091f4d76cf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ief3b5e8fee2d099a90990de9303f34d600235d989d25a30b5a7e2654c18b5c3c;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia2233f4704a9724ec75efe5e31af6807f8f1529f641ec05d053d6a12308f485b;
reg [MAX_SUM_WDTH_LONG-1:0]    I6754b9c9cc470509e67ba88c2669e1f70666489af9ca14de9fd4e4328d18e245;
reg [MAX_SUM_WDTH_LONG-1:0]    I133d5432ba2f64f1ad612b2505fb95ce91962b6ac761dcd0e92f75d1b663d7b6;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifb664074b1a8bb954cb940a11ae4e7de1278edf3614b861ccd83dfaef95319c2;
reg [MAX_SUM_WDTH_LONG-1:0]    I76ca3c17438c05fc53f6f7075ff7404c0838f62472ffebd41a61afb1f3ea5dbe;
reg [MAX_SUM_WDTH_LONG-1:0]    I27ed900fc3d84c4ab4570c3bb88b5e9a7077389e5fa169cc4e1d606f09c9c755;
reg [MAX_SUM_WDTH_LONG-1:0]    I3ef4c55a4a3281a468daa3233ccdbe660c46a930220b5c9bd3caf6041008bdad;
reg [MAX_SUM_WDTH_LONG-1:0]    I9d323aa17bffd7ea7a66ef99d4d004ce664a0e7e5388ed24a4d45c69a4d9b396;
reg [MAX_SUM_WDTH_LONG-1:0]    I8e6a3df905c8c5778e1fd6e75b091c545389651762d9cb3e0d21b20d8dcee6ae;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic935d033e29fa4baba415347d379eeb1645c65388d3c7c9858ae48f5a098e2bd;
reg [MAX_SUM_WDTH_LONG-1:0]    I1f212ee134daea9d568f52fcdce6452048326c2dc243c60d25ee71b95ffea50d;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a25f0d4a6f0fa33f493d9aec6fc7a318a826b3885a3cccf04e9b1a85bec345e;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifbee83b3613941d8ba27021c2fd37d0990a8af8fa3e0399f0f1f8a92ae18d273;
reg [MAX_SUM_WDTH_LONG-1:0]    Ia1c056993094512262fa3f3d38a2a46cd43eb08114e1af8c48ce2f6705d7297b;
reg [MAX_SUM_WDTH_LONG-1:0]    I61e29bdef580f4f1057d7b4ffb5bbf37c67d3b8107d7979c2fce643282c7d861;
reg [MAX_SUM_WDTH_LONG-1:0]    Ib07a3587e3bfa70ff5dcb296b8595c5d15cb8a94efb13c3e5cc92cd3be3605ac;
reg [MAX_SUM_WDTH_LONG-1:0]    I8c443a2690956ee9d0171ca05534d698f75563cd74ec9f4de33c7e8dabe8105a;
reg [MAX_SUM_WDTH_LONG-1:0]    I5dcbde9462714577263040534f0560b0c126ba001e959add92d0529cbc94bd9b;
reg [MAX_SUM_WDTH_LONG-1:0]    I3872eb448ad521cf99b3a9d07ecde078320dcaaac45bd387137deaf5dec956b3;
reg [MAX_SUM_WDTH_LONG-1:0]    I144443166f296f7fdfd616492bb4b1fe44e0353fa6b0fc822b3aec0c1ea0c894;
reg [MAX_SUM_WDTH_LONG-1:0]    I5445f1e35f9039ef623a77ce395c2a888153749fe8226e9b844b271c1c69d760;
reg [MAX_SUM_WDTH_LONG-1:0]    I5d9ebd6a6829c49b0e41f700d29bf8acf06a5dd87192846e5ca204ea8bf563eb;
reg [MAX_SUM_WDTH_LONG-1:0]    I7e26d67803410d5079a43dbf6053aee09ff9b0242133282679c3beffd05aae02;
reg [MAX_SUM_WDTH_LONG-1:0]    I685960b47e49f3ff64eca0e1f26387605e48d325d533550beca6bd6d0f3abbd3;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf75218ad23cd1505d2d69d09c0305642a8be48b8a3b7aca4aa4d01a564ddebf;
reg [MAX_SUM_WDTH_LONG-1:0]    Ic9adc8e66938cafc1f6974ab9e2fd71a29bcd6520e6fca93ce7bab4815494ed6;
reg [MAX_SUM_WDTH_LONG-1:0]    I4f8e5bee14ab1e584593fc15140a36cf071f2949f1bc86fc3fb7dbfdeea7343c;
reg [MAX_SUM_WDTH_LONG-1:0]    Idbadcb95f603dca2fe62a931973c10429cefef4d6cad0b8e46cf34b2f7c7907b;
reg [MAX_SUM_WDTH_LONG-1:0]    I9f94e32610a6e83f5ca5d8eb0ad81277c7226ae8ffa7f1e734959a614bf1edd1;
reg [MAX_SUM_WDTH_LONG-1:0]    Ie023df7145a8643ec413fd62bad9e4dafc719f7c882ae969eaccbce255ca7748;
reg [MAX_SUM_WDTH_LONG-1:0]    I3a210f2cb408bb61efba033b0ea8f1cda9a3341500248e1443840c24dfe04cea;
reg [MAX_SUM_WDTH_LONG-1:0]    Ifd9d392bdf654a9146eebb9a670b75f4d74807786708350ceef7c79d54805ccc;
reg [MAX_SUM_WDTH_LONG-1:0]    I3cf51d0ae95d4e3f7d0809785f84c5d25153742e5dd0d370235828d4f9c0d1cf;
reg [MAX_SUM_WDTH_LONG-1:0]    I4fc7c4344699ed94536cb79d86f697e9da22498a2938b10360763aa9bad9da33;
reg [MAX_SUM_WDTH_LONG-1:0]    If7b4cbde972a67fae839c5bc9ddfd64dc244041f6dd60f95c5329105ae08e460;
reg [MAX_SUM_WDTH_LONG-1:0]    Icf608ba43019dffad0c708d49076088f2a4b5e126e76b3b2fefa5a0f1edeac7b;
reg [MAX_SUM_WDTH_LONG-1:0]    I0a5867bf6971ed11db3a6dc9af8cb356352990bbc3032878e82b6cb2ca8c402b;
reg [MAX_SUM_WDTH_LONG-1:0]    I56253c88487a75fb5f830a66c0dd3172ff25795a2509eaf5367fe045f9e12b61;
reg [MAX_SUM_WDTH_LONG-1:0]    I199abcfe7a0dfbaa58ab1dbbb16223bd434b4ce5ed3a65633d506d668aa76f8c;
reg [MAX_SUM_WDTH_LONG-1:0]    I2ff52a8e46c22b626ca488ae87c88360d413ad08dfaa6701fe7b237d42c2cbe7;
reg [MAX_SUM_WDTH_LONG-1:0]    Ide088b881c7dabf6e2fab61eb4e5db3ea3750d7b72eb26cb79877bc23429efbe;
reg [MAX_SUM_WDTH_LONG-1:0]    I5df56a6a00d4d8ca1c6b1a79e5f0e674482cb9541d86dd49c2ac361d86dcea1a;
reg [MAX_SUM_WDTH_LONG-1:0]    I16b3b3cdfef91e9cd5ab763bbcbe2188e61f45183118f5c735eff60965fe4138;
reg [MAX_SUM_WDTH_LONG-1:0]    I78e49a2727c2f25a14e0f8937e6241f54246c8f42a643dc569f0249384909fb1;
reg [MAX_SUM_WDTH_LONG-1:0]    I6563fc7a6bd595720441778baa975487126f50343c92ccba99218e274cf40336;
reg [MAX_SUM_WDTH_LONG-1:0]    Idc94a4d308c2e301c3d3524f1e20817f9b666827f340874b5adc763970f2efdc;
reg [MAX_SUM_WDTH_LONG-1:0]    I3167835472a3c4db7f1b7fbc1895c44e547122e9ad273066e6bdd43bccde11cb;
reg                           I94dc663f1bd5ef375a365e9407e700bfb552748c9608227592046d149ff0ef4b;
reg                           Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b;
reg                           I2009e43b9f7d79470526e490ce29be9e5d932a3c25647eb8e903114c5696298d;
reg                           If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458;
reg                           Ie6f0821795a2d09a9d5d9fee0deb445f74581e2f81076cf0395d62fcc7ecd5c9;
reg                           I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0;
reg                           I47e3e3ab4fcba3cc4478ddd5e0ff92bb41fc8fb0403411b2b588ca51686b978d;
reg                           Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e;
reg                           Id11097cace1e3bda4cdc1e833708180e784d09c9fbea9e735a2ad96e473e9494;

reg                           I6d0b0c1a3968ec36626f19660bedfe0a538a7835edd2a21dd3f4ce0fe2c5c86b;

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          I94dc663f1bd5ef375a365e9407e700bfb552748c9608227592046d149ff0ef4b <= 1'b0;
          Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b <= 1'b0;
          I2009e43b9f7d79470526e490ce29be9e5d932a3c25647eb8e903114c5696298d <= 1'b0;
          If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458 <= 1'b0;
          Ie6f0821795a2d09a9d5d9fee0deb445f74581e2f81076cf0395d62fcc7ecd5c9 <= 1'b0;
          I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0 <= 1'b0;
          I47e3e3ab4fcba3cc4478ddd5e0ff92bb41fc8fb0403411b2b588ca51686b978d <= 1'b0;
          Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e <= 1'b0;
          Id11097cace1e3bda4cdc1e833708180e784d09c9fbea9e735a2ad96e473e9494 <= 1'b0;
       end else begin
          I94dc663f1bd5ef375a365e9407e700bfb552748c9608227592046d149ff0ef4b <= start_dec | iter_start_int;
          Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b <= start_dec | iter_start_int;//I94dc663f1bd5ef375a365e9407e700bfb552748c9608227592046d149ff0ef4b;
          I2009e43b9f7d79470526e490ce29be9e5d932a3c25647eb8e903114c5696298d <= Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b;
          If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458 <= I2009e43b9f7d79470526e490ce29be9e5d932a3c25647eb8e903114c5696298d;
          Ie6f0821795a2d09a9d5d9fee0deb445f74581e2f81076cf0395d62fcc7ecd5c9 <= If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458;
          I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0 <= Ie6f0821795a2d09a9d5d9fee0deb445f74581e2f81076cf0395d62fcc7ecd5c9 && ~converged_loops_ended ;
          I47e3e3ab4fcba3cc4478ddd5e0ff92bb41fc8fb0403411b2b588ca51686b978d <= I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0;
          Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e <= I47e3e3ab4fcba3cc4478ddd5e0ff92bb41fc8fb0403411b2b588ca51686b978d;
          Id11097cace1e3bda4cdc1e833708180e784d09c9fbea9e735a2ad96e473e9494 <= Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e;
       end
   end

// `include "GF2_LDPC_fgallag_inc_all.sv"
// `include "GF2_LDPC_flogtanh_inc_all.sv"

function reg [MAX_SUM_WDTH_LONG-1:0] I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af ( reg [31 :0] I24de34e5237762ee081db8bafa630c1f9d05a34a83f96a2eb34811d098d3f5ec);
     `include "GF2_LDPC_flogtanh_inc_inc_all.sv"
     flogtanh_sel = I24de34e5237762ee081db8bafa630c1f9d05a34a83f96a2eb34811d098d3f5ec;
     `include "GF2_LDPC_flogtanh.sv"
     return Ica91d9bac0dd49c3d4a33cbeec278026d5f4b3f1e4fdf2d3d75f4d666e11a0b2[0];
endfunction : I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af

function reg [MAX_SUM_WDTH_LONG-1:0] Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f ( reg [31 :0] I24de34e5237762ee081db8bafa630c1f9d05a34a83f96a2eb34811d098d3f5ec);
     `include "GF2_LDPC_fgallag_inc_inc_all.sv"
     fgallag_sel = I24de34e5237762ee081db8bafa630c1f9d05a34a83f96a2eb34811d098d3f5ec;
     `include "GF2_LDPC_fgallag.sv"
     return I2921115a104a4c6799b85673837b12992d6251292ee3f5f63bf7126c12eac61b[0];
endfunction : Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f




   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          I96fb06aca6108479f7e21e1835a091a9060c2925cc6320c8ed71a0a0092bdeab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie000dee1e3953811fe9424588b71a7dbc88f41ec69afd16e17e8fabf141c31ec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie873b138e19cd7f7e8afa8bd8f8c4610b65d0fcd647e76d880d25f6fe36c54ef  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8ab1772a3bc752331b0bf62069643cadb48bc13bbb06ad3eddc68ac603d73654  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4bce49360270b653e45b914c493ca8e5b74beb0b6b85838bb3b54f1f39389fe3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibb4ff9ffdb2771ff640bf958798f8447a0dbcf15ed0ef9f82068826ec621de77  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia4691d32d9e84827a250e0b3d6ea8142c24c9df4ade01c19583e6cfca06cd990  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3a1380b85cc7f797ff92d02b7081d1ec3ba069aac74162ca059c399daa10690d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I14919dedf2b4d4caae8efa1726435d1946f48e1e9b1052133bebe8affeb3556d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I852a201bdaecd968b6f9c9b6bd64dc8035a17fb92ffc806a690781666354b069  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I345c0aef41ee2863a96a076a78d92c7498f50ef90e82e75565df1d1f38a08161  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifb94a220081758ce91634fef64be084898a662f7c0e8cc9f86859bf3852b3efe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5f1b294a0702ab37f94304ae67fe91abc04c397dd682d371126a7ceacf7c43ec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I81aa911c9f6f4bd88314aa3c5310efef6c40219ca93521bbea3c1afcea7bb48f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I97f674eaee005fc7a54ccb648f5a0a67cec041e895d62eacbcc9a37068b912a7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7628fd0a5ee3ec547c1b4798a4d76de651807424cd18f0b3b8a3bea849e6fe0d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1d8a992801d3f6a457848578ce286b496d4e2a69937344bdcbab4e8b1af1fe4e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia28f68b737aaaaa6b98aa5e9696b937e564754edef217740c414c16fe2e485b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I099e314496f03784e5504a35292defa79dc063aa81e6aa8764802f7fe3a47114  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id4bcb557769f043a7275ab01d6d9794d4cbbd9309be38f58acc307a1e693f347  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id1bb830ea0f92a1c0ed0addc915fc85198e4744c4bf7369b4ee1f7131f5f8542  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I31009872a3e84f78bbf1f12a7da708c45e3b708bd943b6f4561ad436164b12d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idd9957e5b52c4d33e24910559d8203415afdf467bbe1c9de950145282c7eacf0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a09910e62aa0cf665f69be80c9ad61f2d31115012314b8188cf79fae365626c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3d6f6b104bd2ffb35ea6782748bb777ec7eceae47ef2e1d18d37d1677d56cb80  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id5055b759fe480d476c4bf08c420a5dafe9e65cb03c6d6991c1d225af0a51d7b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I93e543ef3d58bc8bd48a279299dadae1d7f4528c3d09d7106b969e15565d3a15  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib6ff050679c6366efde7b9809fcf42051f107c18863bcea79d41b5fee0603e9c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iba81256fd46cc69f1367fc6ed7b712d2695e099c52b476f9b39f0a13404dceaa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I608b794037b45c46a29ea01e378b63a1f267c4b489b0866fe2f6090936fa9d44  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic48347f5264e8e479996a8dba0171a108b602be1e1d24b2fcb43cd2bdb82f61d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib62b5b3c80d193b97bd6b5c0d5678e424026381949c3f24546d367df930cbcae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia7900b5a01cfc1c4db79ca653f072956c13e2040cbd94cf07de2f1d969222fa8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1aa136009f34c39a8dbc39b4444642cd09c9cd2f01bd6310287d4ddc9bedad85  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic195e053a186bcb0e653c0ddec75c57d1b3210c583162dd90978858c98fa53f2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic859d34db6baa83e73a8627c251c877e93f15653973d0634c42a8ffc9f628bae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibeb23788ce301c724494a2852312b38344c27416a5604c0145fa330ccd1f290d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5ccf8e87b0b8e8ce9bdf4b3329e4458a628f2568184f82b998ac62ea28bc0307  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaea7277e745e05f803325e0f19dbc5a54234878a9a3cb2cedcc013e3942e9cc0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic94e7c887d7f24b573b470820c36fe8a0fef750e2c46675f8867d78f2100f1f9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifa0b8243f5ab6adb88a70fc1245e3480ea3fb3f3af846fdefd0613ca91d7b122  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia00cd24df6e6b22b466e1492500f1948b3ba3d70bdca407d1c22b4dfaf374eb7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8b41f817a4008df0994e2efa6b33eb847e82b031082f90a767467ffc03cfdb93  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8d91c857f2c8154bb09d456ff73ebdf81e3b7d9bd1c57c2e6b8c2de74e55cf48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id0f930aa222bd91b8a7d5f80a38d84993a63fa1c6aca3d37ed259294e08869d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I58598429d44ad951f91139a213d3b0bdacac6d71f1b9753886dfe1d39d0024ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3cca3cf08c967f80e7e255a590bb9c442abc535cd529f7ff304f25d5519dab04  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I42d1b7202048c81ca3a8bba0dbbce65501cb7a519fde37085c68d01db7edd635  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I07bdf8f629cfc9c094023be167a717880dc3a42099b01bffb431036521cd6019  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifaa925832248fd0e2f5841096d9618c2fdaa3c63a3130b57f493782f96473088  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c22aed0ed8abb0cb8906a35a4d44cfd7cc68b2924e474680a2eb6cf7caf5582  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I31ca3705bdc7e063c61023d93193b3ced40cf440afd817d0d730f6c8d37f8b92  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I789461a909fa4abaf3840dfca4f63bfa63fdab389e149fddb7d8ae2b876dc912  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ff3298d93471156b56cfbbea17c8dc0405bfe8654e9f830bb33bc6c9a649b3e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9eb30c75f8d71ade925633d7c8bc6b948ae519cdff33ddb885761bf72a8b0869  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5456c559bdce4d65af540e4c71c19e44227c62e5c129b7de968ac7f311dd76f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I98e4b84e98742d38b206ac059ad123966ee63903c616b9c31b4ba9615edb9f40  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I40d7eae63827c6efe2ac480c8eb9f8a8f77bbfa845caae02d137397c9da822a9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I30a9d5330fac5c3ec7b63cfab0edcef0eda61dddb23d2aabf733b9982c12b4ad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icbdf29918b91006ffdc8b68c707840ee6bb9c27779dabd372e2033888743409f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7f6b89a61d6313029102fc48e92a54ffdece30e9eac1191d840c488be69d8223  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9471414594b824d60836981bf4b9931c135520ad1ae7dea177e0bc591c2572c2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0e9135a0817e96971dc8c4fe6eec717a563c44738f7e38d5bfb2f4dda8c77876  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0847713503570d7ab3efee12577ba27aa81869a22b14ec8a244fbd4665d566f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7b529f16d1499766369f75cde5a356cb12c06d21f42a10932edc6d54146735a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1b93b1b2c5f55e2267a4deb4f75ca91039d6893af8e082ea85b7a5e9354117e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7200758287b0c7ed92552ced989756e1d49b5418181b9e36421da7e2694ed3a2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I96e7a523360a0cc0f3abfea09a566658e5e9f3316c3c412f99fd6340d1b64235  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic4839247bb24d460ee6d963d31fc390e8d9d679cd73f058d94ec34a18ceb39c0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I23ef4f4232fa0d8813a25ddca38a2745fb660c05dbe9ddc2cc33c47d45b3fecf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id5e78e4ed6db0562ed51d1da1f34242f54def8255088c3a1ccf0221ee8fa153f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I17cdc222663e370d6ef2539ad03c45a7949d9606583c17568a24c528a3e8c12f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I65e452247faa2c9d6b01dcbbebd5e8c31884c88e70dc8ec76d55aac7e77e2d46  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib0641eb8fe554f69ebb57e8e900f995c07bddadffd25c01781ba234b87af4a94  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee9c2c6a9b8e84402eb1e0de611c1cb8ae1e802226f2c07833bafaba74f1ac15  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I443435c78145236b927711299e8bedd0d29a743e3784ac22f70b2284b6be11c1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a86387a3136768ab52d320fae7fe63c7c74bb5541d18889faa263c71b2bfce6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0c4bcb29e2939b889fb7a5a7b62b49a3eeb3ee6f4555518c9059cb34dfebc7a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3de9fbe37d08009f5fa66bf7c59debe7da836dc078e212968afdc608b100e3bd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7c6d90cd79e1b85ce9a5452570cfeec8faf9ce3e6bc886f66495ec2a66fc8c7e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I57d80f41498f8d7b91410dc02e646a45a3f05d45e9b5871ae95d6432ecd2af56  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ief90cf0b0997823c3071eb46b636e384077579beae3d85d29e639a7719763396  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I295d7aef060ca978805bdf65138e5bf134551eda9c396a22165a77a3091dfd28  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I73a855a590363c762c34008e77f73f961950c0dd71b795acab3adf40c4540453  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie38c638da580ca7d25fc0754497163d0369f31a6cdb4bd26663a759b74efd588  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c635a0b11af3be4774428af79ff5cbe6a32ede6ad03ac197ecbb3ca2ba78f8f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I34a89a8aa68b1657dc7137437574877b170659ebdbcc93a772989e2b8b5be31f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9f9d895211b42c2c9d491349dbe7aafbad775942920197105c34837dba6563a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11c6d693bd6c019722571e1aa6eea0507f351a89cfc6d16f8fc51997981aea81  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib53bac100fd49f57a5185ff4ad973dfe8eaef6de1937bb32d9246dae9459442b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7ce5fe43a760b5a43815388233952e1bfe5d8b5a7c002f26ae2d462129aad434  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3a2c9aabb8b064f82bd6f6571bdebdd704abb7526f4977a7b98613f883fdc62a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I52f4d169be660862052b60924958cc9a0eb99b1454608fc48d47192452f8b390  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iade009d6c5b9e00f5459c53b0c254dda356081e6965366db7b7ac42a992e3ae7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I52dd625c97050874c15b1980a389843c4a7a890d73f6efb003c4324c029772aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11bf8ca77f64484279bd3f36febe1c6869fb79b4585a800449a0e5c683c6aa18  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I255a6c7b69c31d60711a86b1f0da51040ab60c48952002406e028a200a835049  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I24bc395a7644f2a2d7702656737c32662f8c2e8a7e2b2d4c1bca200dcdf49219  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia84166c5479fb08b9d5bafbf3446230d231e77cb1a3034b53477e2f0632ca74a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I544bba815490c8592dda0fd85cb612828256c09ba1431bc2632b74cc9cd2aa29  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7b8225b7ff4972426858a8550dc67a231d85fe94426bf0812906f1aee0e2d097  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3358739f5e55263208e661a339d6b29f188f07ef07e2ee7a63a24011a4f8568f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5eff39d324b6a8910fad41786d651086c622d331987e649ba4b3baae11ca40ce  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a5c4f290852b8c1baa90ae00400045825f13c24b546dc4a7848f91824185f7c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9af65d3592633577409561b2069e30c73196d1a4798cb92f4d2f14db8771895c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie2261f6d4e2c2ce04997cd365593486e02a7d85106b9c3b568ccdfcda7a9c352  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icf0b2747a9e17f2d2672f7a17111c6bf54bed7d8fedcb5260f25fdc4280ae727  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifb6bf654293ed3bacd2a4ffc883b8ca5e4dedea39e338bd1a30b21e8f8df2f62  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0f4ede6017039c42f04051822cfc539cbcacd77427efe92d393ade1c10a46462  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I23e0423ae4012d108a4e6a495814e0e6f920fa6dcab900bb35cba7b95f590c9b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I571233769cc63838bcc3d61e7a5e95805c3f4116c0053dfe86831eafff7c32fe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7fbf7b7f7a1f0155cb188ee4219620cb35a2fcf98d2687cddfa2508273b70154  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f56f225d6fa40e0469f803c2f72ca27e9c45768ad2af9af9ad10e529e249aa0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I634dc6f7c843c6e4c63ce6a21b9cd7a386600d1155c0696988403fc1ab790217  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieedfb1902d1f76f95f5f971b578c2440fa5de47dd78e9dc70c35698f813048cb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I88272c473a90efa576a83d0c277090f5814599e5aa192b878cde74215909c46b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia3e877a9f66cb7582b125e56b7c3f79601eb8e700f54e14f967a4d9df9b5725d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie278ca9a470ffe4ac78bc335aec472b66707cf02bd91256aff2e7c73b5d2c6b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5ef535b2e573d96fd518cbd837132928a2a0c6a25d4eb3c360f1cc0aed89656c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic486b9953b158eae95a2d8914f8144e669e056675946d245c8239bfc249a16ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id89c8a47964d1e4aa4bb9e96a79092cf7fb55eee5808d6323ecbdecf8926adcd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id1e80f29821e7ae727d759f44b21e84843025c938468caf7c8adfba52f1cae43  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7530c712ec14c8fe97d1699177ef642847c5c1ce6185d1eab39b8416b562b454  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I41b365f8c613bf86dc5e2ed41719ec6823046127babf87a083503ebcfd38ae75  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If9bd4d7f3740f15bdf597de00eecf1cbf2e3b4efdbacbbad889c0946a6b34a24  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I31c470f2adda0a23b85c3245646a168f2478bfdff11a434c1455be20db703c64  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9fa9c98579041b6735eb78f7b3727824dd61991c6a6d91a158c6ac65cb20b05d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9fc6fbd6f2f888b9750fa59a966971aa6ba6fe4eee8c8f3ed4c3ea60141a7d23  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8c133563a8b5e359a6a45a7f3b4e939fc84766f9fa09634d18e5d2101d0c0645  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I84238bd7e53e0dd7ba07efd813661c8cd1648b76c44665dfe51fd07dfaa9b249  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6c3a9695a1c1d22809b1378e82cbdbebc1ca78428194df50cce0a69d6a159398  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4d032ff7482be75de7d2b816ddb2bebfa9e896e45fdade2b5f81b35c003a59ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6b4d2a32c92c22b1cfe81ee6620c69af1850621deea406d75f098da0542843e8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0964979ac559942d1da1c41ecb3d9e94c6c7c0da3d16177cf2379db8f37aa65  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I236cce67d0aea9f9c8d5ea3c39cb598d55f734b44ad6e3972e7f6b91d56001fe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iceb8741c9680982b02ba9fa2dd76d3b45155ca5f688b70c41d66f3b3690dce42  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iac9f4a2fa823ae63e73b655020376580991cd4b2b3123204a757afeefe35a10f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifb57457918458a6aa9c5df68dbb83243fbc49b3b7037575f43749dfe1bef373a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I91589fd8a2ab91f079bb41631c44926b2c6f83b82448d758d97578c314d0b76c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic20b5a20229313d70c01a5f53e13e96095c1d8695144668e66efdc81efdd8374  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I53e90d4a2bbfaffcf92f2e9fd80c491e61990aa575337df13d24211a558315a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie57b3acbbf1d1593e02ad38bc0e07bb84db2655f9282adb3ac5edc311e882641  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I632095e999af63661b01bfe8bad0078cfc2e74217253d3971230968c235bc526  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a66a98136fb7fe52fd830d869dc53a3855a545aedc1d16927f76bc12e319060  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifea15bb5031583fe42f92f554866179105e46b1eac3c6b691958a998c26ac2da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8b2c2b27add863ad56639a306f803b656ee8f91170e649d29aedc5321181f857  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie3290070e785df28e64ff4df124d14c370c9edb924d5f35b059a6c82e8373f91  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I02ed3128371185efeae1e27046aa378006ec78d7c458dcba137f69c29c4363bc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8dcb7a5498da4a9d3e4a76923e84c88a30ec174503cd435864a066ff0ff464ba  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I94024b61447a332a2c36a75bbf305f3fd80606bfbfcc4ee8c5783e3910e9840b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibcddbd4e851466c5ff49f13244c2478ab6c089e6d8ad294cdfbdc8451ac6a895  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I50ff347e89fb452beb071f112e4a51e074cb3d66bd903552db23c17670286e7b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8b5ee5d271abdbdc518ce02f900da21e858d3e2530585fd859690a1a71502434  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I54e64fd01d9aff7ddfc4babeff6703891da38578bb141d250c4ef5949d818cfb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I448065f71638c5abddd1eba1fcf567566281d5b4b23ec4ff2d2208d32a506fbf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6ed6ee11f6983e96e7ccc4e4be6ed8c4ed166ca9075b9cd218f26f018ad2140f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0678dba3dc1a3400ab26e223257bf71c03f0e8d284810653b5e507fe964427f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If34d8ceb2732716c923a7f250495970948ae431d5f1e0a025618c1070940ec39  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I60014273d45dd5019a1b82bdc0a65e44d9a16368d996c8c9ff312fe27e236171  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If16869134ec7e59b567e29a1125f0d27eff7a3c612240e25462e2ee84a7e0104  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8d95c0be0c84d3ee590f8e77065a6ef224e0a75b50aeadea980f9ef4b8d25001  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I28940d6e8fc5937055f8f50c0d65ac9fd892bdc9f0f2a571808f930c8ad21717  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifbf3cda7e0639ad343a64c5b3d2f45017f1d280bf72c96520cbf272104c90ad9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4aabce2cc01e829bb9c3d6a984cf2b5bf9230cf3913db788c47a932ddf71b869  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic9dc8459f6cd65f223a6386c82f754469ef74fbab59ded4fd1370fb69136c847  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib22de4dadb6e63ea49c52cd8bc86dadfd7b73a002dd8e726a9cf1b7b299a8c46  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id6c8c2ebab66fb903f108466c8d15060ed1328fe9a979858569c39069bf050c7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I385f4177f3a22b6fa4a6352d164c7d54c94b980806080c51d00a65f030966110  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibcf016cc83d0fcc2c731aa53147c199b32b3dc7a9f1a255e1a0e31615077205f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7e7be31550be1cacb2acdb27d5120769dd7a0a49efb833051ceb83c8cf691e21  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I26d08096b43367ba37b8f6dcd919bf4ecb9c660a39f2c0ae29f655e42b88887a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c200a5ade27683d4afd55e06371f9880a7bb99259e2ccda5c368fe46bb385bd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I92d28f6c97dab90de260df37f619e0a9000db48e278327a5c5d1528a34bb6dd2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib053c04dd4e330e6784846706317bb6c8b12f9b36a57ee12807bff7de8ba7f0c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0f71479f871309f1717e7a1a2372ebfff4623c315cc31914588df3896740a074  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If49d6a59c1d539e369406ee4e8a2ebb30199f46c335584e62921f98fd811001d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I051f072f564eefd657cb4d59c1c851b56df2e70861d875f3b4c9b95e8945db08  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifc8302f040679d23faab1ed8387a8a3aec85aba86ba9a78d3ca903126266af4e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2747ce9b7349ed89e3265df62bb0d0e612706d8c1b61e30a2878094662da8ff1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3619e836fee4be75d6700a0e72e84df3a5a61003227363b8c4d348b8353075e0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id658b37d70ac8e3a324133f475a77c7948231571aa66ea0dd11b6460fca011a3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I737ae96fe290087c8ae686b90b2ac94df2185f7ad8b4252a6ec850278ba5ea9d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I18777be7a1745485d18289e0b4a6e43e8a2e6758be0967b8cea04a3b0faf973f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c30d2957a73fc51bb7044b869e28e0a8f6e0378a6098ee5e244efb43ab6a690  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I69f7964c2f630ef03f49c2a6cac12420e0998397470245e6afaed2546b33775c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6f63c71eab6c2d7e3eb41fd78c9e18d6362d2dd4100c72b43d3e4b9d06663165  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I23c91b29deaa2df1f4d96e343f6fb852a2b594937a4f62dc4be1fcbe0347c439  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8411087f9f6fa41d454a74dc89e5152e5e8edfa501c8753bd0735cec3789f14b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I119a98150511650722429eab31b5785e99128641bad59a3cb31e42158a648c48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I28a2b1ada19dc69ebe4949a75633b2f543159d2d1cc169f3bb6070c1419878e0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibbbf3f4aa7f74c37a0e8ac8a675ac9a9fec748ac720e6a78e9cf937dd089b8e3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I59a4b1b33d114a1b5bdd708e1f856f4bf729c6b86a4064967ca1faf779189164  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9b13cfb3566db96edc7c018b88f158faa57e4db029e3982290989c6fc08163b2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8a1ba53134dcd1141a6f03dbed0f18ff7be9728dd9a6d6b138ff266c5307ba24  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifd2ca31ff3eec501f34892055a36979681d27574ed8007e4df5cc0109b71bd89  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6b2620e847ea73b8618ac7bdcd8236c4278de3bef0bf1511ee9779306438fa38  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id2cf59876d070e0f34ee834d2691f7fbdb039bc9273329e2ce8eddfe736f0a45  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iae213c2ac7729f8efe23deca256bf56f030403ef6ac00a3bc181414b6a3aa75e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I08e50de7e2aae48cc03a9959d08cab30d3c1c2ba8c4ef0799645787b0c09473c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibf22dd3f14f19c3fc769966f72e8ec980dc79c2991f69d03ca2defb7f720f880  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibdd37577b403da9aa72ec3f4707379b1151c0b15edbfc4fd304c4e35c1672da6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8e23f89e84e219d5351bdfd4aab58f61c1cb310cc731164c6e0dd2eac37b07af  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3baaba73f51f47e6a3f2310f692de9f7b9a871c65605e14d204d6965153ff4f0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I82d316ed1475017844ea73f32085b755d17c9fdafd8191df2e363496e1950869  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id9e3ea08b52843b4a9426b735967bd4ac3d49bd67ab8fc85688b0f55e6df186a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I77e34c24ea46e99b6bfc0f960d428d6ba3ea4f9261d5a183d83c386f259ab431  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I930ad334ce972f0b5dbddf698f6101a196d8072e90d8144b31ce3f4b48a73e59  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4c0096e7bbf30db97520f824e05dbc28e6d1db344202349993fc68cbc95d6585  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I75c796f56576dfba821e867b0de1a871ef35851371c3aa422532bd287f02ee11  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieee1d2436dbda6f58f19df70b691a4ff28d37db8ccc12e04413e45f80d7124e0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I65b0824920910c82c7d677c2dcf4216e86940b3edc0b3da85d8f65505f58ad48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I169d92aaa7eb4f8516e38745955b91d8f6e0ff43cb212186293bb78884282978  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I492e47d35231729b266a9f31aba61a3ac2c93a9786a20f6a152d342cd1d0b911  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2624a2d841eeb09774127e5d709364f803826266b46f0fc3122fcdcf0aa129e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6414b3aff6031e10856953f6b15ffdb0971aeb680d784a7199386be15624ff6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf94ae58c1d9c9206d02651cd03cf2e02bba505f76b849158530a38382396ffa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0a40c2a77389cda4a8333aeaecf37a2595fbda87854a43162ad1299544bd9e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If692b993dc571ec401ce86f38a18ea4f96a797b00c04699ce83ce875b7c31730  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id5a74d0be90678a7b69691c10e4ab75b47914e213e67eae2f20d4b58e8a8d9ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I47b54f01ac82a9eb80a681633a06c4e1d432d358091e9d079f74484f40ab3e09  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6201d3c2d85bffa03f368b5862fba1b2e0ce3735fcc8711cb8107adf16ccdeb9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifcc25cd8dc442c6720ac0f764b432530aa63681953d8ba16b441892ff5966bfa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I256cb35fd6d4e6c6e1c1a9b42dcbc307f858e5f9525acee9fa7af42c820664f2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I67183da8c2763243a285b7cd41d838337f98eb6e59feaaa0a9150bcd6c29877b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I730fa6d01ade8f1439b29b955c5cff62700a90e523a4f4208ca2f9978e59afcd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I37084afdf6695d3b8fb0530643c8b03deb2499f4f68ead04e3b5b79aa4467f73  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee510842ece3717ba6eefc3ccd844e97a9718788683d4c7ceaefa6ca0030585b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I53d3de58d6308b770e4a8884447a5f0b92931c8d83c62c86714b6e539b498894  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e8142c7ece070c02ed90211fbeb423bc2a4ab19fae011793be99c68ff103705  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I425913b12fc3c865d95f1caead00d8c49de08765b634aa444243f4a03a53d0df  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibe0fac26b5e106fc1753aeb842e8a04067fc91c95e358b1caa58db8192381837  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibadfd4f0852067e83ba6f0d57699585ae20eb542d1ad8f2cce3bda0d043ff2e0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ife27bd449bf6acad3f06d6e337bfc29c612ba6b3f06927e6f9699ab24d1e836e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie130bec82505842b184f5dd86865ab095110bc65e59662767e152f427dd7462c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2abc1178fa35959d8eb41342a7d7289e29054439c7bc06adc61f3a1d2e55bd6f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id27dfca888552262f492b81fd23b881938f66eb15f7ab21afb210fc6056fa09f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia96c921ce4e0590c903d02dc69790c6af52898da90f4766121fa7b31e0ce6190  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idf239af48228dc01198fdd7240b8282cf247cbc6969403dd994aeac0e5f81898  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6687de5f8cb258492154a67fd3a3d5ee88d97a4db1c6c273ad158d5205ae3b48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib924c4eaf872874debc3b6ee65921f0381331e1421cbfc3bd17e8caf273049cb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If53d34fa90e564a24f6e116baa8a7934ec4c51c5f0bce8160f0f389391792fe9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If0fe01f34db565bf669e2df82579abb4d3629e8bb001bbf874b9b76f8f780a37  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I61f7e06790f5516eba113bb79388fb515faa1b3a3bf06598a07f534ce2845618  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id6b81456b5d3050b4e1fe80ccc8f992cf56eb0f08a1d29ec1e7cabe1baeb0872  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaa0b6d0f2fe24db548975f410ac5b79f687b7646169247f3891ce9e4644ee0fa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I45ade5cafdcd254cc640ea8725da6961717fd6c50f747242aab6976ace4e8f10  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie2e727d2073eda2be7642a6a2937cd3c4e553d8bb6ec56d914231b5bfb12405b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1aadd9b378df1ab58a1b1af097539d1407636833d9c2d8b08c8f70be326fe199  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If83264f9ff9f7b77429559aff8b14fce54040210c6ba3476b77824c28b95bea9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1cf0e3016bbd2d8e5debffedb198273a2d019ce75f2f8352a285d17264d262f0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If9628510f239b2275efec7ce187b8eb7360beb042a425934ac81632815361368  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7d0cbdb63988e88f9f3f69b35029cb2078b97b6cc9008644b2721eda7fb6cfad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iea2bd90043dd35ae24830a90ed10d12869de66637ab0237a1ad459fa916b57af  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0f54db0f4bdec3ff62a8f1b5f4974982e3600a906dcfc79789fb9fac058c353c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9a4f77c8ba9a40c1b543070a42451ed37c0f22850a4734cdda393e69c7b54733  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icdea1f407aaefacb918babc28247d540a8a52d513d26d7fbb5e81a41797e7555  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I83ec3e2a8ec621acd2afe475255e144f2158e1941ec685a346b75fc471b9cb76  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I25600d0eb62c066eda0baba4269851387918088406d117377eb8bcc2e080e426  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If45b8fca9a85788040c10a47569139b44384357512af96ee7bd8cd98d88f8f0f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I926233df0c5e8461173cedabbf49fead4b0ab577d82f2585af3a1fb6e3130e21  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I979c6bc2b8486315e3db6888ef068b88396857d05a62470d4f3c33833cfde130  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If2b1e365b8ee6d4afa8536f5c2f5c80d31e86ab6729b26795614d75a6a18ef42  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I50e7a3df23a8147b9a87cb5e38d44bce7613b2a717d1e3a8bda1171f9522997f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3d6bb14416567aa7b8883b3d1778b55c251a22ed42b09bb3cbae6a5210cf11f0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I54b0a17c9919d856bb3ed7cbbd8e42fd4ffa33ce8c32d45e4be1e28b71426ee5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a6a17ada186c2bb60e521443c0a5a0248d03242c4ae01b751fcce4abe853065  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I33d759e40b55a0d83119f5c19cf87e6e3181c7e3eed94eec60fb52f9c376addd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I84920b6036437109dbc48865b69f249d82da5c7288a7eb7744ea7ea567e03657  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I78f0dcc6533ef218ce6959768639c983d2119dd518e988eb3dcd6f0b4de98c82  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If64a23ad02d1da21fe63cb33f95d37c576739eb181b0fe50d7a5101817b4ede9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id4cd4fdc9fdb1198c2894543e212f665c925298f1c92b4da9c432eca9442963d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2e15c5739b990462c8a17b590fb7d60ac9c7e6648b79e75697139f55221fbcc5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I294ca1e2c287bbe18783f7043149078d4fcc1c59e24792d75655fb29a36e33d4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ideae854591637828f033505e4fc9dee34d82369d02f7680ef6887c597ac1ac82  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I597d0e1b64b5d47502804c7ba47fd0c17322bfdbd4d332b11f9742713f76855f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icad68e9babee274d9a5b79cf432d9e2a1938e06f51aeb564af6936972b3f8e54  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I15b5266ec781a5ae11540d23bf8b1a0b2eb45d94ab6f367a872885ff3207d5a9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5c1a09aa19ef4bb254881dd92543acf840270aa36ad4e0f5f63a6182a4c93a1d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9afcfde9391d485e865b08f9b8ff69cc2ecaace5f5e26e27b7e1775b625722c0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibe932d914d189b275138de8d6f3ffb914940d4b2bbecb574fba3c6aed885c44e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie2abebb2c2604e435cea102275e0726254ad91df1973aece477e1e5315f82d0b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8befad7180232073f2f7db5a3f546a5a1af79b21cc9cb00a13e266db4eebba48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3a9293b8f323c7e097a099fa6beb33ca299723796aec9396365d43334eb55e35  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I52698fa0d5291f0dc20fb5f24c33e968ea63f47765bb7d231720330b624b2fae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id8d0e36ce1faa76feb8cbe0331f2179ddfc066b70e93e990b5d5bce17f505440  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaef8ec1714d2faf3d3b947db31b7975161077ca31fee04842efc1f7159104d30  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id8da43222903044cc48243a7bcce7864e66d151673396879258ee4af7008a706  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8eb86c8d64d83d4ac46667af42b6383e4d165459475ec6be9d547a70ef0248af  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaf205cfa67ea9b2c39d6705da465f081eb75c326c1d80e63e1331a098ca9a4ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I16ffb13aa3dfd9da5da39d9b2246d5ab46fd0fdb7c02781abf4d8bd754bbbdf3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9a15ed1b2fa413056071c97b4f003717902f38d29805752222c45cbb2cf58109  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a10084ceb62d383dbc5871a208fc087b23de418b2c780813ae950bf4e594c96  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I63f5ecb10fc3ed9bd8bf79403afed8ab1a70600ceb1e755de0d44af98495ea88  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I377aa224e1817d2ab5cb02a5a290a723621782607fcd59b319d8cec1b092bc1b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib1310cd21337a1faa061ffd12a2670171f582e03471ab315b90de9f8fc30959a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iabc9fc6e9581216af19559d8e709ea0842cba4f29f3fdfb05bd71d6d9f7594ae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id165331f616d7e8f347cbe46daff955009fef6f8c0310c64c01dd35990231279  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If17c7df712b5dd40132ac60628bd514bc70092122a0cb89ba7d4559439779fc9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9d7506b5ed3de0e32e821ce6ddd1c28aed177910ccacc4d4aa2a8ee57212d162  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I734136c95a40c62745d684fc7e8cd1114b883c6209df11cfe01b9174cffc720a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibae97ff31fce14dd0506fdfe7407fd6260f7cf8584a01da77312b1aa48594be0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iea011619fa5b0fb7d22dc4bb4ce3fcc4856dfc7286ff393fb329ac0d7e348207  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I954e0367a6f3af96a7e033da51e7256543d7eabd37191d4b03f3077567cb629f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e6d7d9769dc32e1e014951538f1cd1014e9d07b675e6369e88ad5a6fd400787  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iac4172f940fcbc93db2047b26fece588f3fa63ef255ef404beb5e6ea016b2ba3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0e9a7c6c53b89ca2685615c270e8ef3d3f51fad8619953972e1037edfe633834  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib99b447a19aa10415461faaa8d8026b0073582bd078930f2cdf0f531259d9c50  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icd30277c9d839d833f27f571231dd138497796d3e7818460d836a48b87e34d03  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2862bdd9be64c24d98e80e8b662a7c97c70943bab3d49cc8d39443abcd5c2c3c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f73c51d25db7485bf4a0d63f95f14fc0661431870ce704f70cbb787eb336f09  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2647390c3800518f2251794a7ee4aa2d71ca9589534cf73eda0accbd2b3342da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie05c1da46b594d3c94aac179f6c98334d0d667cea08108719b44541b7b0a2049  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1bfa3da571b0e3d943ec7b9a8c641283e080bcc6502fa8317ced3c0a6eb2c4cf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idfa7c6c8248be1a2f8a95c6c74a71be3126e039a31f4e16e0b964476c6d47953  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5c43417b1bd96dfedeb36f6d3405fc7f6b73c11a55f21ebe6ffd675e991a13c3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71f31c9a9943d9fd422d00aa01888aac32dd8b34236bdd9bdf3e660413a3512a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icc43ea934f0c07465170977b52d2f402fe155ef77f3ca27119fa665a1d918694  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I78abc91706fec0893eee10a69916f7247b718169155038bdc0bb6f8661ed1c3a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia428f915c49f84567006696ba3f5c783035325755b4fefcf74d65aaae1f3d3c9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If270910122bcee1c18cc592dba9b38c026f792d8d1472400a09edee9d7633e22  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1517acf28729695d689aced1c7eb358d9acfc4453fedf95a76fc22c972550c63  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8ca8dfb7a3a8ecb9eac34d1d1ef4768d31b86a757cb7b9ce61ef159816ceea7f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2cb1ae23e53b89ca0fd3d1df98b32d5b9e478e9eb579b0875981a6b056e8ef4e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1a2646b8251f83855c3fe8f6172f36500201ce43b9b5ba2cf0f25fd5d540e89c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1d9a8ff2514f112838c7e4f568303dfcac3f86d94003ec4f1a40a35b79ee8ef6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I83c8ad082be8fe1a71adac4f41a3bd7019d2df299d19f8e5a293367e49b04fa5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idc29625b375c44e890e371217aaa25d5fda337ba8177fcceca881adc72292a3b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6e88f83ef5bc5f950a4bcb904ffede2603201e72e362aedb8db04412f7bc2bd5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7ff25e517e328eda581e7637a2114a7cffe873df520114410c0487e503c01aa6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I463662fa980f8a5e4be086aa5f37db53b1d6ea8dfe11725b8c407f779a168998  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8db02445666e4aa12d7e495ba28ca0eae6ef411094d30330e91eb9eb03b38aa7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8c971b4c1be575fe328c0a4a9ecc5dc75f08d36f65aa58642976d971a6c316d7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I09e6d011dacfba2800f9ade6a495076a67e4acc6a944fd649a7c382422e8fa6a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I76599c709cdbb3f3cfe4071b96fb7dcdf8e072fe85ad5c8e7bbabd4f6182303a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0d9bc57dbbebd429ee5a5e5dabc1cd0bd9f4de95a920346b9e61cee83969ba0f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I91716015389a9d3b1d0cc77327f439e02e54be0d3524b2cdbeed886eea673b10  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibc3e77c4d6cb28599b7a21c7992802beffb168f54d8dfa650750ffdc6730df29  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I34f861f0a748b0ad1550db8ce40149dc638194b0089cf22e2380a39a49f8c902  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibadbb4e272ab1105914763e2790898c8e37a553a1b6726e8818431bf5209b369  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I308f551a8479d066b2a4b473206e8f407082cf83b37a376e6b0e1454f7ea2635  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I58c6fbcd5f77398c3514e6a850bb69d9f57880a387f10132aa63079c0a1f4857  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia9d25b6cb880b9a00c9bb27bdb80c08988eee46afccbd578659eb98301fbb8a8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ied710d5ba03554d4103468029a9d895c25c10765b6e3d73bbdebc54d7cc7d8db  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id7dcf87d2a40e82e7f01327d834d5207ae5873a7e5133c3dddead9d0cb9703f9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I982c94b61dff8249f2f3055f60da6e2c2b0b56c403f151168b28a5a211aa6428  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I710a57e6c5c8e228325430ba2a5fc32ed9da101d76ccf1d8c9f3397859b39ef3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2cb87b14b006ce6a36ee5439eb18a4287c5b9ae79748faee259c0435d0dac81c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ife00518e7b24a5de694b56a32211898b3c23d2dbd2df91a4197216c23fb5aa7b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ica9ef16b19711ccdfe32e34eed347b590635f1ba7983272eb02f980f80642254  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9331a9d6610ae5cb77aa3d477fce0c0ad7378a884c86c4872a1573f2d8a90d8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I48d9ec419ebe83e2a5a8281e7beac36acc9e554b86b154736dc51ff940f5348d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iab97067540ba8c9551711cdbff0c6aa3993534d3e8b352bda090a0997c681afa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I25c667a6616c9a94f6618166c99298b28d897f9ac8276bb85816e4b42582cdfe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2d2137ac29a7c23160dedc43e9caf010f72f7d08b057e49fcac89984e616fa5a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11775c069ab4acd951a3ca47bfa65c7632a6a8a369bb103d0bb719806dfe0c57  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6e418efd4b385b2a298c1c53d344e35f593e8380d1c27d7cb62cfe35223121c8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifd66abca1532f04fc777617d91cd2d5f4d4fee35c3f075e91639a196780168d8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6dcc482b16866339b78b922f9a7ec0f4a0ef311c353e6a4e107dfcc351abbb23  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8c8bc477ddc4000dde6459d7cbc4ba665fd4ecd97242d9f9fe97ca6825bb033b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I54da11ab334a3942047eb5953935aedd00ef1a24bb5361fba51504632ae61831  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide2ca364c5742f786e5408980fbe12322ebcc2920fd99ed322112d3623d9e372  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6024b75d70e3da7df4e532e712df56a8bed06352ba0a545ec355f59473929d41  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia79355adc994f77e150b93a3e38c8bd6f0a5848a212ac64559cf1210ee0d11d7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1b68e82cfc8606d3a9325ff2da047f345e2f34b44eb428bf2a3bdcf42a6e869e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia1d4bd5d90332afbfaaac3cd0d8f5fcbc626ec4adbb0b0f16fc80923925f703f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I87af49f5f04df14686aef62aa27c16723af3ad05398f00e29788666b27784de5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic1211f3a0703e281ce073a20afbabe9b2a698d1cf74f07f099d21fd89ffc8908  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2985f4f17b726f40ab6609b57a796727fe46605944c5e25c594caa8dfbea9f58  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6f7aa66db409365eac05a200d0a0f1d2b25e9c37ba4a7db3b58a7298af0fd6e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib1e319af12dcd98c09841e8b06e7af86f2569bd7afeb1718bbbd26e30f65c464  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I30e28a0e32497e3137bb689fdbde46389bc490300e15be88612f28eff07976e6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0b525cae7fe005cf25a07cb0b1486152d726fc74aa55f03480f10af97379953b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3df4fc0f2f099890a34d7b376328da6460d429e2516a5f8fd1aee5a8fee835df  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib1b15c9e15e963cc4f2e9caa1b6b132e338947224b705b51ebe710d7e0f661d7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id364040d3b9f1ebf34ae3fdf7465d955b49d7a2f4709219f76229766d6df98a4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7cd9dadb64725f4217f1330c893724a7537a616ef41d9dc49fd2794125e0dc3d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibdd77bf8b31352e365f7e6440a57247a8ba62e667b000c1347165bb39f3c7c2b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I35e7fd3f09acca79a1003b0a4b7ac62c4a2be93bcf333abbfb13a5eefd7d5eaf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7e269b2e2d9ec70c47570bad75bce0ddf53e85e3cb4ba87f784ca520c5ff1084  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0c23517b9814053cd1f89a8b80a64fcff6ae65937dc97199c0b79ba8f7a34ff3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I73ecf8ab6430c6343bf7596e671ce01a3e3e7499813ed75c583a7103147b0bb7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib7f659da098e577e33fc0f5da1c03f6d3e68b3883ad7888152d2e8684a6177f3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3386ee46348e8c4359b1ea2153bc64afbe76f2b6bc9a312629b8c52762a22873  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8c2fe0c8cb55f09e4dcdbaa3960acfd815764161f53c6234273dffe4558644cf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idc64cee034c1ee132335ae593844b2c46e3f1b1b2cda8699940df311735a32a0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c7699448a10638886eaa021495d4c7cc378fe1e9b0aafccda001c15484b9419  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I45b03b0185f9efbc11c707a64fda9203cc82ec2fbaee7ff34610c74d7cc1132b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3097f16921e899a99f2a2b013a3f6d339ac9672fa5e17655ceba4de2d506e151  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If0d62663c8a08719b83a27c76fa62525eb14d452d4ff0f33e94c67f58d7c86f9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifedfb1db4b16b86149f5eb8b0adf06499331d423c368c0077c738a190a1814f0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ice24cd0bd76a7d12a0199df195b34f41f7f72f037177656693b3154d102ba729  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6148a04ce3733485aeb6c4d20b6117eea37a510aba76ac29e82d44980bec0934  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6391e6b0ad4d9fe4136b90a57d121f2b5f16ed4662429f1b85677591fee37a6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5dfc39b913b8e0d00491e3f7f45b6b467a517b5e87baa065097e28e6d695500a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie538f6d2c778992e2324a9adbde215acaf7b8dc3a72a9230d4fba2332f3cab67  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I03929e638a59a35fc0168772ca06f7a502352e03525042ce6d49cf9ecb671093  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieb5e001b45961175497657da7a0340c2a15b6d8de1b72ad68ac3aa7f96a47af0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6d58dbbb9b18e4b347b34e548c70a9bc0d819986fb3a6bcc3ff8a67c1fce9c9f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I82772b528a8c156f2932a23a720f8446f3062e9605839897b4652bb2936fca1d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idb259e613b71ccde839570ff2e7f21a9cb7bf676ffd4aadfb08d6a963bea9640  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie9b1b4412060f1e9acccc1f3ff897bce33f24fea3bfc91266f9e42c1f38aaaad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I259a9b6041f341013e6ea0706c4e9ef9a77148bc003b3f0cf9593ebd915b30c1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I41a57b30ab1dd9c40a723f99315558a47412465aa3fe967250572e8373aa7180  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I42968c25ee2870f891f69991ae3ad8bc1c3acde2f8f4d6c0cacc48f562399c37  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I44103a07ffcd818c0d9280b96ba08c32f96edc83a981ec9748ed3d6e9c061d62  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c886223618a03ba9e18de68462ddcc522338cd26d24b5e126da9da1df1339f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iac242fc0dcf37a86cc334319d77aaae46dd223017f2a6489c4e33314eabc9874  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3225ba7b6d0e0c7a94dfbc8e074ade02b79a66f6aaf97580a451c2d1781a625c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I25779b63a47c05d4588d4b33fecaff61647609a62fcc90f0f541c6b30ea9342c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I05bd9a1d7818f4945ddc448149dee571e80dca8b6eba7ab79b17b6f84d3f35f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I17eff5960d8d41f0832a48fe9a3ae0dfeef1bfc44b73eff506fe1d3813398d15  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1b02edd5d00090446500b1dbf66a7e674de978c068b81ff0b0fb7abb9ffb1654  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c865426b0f044469b391bbc13f977fdd19dc89c908574ba289388e382d55cbc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2e557a901de23b8442e8002b3560bbf9cb8592b7bfb7a6e2f8aad12843a5a041  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I469f4965961eacfe3dd0cb82fce4905e19e6695d71bec95956e8209d2ae39ba1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6e148041c3612c795f1eb1513a9eba29e0509f02f94971fed189dd9f03d54a4c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2f687e6270528a72aa2f9f9cc0a5a6368f8eef358270329cc40b56abc0e4a35e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I661bc8acd80497efe43e3d6fd92bc4107b1ca63eaf162cff5695b35f8d4a7e26  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic72f2f8a61b8ecf8960d476bcf8fbbfd4389e932377679286e7182cc12c418c8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I823e337e6437e5ba36ecaf0b1ac6b7a4e74cd2ed7019dd5447355626a8877d89  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1622b11941b00f6d2ecd90320158533a66501a6ddb78defb4464a937f132c232  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9ab473d34fac3327f03768e14c7bb20056aa8a3dd31520d385552eb6d214f890  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iedf1b21de2a0eb04c4a64f9eb34e2b0b3a152d90b1938b61ca45c880eab16ab6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibe3e6de02f0c30287dd89b07be5254ff70d9683389574d02f1423e792bd2d534  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iad8ee4f6cd13a9f415cd3519de0179a66cfc993a840b3101cee554b55c0e7e7a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I15123100f4377e14c62cf47fb1fb652badc3bd0e8f0ab4b970a0bece065a6380  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic0a892c18037ef674c8d94cdfc94cfca47d977ca2da9e678303255b96575f022  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c316e8b8cb6b499a7a8fbb513b3067829197cfacee877c35874a2ec686ada4a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib3a2af9bef5f5d8d7228a3b49a5e0d4a37a33117e057078a552588a24d46addc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia042bc20eb6866de0ab9ca9154f0db63f7d4ad84d553be858a0be88fbb8f7f33  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5b4ba308b0fc2946fb11b66aa5c24c7b5cb2a21955116b97f3790de65cd2a064  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I005ecc3a38317079c7bc5008817e11017c33671f77364ad9a07d0eff1e0ebf0b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib63856036797d30e60f13453da509ace15e3324c25bdfdea5aa495d592e2006a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia9bf10fecfe62530ea6be4687ecf78a2ac08c6fc6e38328c2d64a80cb5a3d72b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie1447c9e1eb4ed110e6b0353bc5dd2cd14ec645355c3cf897df6f6c5808475ad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic8f640e7a0c71ddb20a985259b5e48746d28d2898383765c3b78c577f281d27f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3b1d695a626aefa8e5b146c7f7f26a8da119680783da7afb019209ac9fd719aa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1d91c7e9c2f99df4e0523b7e01b6fa6ea3930382238ccfbc07201b7d3edcc969  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7c1e9623dc53c8aa8611b46c0375994510a97c4d49d0b091964cbe4671acf1d6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1b5d096081c0190c0ce6a674de1afee9ccd766a9cfab0637a0aec33199061bbf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If145a331c8a8abde8c26d2571cc8b38e1eaf2768a4658d350cb602bf8614a521  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I86e764dc3320206d9b52013c2d735ff4d27bf6e4a82227486e64b4ceb68dfe8a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4a98524c02346f4b9468666ffaa9d996b9b868a5a8730264d798d7a66b7454bc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1187dbcc72f33b4cc3442982af526be4cfca1b5ac65be943d4ec380421632117  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I73ce2860dd9aa9ca2c0d541a6ae1e5069badd35988d922cffb6aef0038cde662  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iea2dd4d33966d53ae739a16876ac2cf04e1d95374a5af68e59a5703dfef2aa79  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic0a386f5301913434a3d6aaea1d56d6acb3484fababb7b8831d09563bd8842cb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia8a4fca33add1c3c58b04eafe9d023751882f409c5d2905f77aae3fef8c2b008  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9cd4ac82c1e6f2dab27efa85314df34a40d8747959eba18330bd424a38debece  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9bcd5f3f4630ce7a24ea4479c9ddfce59ed809dfaad9d767e80295c41b332f4a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iac7a05e270cb898af4ba32c16445d0dbdffdafdcc5fae209f09367abcff9d6b7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iad7f008b5f08f3ba94a0832261fb4add17f0897e3c7d54a250377b813e284331  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic072a2fb2ce65ca734c05e747f12ad094cc5aaf9267dd94dba345b5c7b11dcdc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic20328b806ccf89387180fe6d88ba762051c6bc2c7f82494129e8c3600108804  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11855780f53e8711f8eca9370af31f472dffd126c02cfce8154a959f33c68af6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I39b8420e976cbdf011232d83446a5cb92c2ba58577792c9c61dd71358205e936  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibca01267ba9d7e2fe9f8df34a548836390ba12b9b782f16ba40965c00735213a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I105a7d84244a0d9143b9b2a3c64ea6964f7e1f43b7f8f5cb15d579885bbf746f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1b0f11f3bca53713a53e2ed18fb81f5a25c7151c874be612677f5204bca28093  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I434991f7c09dac3a7bd42fce3073dcbcf8b1c6579822074548ea94fdf1ef4eaa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7fec897140c79264b7b7b7f3ae228ed090ff69351985c07d317ff9c0cab1e58c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I82bc7aad8e3adf5b7bd03d9fdac6eea60cb800e4502e3af7bdc9d49139563fd0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I218ab164221d559f1e8bc2a13f06a7593eb4133134762698eec270be5d4c3906  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4135dbaf658fb73b41800cd275824d1c9f410ab1b6e555b6c4c8df12f96c5861  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ief38674752576e92e90fbe2a7abcfc952274123875a95657dd42c910133cccde  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I783b89f0c1e5463646e0fceb976f2b27aac523a677eff6e597e434672b0daac1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib0ee967a174d7c841ebe71e144d6303bfc80a6083ff6ad745c76d488dea66d9e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iea7b69c43ca4b3707d3bfddf19b27616b8686df915734ba86d3685127bfbf39a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id36acaa2c9161668c95e2cc3e6e852e9243ca7f486ca6c2ae4d124b1a8ddb522  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I325ec6d7bab5ccd6e9c4a7e9b02a3b8c30072df123bf6318bd97f1e8766457c8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I07c37e958136be68b3d658649964c73ca78160582248da1d45eb9ee82c1f679b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie17e17c22c7215d0482ba310638db13a96c0943216f9ebaf53c0c29c69971b23  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie44aa17133d02266160c8fd6f75716f8bc4a3775356cd1ef0f495b13145ba864  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idaf1699bc7916d99a2a5ce0174383c189dca6d7537734b19dc379bd634d0d209  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I64aaf806ebf0ead2a4836251dccd62a394b984823592340be94f4ea02e12d766  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I152b3a1e710e5a39bac6338591c6597ee2a38fc25555f563beb7a1a967bf4e94  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9ede22dbb56f48c045a1b5a05945124fb97b6ca7e355dd8d9dcfdef6e623b953  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I30e30c2bee3bac86dd68fe8364f818ab63e91d65c4fa1ef45fcfd03c9df87cc5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic0bef9008769fe36d726cf80506004d66e7c843a046653201c9bc2c816115c28  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I252a77c3eaec2d6accaee6de3ba5d0b354636e2a2aef4992eca0e2a74eb4d25f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5fa628cdc28fdeb96014a4d2c2d06b092136cf2a14a0420bd5d3861b83687413  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If258ff7e66143201e30b3fd451e1b8e2ec9e46596c2653ec836617c093f28018  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id160a3b60a3c7a3ad93044461ade9ccf0b7a627efa4b1bba84a2ea0d4fbdb551  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia42e25bf722566321268c83de181d196619f062381c7fdb381ab5f6aeba6589b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f96b4022f127e7d965786f2cac8ee6afdbee96980608c876c6b699495f80b0f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a2505f0de03f3e2d303fd207ee819f5a1777b650930b87a235ab3cca5de6e87  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8600d4c5861319be0efba19d9b66ad483aa7bf648f2132c1a339157c43920c18  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic551d228c593c4304b4ef79a965ac1d9081774282af09d79cd587ef9abcd6003  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I01d7d3d20ba0eab63d519ae054b6c22c5be4000c846a6a4883ffbbddee37663e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4177cb2b0a83442a271f59bf4f758851d5146ee00d76a1177c9a34d4208b7c09  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5df828301af902c72794032c0e55d8e7548c9b2277b2edc77f53796ff8e04804  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id595e96924941a80a6ade8778fcbcef39b07a62fa1d7350fe50182fdae302556  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iefbb3d08b0b2fc51d2f6b60b25b8143f3f88a705e770396e2f6d050632ded97e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71c3a88492c33461f93d43680f11eae8ef3e9402a4b931c5d31f959a2f8c147e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7a7bbb1d7d9b77199c0b29fda08f8a63112052ffb0a502a05586ced336e13c62  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie1657c5216d7c6e743a23819c08b7c7f2fc8a56793e1bc67fa5c5f3b37976641  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icac36c9706c9e063b771faf556f6699e280687be228aebf6ce71f5ae775a9754  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8b3bb7a4701d3ef22c71a9631482e13afc2ff80f40e2f0ae75cb2211af5ce6d9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6a24b9c3ea194d09d619dff007c4c6f53a3cbbbae5c9d3ba718bc3546eaad989  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic7af968d25c444d210ebbc7ae563688f4f8a48f38035ce5bccee100e10555047  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icb61d0767612534695d9de0380a1febbda612604f373afa55f0339c7a679e99e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I58d2fcb7085fddc9250ca075b010afdc2d019c4091f5d115d9520586224a1ae8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4e5dfe1c7112e24769a5e6aa86584c09ed659fa5d05af38d18183db31189a3a7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iff97998b0778cb649d03228ed3acc81c1b3a97f6bc47041c423120b1311112d0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I422fb05bbac12ca5df13eb7c0c3fd96a4e819de9669ccd64d40060b5db3f3421  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I782d29ca9e53ffe86cec8809d7d413c9c5ebd9edb6a0d76db2d0c321312d224a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0705e6f1954b14f35dd7fa8a64370c2f9e6e39b6e265857e72946815d1f994fe  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3f9e2f1be98a5d14a8b79b252e9b5a2b3a09304f27a3526a4a66b365b682787c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I134dfd9d579ba8b2d72bf1c47119a086fcfb6b7d591cc2c5558e451f57636d0c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5f4870fc880aac0f84130a26e3cd493954ea49eb3804dd17a91b2ba1cea599f3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I918037e81d2f9c05c6a8b94c64724b1d0ec8afafe5666df433fee3e296171f54  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I136f70cfdde5473f8944efa2b1093ed76f82dd06a341413ee2a56054ebef5fd2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic02dae50f30bea04d63949eadbcf892ce936efc5373a6185668a20311dd59f4f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I54296c97ecd9a699f171f4d7271c761aeea50255010a0a90d2dabc16a0cbef79  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I50a310ea41e0637bf28b5f56cf11560bc936e15c73acee063c60668bfa905fed  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I25d2b0d3ff7f684e508a62271f3d29c729dc46478248627013dd91075f8d2146  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7f9f83601cb61fece60f94c3120b43ca0c737ee36b8c67ccc917d3a428d8750a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If4fa37977e1db59d1bd7a30b2b0919c997b6e25e0438e01b62dc273d10497867  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I66291192ca8d81c8e3f667651d5201cb41b6872f73283d13c6718159b008d8cf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4bfef3f43cb1a77ce8b2bf4b26160a161e7f28308b8d2817e6e2840f09463e37  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0aafab9f9205eb4a8c16e213e116d949a5c625f7cb2b0f3d124deb80aad2c6c7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9095fb177f965807ae5a73a45c76b1c0b6300c6800b17259e5836adea5a78ec8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3780e5266741d9a9435818f002588f4c44ae518b77a30ede57a3823e1e1e5867  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I360ab21cba3dfd419f0ca83f85d9633b918c3d24a00214399b0465d7106466ad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2c061ca6ba4299d676b5c6f1e1cc920bc1104e7ac730d207949b952d1a98300f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ief44fc6df0864dd0766877e0d673847250f53ab137cd9029916ab7149446f9c2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I353e1673347daf260e61fbba813cd14f83c52ce3f6e5168c0fa6308d41e93590  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idf77a6217d51b2439f71afbf5956a52a241f2bf8722f54cb166d83c3b45f6721  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8ea9b55580c15fa584fb934e010debd92e2e893630de456e85036d583921011b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic36cf3da50983e4168cc0a31ec0a86c171714355c0fab18398b8daf57bee1a45  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7469c1791d81d0924eb0faa6303565dc78fe9eb371fa13039ff89b92b7f51a6b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9b8a4dcee9668bb71803c25e0ece0eebbf704eb29cfa7b91c47cf48d61076803  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icf4d3544466d430d71abf2513cfbc16b575af540d369d405ed831753f304673c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0568efb50e0bb85c39c9ac6d2ab3474ab38799257dac5693085eeb0d74859ade  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If072f43c0b06c41c30d9bc40dae674ad9052e5533b1308adb97cff2e03821bab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2f05dd0209278c1e661998552da73728c1521c024a7d26f4652d4f151c6e5f80  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I17dbb17fb2770beac552dafeb238c5e8e7a948c35c7c543508e652cbcda01dee  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I68ed84b705e3c00d0fb66182d6eeb93f43999532d713f81fab39a36259e0e7da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9d1a378e4d5703b65f197cb76a1982cc10e0c17654eabcf10d9df091086d8acd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iba503643311c9dc3366b9bb843dcc1ee2f0243c4cf78004a660fca224b36c5f2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I05806fb5d45e4d6f569c12116644b625b7ba071eb052ab97525f06fca03dd88b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib2630bec8f9f78489ca6cfe0bf25746b720aa422b9d529d67d6dde2d045d9c3c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic57569daaae5eb0e66117615c8c6043b5f76b114b5c34b0df50445f66a22849e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5cbbcfd1cfc35b3e78d01b29831195106ebd9ba5907f44dee6761c2b047c4a60  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6dc5ebe003a649f0e4106dc27f25387651d43259f0ddafad10411795ee48b40c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I238a5c9cd1dcce0d745817081a4b240f74de3de6f18a3abcc42cafbb19a0ad69  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I53c29303c76ac3c1c02fc9a74eaff9595153ba06d67c08e07790c58e53b674f1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia92993e9a66294adf7a4dbe1ea88a9e8be6367da1c05b8df343b3c7a38bfd8b6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I329448311438699d3d590bba6ab4bfc9cead805f96015b77617f42d957bde7d5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I717aab2686adb8a0688009c23d92aa4475e240ec0747735e6fee5e196a50c444  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I13a54b612481fe0fdfe8b52909179bb82298c2bff4f10adc4f41215fa4396311  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I26a27b64a7aafdbcf4a6d058181fb84e0e16767f4bd7a9c45211c4c1246d3b9e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie46448d24890ed6ffa2736abb97331dc3ed219b9324bc0e8453eed6aa2a4806c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8ab86da421b01a03999daa91e41ae95ff58c6bc38566a3deff72633a5ad1cc18  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I20ddfee724da47731a2062b2732598b429c42f7d22bcfb300dc084de362a2bdb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8d8dbd62189397b5e9189ead2126a615d5b6cea393901e21cd89c255d6672615  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie79db7f22cab9cd57482ce0141d83d5c1ff720a7c3dca2c3664feb4a1e2f4850  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idcdcb2dd5e2f2aff0d7b362ddb4ae1ee4db08edc2c3df3589a7143bafeec0bcf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I525b9b85b14df7a6533a7e54bdc9bf40a303c890a4a410251c8d556d38b33125  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I65afc937c55081dabf16dbfd02eb03c97204efbdcfbb523609571bb32d537d5e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I45a11cd2f581121ac03fe112ec78bd07c070673712fe6112a3e4fb4eba298e27  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9342de9fe82f2273da138f99da619acf144edf1f9c33682fe3b1a09d0121c4d1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If6cd81d168d83d5f6a7ca18051bbbcea5c7a9e017cfffcf72f31f73275c3a4d4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie2c7966ff2c1e84a7ae016f31b0f8b9ca7aa42eec03467c7e3dda37dc34f070c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I468b28bee4fe1c0d20fe7abd9338bf844ce0a2e322ed6b6de11e2ac621572c48  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I08c55e08731cbdc9703e607b481a65177e7e1e242fdab9bfb014964bb0d1d22c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6c252caff8f1ab047efc25a950ce3e3ffb47a5b779e37a667c48bc1487528218  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2ade6ee1b52da04fce9491cad314947a07eb9aaa8b0a430db2f96e2d290384dc  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If6e953221a61b86b1fc339b69af853f6ad538b60770f2f7b880d7aa15bd625b3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6c6885b180013a16955ddefa0dc75c25ac85fb76059df9bf8b63af72c8c1fb4d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I907aa3f6584035b934017a601019d35f353b3f99c7573bef60fad167f9d9ffe0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7ae7cc2f052d37b650c0abeccd841b1b18abb4049c976fbdbab72ea579a5d206  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5c0776e9826af1a98810296a7cb86adde5b1b41c434e6040bc6a5a30172d1bf7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia244be7d571a1e41348c37534a23f7cc942b689cbcd5dff8c10043325b80e322  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I14730b2825dc07428388347472491ef3abe06da3bcea9b7dc9c919079c22325c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I22670670d7018cb361ca0ffd92516837302d5528c26915b62d22505471ab7384  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibc34c6979b8f5adc5421ca8603b6dca91161055286758ac10d0c612263077758  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id39c55c4f0df8a0d8ee4f8b47f3de8cebf5343bf75521edfe38a695565eea926  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I06a5cdf2e430e40b5c08ab617356f6b4b0389236041b77e2a57d9d314bfe77f3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I22c3d90c4ad5f41054f9b3dc7ddae143f567182c7fc695c5cd087f126ccdbcf8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I533d6897ed500a803f6f6468e36a2a922495b3effbeb405b47ffb7a5f4d82c89  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib8d3655f6360b2b189b79353d38c9c9989af811109144d45af0f8b68a3276149  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6b264ac5221269381b155a30c051523f4488ecdc6eb2cf60da80a8b84c49bd96  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5c3a945e8bd4c55e9cb38d19100b13668bd652bc1162d16b30f1562a6595a032  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ief691d56b56a000651b0a4c6cc9f26bc44da82f4a6382550d96ea4101b81ecb9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icf55933dce8b9f95a57d7d019c9b29f72e08454428013009cf0e4d2c5b6edf0b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5b0da0701e7399ca2e668c1602f494f41127e4c90e6fa91632da0016e7b395e9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6106f96669a63f337b78a6bad5894881230f0ab6467c23ec877cf27a5bc76cb6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I566a76fd27d46125a614f5e0c72dff06a0c1d836c7fe4a2c4086129386b34dde  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic754ed4f2d29b948b422876f371df4f89b86976e25183ce1b9f664e1a9b19f56  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id7310932ca8964fd49adc052220c04855b028e29fb7a48521a36e2dbe1d6d5f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibae8222f76059e8f61dff938a64e23080eb668880ac50ecbb50de852472a22ad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I09673e64aaf6f35dbf4aae16ffba969d08a800d32ab25413bfcdbd540d7b01f3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3ae1a42457a669272eeff1bc293c80c67239ef6b725a09eacb82b06ec84edd65  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5b4c4554a78c551dd34a93ceb225237a2d2540a0e05311c4595bdaa5a4cb14ea  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If27288056468d3ef3052303952f2e4be67796c40d6224383047d71d996f98cf3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I12dfae8d4c1a0612c6d65c6f5493247af5e06ca1d8c72dc28f9ca41b0bbc6ea3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I295da244d8dab1563a5947230e49171eb905c3758c289526ff6d3e0c3efcebbb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I89cf2ce418b6d96c0e2b9c8e82167a47d40ade45a8f08255a1b849a9df9e6d06  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I47ba4d6ad7b1889cb52ff7a1d42176e166270e39a1d2875f3a0cd260a1fc92ab  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I08240dfbc0f698324c1ffdb8e769016bb8b947fb0b8dbb72839375cdb4cc47e1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia9ea47bb0829c979af002fb7aa0e22072671c2876bcdf79365ff2b3691172149  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I58df4f7ee4282cdb7bb80c9f1d907ff37590b1db22994f3a07b521132ab80087  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iadfdcb3c0764107a2b0deaaf039babe6a08f1018f3718f5539718ed6a5aa962d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia2417744c8f15898d5d951e15cdf8c03d932cdac6acd27e32045e0fbfbfe4f30  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6d70d8c6d44eb58daff53226cbb59eb647b6dec6bed37021a64e16ac5318d484  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ice3b06f04279add8283c8173340c2bfd4b4801d85610179943f070aef508a893  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4fa5ada2d589c7a90e700745aba8e09edcfb0252f532e4c74eb0809c712a36f0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I71c6f88cbabd48d41f42f2b16170c8955b79d20b8a8b211e174d1c1473567ad4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e7e130607ec849c80f9e687f0215ceb767a2650626f20ee44a6fe677fde2299  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4c02563233638e273f05bac3e277c702b38c204fda200dc5ac163662c77a429b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I85d8f259f770b22a380d6eb5ace0281c57f0952506152be05f38482c47334988  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I989259874d3f12b373358db47fed6245f192edac9e7df00531ea7ba75c360d4c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2ef69d9eec4f925b598115d569d2d85a4545871f2ac62635f9b072ba718b595f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If8cefdab8d831c3db83e1ef615ca534f34c58b9903520c7741cafbc84e28d207  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I00e5abb30adb527f6b32257212dc21f9797e9793ebbcc10feae9e524188539d2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9349cba960e03e6068aa27e997993b0c466e040a1ee9e6053536d3346c84214f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I19797110801d39a7970e6d8665215c967071ad9a1bad12c33401b44f595772b7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0d25b3618b50ff21e3f301fe44087368e38fd6b37b6f6fab004824aa9df51f0b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iba62c53d136b455b7d575b868f2ebd2dadc6003981aa2aae72863a0eb812bd1a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6f2e4979fa9229a647a81a4fa3f8b2af809199049d2554ea15fa9a6ba2f90a9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I83d70d4886f48dce0888e203c2c333c76d35f0c73767dd9443ec8fa4790ecb09  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3f92074e96f2c2711248b1d770b4ad718a565a323e6fe4ebb379e6494039af47  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia478acf4034b69d392277c3d5c6683346547ff26d418b3a6c36a3f9a56e3cfe0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I06186aec49594899011a9d7bce163a3a43ec094d7c92033df033594ed5eb43ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icd8ef17fc44642a3c86a1cb62727eb607e3a4e6d0b021406b9b710ea5c96c06f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2a3d1a32b282fd624497621815c6ff85c904f5f3fb50f18cf345c5a5d7a557ef  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibb57ab5a5468d08c8b299ee67b535b83995e94d6223d0c6d93dba8580906e319  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6fdc128e94d85f0f7f884ee1ff44fdb6de2ad5b93d83c3e36ae235afcd3d23c0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2790277776fa84c3edba2332cf538f8ea3a40c1b06cece7463a3b4757b1fe213  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I068f00aade8307d2a2e2ddb37d7429a04c2f6786232134a041e62733cadb03ac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I07087056bd31363bfb1f76f8fbeb18d1deafd5e4816ca1200d362c0797a77bb4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I01c264f9a89aec9dc11fa16206ffee1c8fb03bcb279e9e9f53fea1e94e9d8b23  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie42f89c20abd223240a9f93a89ce650ed2f581e1ceab0587a4fea2ddf9f4f98f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I44ba42cf2460fce5fde6d8a9fba799517336268d29b5817597d819a9eb83df0e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie4fafd34aeca2efbfd3bfd3bf45f73ceea27b613ed242a43666d85f3680ada44  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I65cb4f1288affe61a7cd9981878d8519db25d724cecbb80eb3932ccedafcd5bb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I577e642ba232b9a606abfddc4d84ce4354744e2f953da3b285e417dbfc5aef16  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic68515eee7d422be9cf8950e48b81d743d5491851d5a117d1f9b70d1d9b55060  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0ca47358f982879bb85bd78f6bc19192a5ed8c62214073342b37b040aea331b2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1606027ef88387f2150285b55cef89212359f49ab1a49fb71e457a3dba0c438a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic09f51154140ef91861243d7b35f05961565b368264d44c8fd5d0f85bd0fa213  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie28425115106f4b2405fad6fb2994a76e64dfa60e7bc165f46ae67411932a1cf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I64862889bfd7d2a15503bc07af594be59cbaa8758863f78311d6f15ecadcc99f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ied4424f3e85f3fb92f4e40bc63909f4e77698a18a1d0ee651e54e4de06ee330f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6c850d46af2f31f4e3d31c3fd2b2d9c7471ccf817b452a4fa2602485f5e7f164  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1a1a9f7ee74e17c4a0d7064ca9fae938002b1b685f3cb6309569081b0d971aed  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib5929b32be13a8436b74dadded1f26d3742e1424b6025d1eacda112bf4749a15  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibcb7809e1db6cb82ba62be017c5b8685cb6f988f85a0d29ce2459f6ac80498dd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idb971d0017094cf8b28e639623f85e6e5fc2c03a1da1e19a1ef87b959fe8e1cf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I89373d12365deb440d5337a2586fcdab81347ca28ff6f261a12e35a235bd23c6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib8f9b76d6cf7a74f0d437f634ce888096a0d6d81d66dc6c60b62a60006b661e9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie55394a5e3d49de60fbc4f33b3f9813b885da2049376036c935e8cd7c85010d7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6240db37d8e82731a264e5e3eeabb88e632dc6445647a26b4abdb142ff44c03  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4dfaddc409bf6d3698f255e55590182c2c8c067e0766311322460720dbd0967d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1dd3e1e1e78d9e24a54fc937e7a25fc0e2514eabd1c1cc662d81ba73aa44680b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I80d4a0cc8b63f2ce0dcb344da5a47c95cc28b5f93d5bc6b77e9b875cdd58db99  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iec19b0b63d20ea69dbcb23411a298bb6e833ee523fdf082f9343a695891a990f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib612f39370c6527c5f6eedb0eb5e7676212642673e940402586e823ddcbfb4c6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifa501efa24e47050960fb3c383458a20f54abcbc5ca45bbe2d15a037670cd5cd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8f088dd043a22011add21694f90df62fe1d2f6670cc72cfee805c9fb49756c77  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id86d515c6d081de87b9ed3c3521ab079e93ee082d8a0b396d44b3b70cac06b9b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4f94812066080b656de1a2807f5f669b2a81085bfc0470f9868bf5945856b451  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia92baf4463c96e210b460ea02d7775353edc6d475d7a315b594b9798cfd17900  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9d4c230c86454c5c5f9ec98917ffc8d23fd19105ef93ba860ac2650bcf43ba4d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia4a28d520896fadbeabee4130dcf862a9542852d87be480b1df2b67817f0ce65  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ide9498000905141bb106efc7e2184bd460d0e59a2270b10d42f981cf3bd514cb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie9a6b0e499ede3f80403e8f9c795ef4e93108ee8db755e12fb931259f1699712  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I362132341c8e8a464a2bc93e7cc5b1d9d7804dd93965614dc340b48fad5c92da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4b3c222863418745872c878545e419ee8f9c531f2cba89d28f0787992b0be8ed  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie39e570f1b5dd9f1ae893af78d81e458d077fcde2aeaba432209269b79785582  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I50ebc7f8f7cf324814b5885b2b18c90bf5007d8030744263d6e66880d836eea0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I326b57b49d3fcfe654c4cb9ebcd6edc0ad7969e3b531f498e3c31270a5c4aa70  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id3898be2185f86831f58bd16651edee3d1bb21fa07b33a1928740ab496404178  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2aa77512781cba636ab96a5d09527e1ac34623ea2bb6c6a8d742bbcf6eff499a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I225543794992ac9aa68ac3eeea38d41077ab5512b9f3b95fbd65a839294088e9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idd1dac44a6f35d558d400160a087fe7628ef80ad72c3962df2b3a3809b89bcdd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic039114ea8ac4120b09973c79fdc044251fc66bdeb18a498dd6ed7265cdfba2a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I21b3fa431ddc4bc8eacfb17a90fdac2bb32e4d0f4d0118715642c37601a1f883  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1c6d953c9a0e96d328cc4b515867b2ac21d2947a85e96be19f38e67a8b15001c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib823a58e9d4db87e4d73a81a772a02435af32a11d3c2265fb8a16021cfe4503d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3427390162b0952481e5f0728a20075c9cfb814431ecbb1a4014d407ab3b3afd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I35a9ae1cf23d8697091de65a1d0678632bd6889ae32408d7658e542a756e95ca  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I37e54e8ae28cf1a36cb9101d5afd4d523ca9a6ae244efe641c547a4114726bea  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9544a194d3d75c6c414169ea2536e111c09711ee602eb3462c4022350906a21e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e4bc72a55efb8462410905dcb2c9a8412e2533ded854d23ca648e0e36802960  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If2cec64e868d25d7fbad45ce4889c6a4cac0084aae00d2aa8963678edbb88875  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I73ad61911b0822e313aab2c484d1699cf2655a42a2bb0a1c9ab36228e41d0f7f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I218255d96e659dc8f60cddd40cac94a56d93556ed609b60157d88b298ec95f0c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11284a18d6115421b4c76054c1a580c41987dec66caa7d5bd9107bbd4ac8bc2c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8516ef195e4ba8f6e29a02ab5ea349a26bb68f6ebb4da847d56c03c942e9c20c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2411dfbbf605c7590bc678373dd20b7241356a433756332f9a3445ba8dad57fb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I69d896cdb2303b99b73c4d6886f2686381230feca86c62fc064a85e4d11266f4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If6ca882e537cdf5f458a2e11b7a11f057a3d2a00923825fe236afa0b0e1442c0  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie35443efbbf821e07284652a4b37347c4cfb959495dafa4fd2f81ffa2edc56db  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id6d0b1fe00e5324e0ed7c37d41ee3e848f9c7dcfb4a85f5da2b82ed4d8942b21  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0a309e8aa7f7e07abd837c99be6d8bb8c29dc1679b449111a02f49442d5cb432  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I416c7ff28cd1d182ba2e08c3882c04d5073a014f7b9b41e56a3850cdc289ffb4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie44d1a587dcdbb709546c6c567988fb0a19c276a1df7aced4c09a029196dfd4b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic2b8d811fd01f5cd88dd60bb1b89b33163b3cbeae48d04e2316f15500c6a1a40  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I85ff9ab4f9a4a3301bb8fcdc7107202263af0c37f091445efb5fa163a6b47a51  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I39ab1bf4bdde9805c5bc7695c4700975d5a6094c40e107b82477192005d9ce21  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I602591ae56f1a42c64e50378841e065e79aee138622a0a571effe20cb48645a3  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If37e9ed3af8a31c989dc6ad554207cd464c591b630ca1e5cf56b2eca57a18d8c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I80099c7b01770cc5f7edb3a3551d8edfe9dccbcd2a12daf8ebbafdfccd141bd4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie479ccbabaa8a00009152557e4de08bd240fd28f1b131c674dafbcc2505711f7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6364406b04427fe3a4cecbed48e12a67cb08dc632b2914b0fe52fab0ca541c0d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I610dd39f1d44d84764b0acd6b3fb1219fb6b6d6ca92e1b226ca76a389bf6c937  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib9f9384ac4ec4bad29fbb4ce683ffda7dcab311135f02b6336e6209f5742fddd  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I60980f76d468775bcc8a7052681fbb6ef4b2243e5e30e5365cda6cf598bd0bde  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I892a754f0322d92126d4731e8066760a24897f93e2afb858ee1393604d2cbb26  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib0f8816eafd3b950f67cfbdb6a44c59ab7c0918979817a4a998d8305da847e72  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I04b55f2c45002f1f1f7a6176773a22730dcfea14662f0badb102ddb60b84cf9d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5edc072d158ac583bd1cdb2449086d4f0b17e36d724f4cfde79820788ce57f31  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ieb128919ed64e331affb6adba798c267e8c3ec924a7ef58f50b1bc0b29702c23  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I90cc372cc2f3b23eaaf2cb32da95ee715af64ca2eaee77195d9813647d2a0d08  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idaf65411d995039ea730b6ee4b5ae727325da17dc79c8664270d60f063828453  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I977557441002c273f9b9b8748ffa9edceadb342e028ceb581c3bbce9af103a74  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icc10ac19a64065f5923ecef4f1353f13c7796c23f2555f8ae6566eb538d77677  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I725c369a5013eeb6b581209bc8a921fccfcf1754137191e26757abdb72ced94b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaa02b7ddfffcecb763aa916a2bc4c3aea58027c89b515c40b72214d9dd44ba21  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If8737fa82b71d9b0e7223baabca7405e148621600bdaef02e65cd7bd175b2d88  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id85c2b905d61bcdc87d500d6ede3ca02d52bc3eaf278f087f27fe6f277c91262  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I5923f41aa444bebfc18d13202747ff84e20a4753bc9cedf697b9ae8ec3418afa  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I4ac498dc826a9dbeaddf2f013ae7116e92dc772ea55987a4661f18e56a4123a8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaadbb1b235a85c555a6f37d003e87a987b7d9b07148207555eb717b7332f67ec  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I6afb533ec993de4f9b04007b355a9cadf08488ee6ca02aec2d7916a4c98a7fad  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I01313177417c899543a67763ede925dea3ee58ef4a31714ad15a7a3746bb5be5  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibd0ba147d1a08acea707b8c60da14ebcc4ad62e67ef26634777b5dae38af6d61  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I1e92e18a915678cc96aa493a00627dffecbd341dc8e022615610061e52c1ac3f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia7b91fa4a1ef16f859ee162b91daedc97927244dc19aaedede898049daf85a19  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I9918d91748722a47f8526008bc3fd4c498bc80205211d5c92acbc511fdb667bf  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I95d109e37a87827de1455b5ec479dda78a0218cb9db245b80710cdb1e8ead67a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia0c7162290e415f24699688e45850c243397b5cccf07daf0398dda04810b0690  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib9dc17b2b9fc7c228eba40cf625a49a27ec16f8c8a91957de14fb6849ea49212  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ied32ced79448b3f92faf0dca1673559e07372ec338e8c51a750be1c6975a298e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaddb000276bde734c13ec1395f06c1b3bf5606ad5cb138579d711cecf26ac88a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I211ada7f9095ced6b3d20f8f7f67b56cd2e73595481ed5d4c08175ca874d16ae  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I0d49182fe7486bcf54c8f68904b4b90436de6f3bc42fab67a4e47f61154e22c4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          If79b91295d25c503f6bf5ca7c6eebd2ebf6807dd9990ce31e844cee0d8f89dac  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iec1d04d20ec09595743b7a35860b5cb2ec862c20da87c6f899284069c60bdd71  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2126b1597a95d7aeb7d20d4e0f4270e1fc5cb0fe6eb5003b05abbb7e5e9a2819  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I72a115d9b3659f31366e1d73d6d9a0793e20be233c3ccab2b513fd79786224bb  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I469b0bcfe9cfc27a8596782bab479f30aedaa132a5cd404feb1fec4b52a17d3a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib4c52550766a2cbe0de236d6783edfb1a6a7cb4c2bb9333a9379e1b75680dad1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaa72101e8c3e7fa248ac4d4336b3847c4f602b6db009e9cd74cdd25251d5178e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic1381219782d18c1cb880970c062eb260d9d3be0b597e1465fc604c0c0c32c68  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icf0c3c82c9e458a347212415d3029f192c40152e8525a20b5c9bfed88ccdb32e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic5a87abf4c6018e9555de321c141d9754a7de91f1743d980e339ff9cebd63b7a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3a27e4e3322c28e7fe85d7e76b7d5477f4d4f6acb8cdb876b9a54cba98b189b9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I11edfeb948852dab396975b53b12d09da7a5fbedc2dae9fe7c687768cfef05b4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I578437932d2d1156445b41a1238e0fd96ab5702bc3158ea337a9e37d14d6731e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3c2c5b5cd798851c7fcb0d0e66ddf81a516ef9bdf4aa4ebd4901532bfb2a651b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I8153d6f17d832da24daaba2909a88f1609e523ad3b6eac7ad42521979aae96da  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic10ea001dcd0b864b987bc3080e95b338c1e91247bb90e884e161c926183fd2b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I61efe7187a1aaa28235dacf68eb1e1dd97e7cb5900862790bb4d5872d7adbd67  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3c710fbd5e4dce0c97eb9da2d8e526f9d44d87fa75088c0421353614e6ef5da9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ie02f677979058dda2291ddb93acd64f4461f6d75f3a33c21dac97129344f7055  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I2b78100b50f7334d563daa27cab8078fa374dca0c438157d1ad44ed3fd9e3456  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Icdfa68bdad11213dbaa576cbf43ca9deeb1f9f24225264eaeeede7d1aba5fd8a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idb39db95234cbfdbbc89fdee230784c703e170b9e932643a5e1b811b24ae021a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7141b42fce475b5502fd33035bf37addde06271b2259e158ba03a66843b66075  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I245e922da0aa5470370db389d5bc9db33327c905528a1740aa015b7ccdfcc29e  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia2ff4d61c4f4fdf29be87b50e206c308cf970cbad2638e86ba8c2be8d025b534  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Idd383630385363471e1b17ea946a61194a3cb287d833af386876c3b4ee66e406  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3daa8702e9dbd047a05e5ea044d14b670c2ae3849526cc514be6a511c5c45c35  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia695c63ae87e9a6742c6fecea648a214f5b24ea2b652bb5d83f35d9a59b94f72  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ifc31b600cbbf26e78cee82cd354c17b872586c1a53ddd132edbd25ce87d8aa9a  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I261e70e693cdbc572e40e81c594f3dac624febb03465bfd0fb864d337e753499  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ia6f7ae0adde8136c7a25f4fed69bbcaa376b5f28cbb4990afabb57a87ec03019  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic40e94217a2d2c13f4b1ad2766ab1ae4e8ded0b5e0a3522dd51ec806c3e9feef  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I78602c68a4a00f530bda7ba1dfa4820b7faeb0edabc636d6a2d8bf97005755d1  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Id8e684d92e6d0b6e10b5e7f7ff9656e6fc67c99edaa59b49e453844ae33d23f6  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ic9d9001a209401fca8a3f28e39c4b89adc8f4e9d225aeffbb5d30893bea1a7b2  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I97f666707f6afacfc6156ef498941fe5feeb7424834b4a283139aefb5f50a68f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ibdaeb96b71f9ccccfe79b1b3bab77122aa32217b58037d80a3183bf888b60c72  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I574e4843ab81be7ad95cb7027fc3284a8780b07fb8a194a9c991997988d7ff8f  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iaa4463f258ed92a2c85fef0790c47e725c555f37c80dbe366d973c9599a5484d  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I7102386e760e34e2d0fc4563b497acec7222bd171333a2169fac800df94ea27c  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iee34d958bf4feec1e5bde8a866a9919f29edd54f1bc51cc9c8216b71101d640b  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I64b0ef6642050de0690c95be2af9606797be36c1656f1306b87ce3e8131c4629  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I23f31ebee34c7f4f9c46fba41d41df176a7465c074ad8527205a5782edab6524  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I628b9674d7d6caaa70c54539241df2e7a4be0441dde1739b442513c6e4ded8a4  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Ib066c9d790586949b27c4cf09dc957e7d28161ab00e8dc6920e4e0cc5ac665d9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I57419941b1979cd06c4fa0e6be943f004dd80da502425ee5b6dabd2239139cd7  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          Iabb5703a54942b1bdcfe2213d2011c659ec812f751dc75943b2ce511c81ffaf9  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I798a6a6074b50fc61bd4e1b4696560abd2e515c86d47f85e9a3077cf6672acc8  <= {(MAX_SUM_WDTH_LONG){1'b0}};
          I3f4a8ec7c554b1f0b9d3d2963b0e3dec4654bf07c5b836f8fd07c639cd19d588  <= {(MAX_SUM_WDTH_LONG){1'b0}};
       end else begin
            // I09394b7939814acd4a58cfd06095eef5e15b8426cc1eaf428c87f25cca6d3777 and If076b994bfc2fa6c6de92c2e43a8779943e97717abb5b9c62225518daff111a0 If86b1f62a8554232b940f4fd9c8d6601aae4767456df3d6cdff55a51f17b5075 I9c19636ddea25f0a13357d01c0aef27a4eb4c7f8cbaf2be35f272273572ce2e5 Ib8d31e852725afb1e26d53bab6095b2bff1749c9275be13ed1c05a56ed31ec09 I0967115f2813a3541eaef77de9d9d5773f1c0c04314b0bbfe4ff3b3b1c55b5d5 Id8198efa3604d164853468608c55efa148bc56e3564d5a30232bf98b8ab43aeb
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[0] ) begin
                    Idd9957e5b52c4d33e24910559d8203415afdf467bbe1c9de950145282c7eacf0  <=  ~I893355bf7ee2fbac8f9873385982e6b24128db3c9934e37db7bb8b576a4ac41e + 1;
                end else begin
                    Idd9957e5b52c4d33e24910559d8203415afdf467bbe1c9de950145282c7eacf0  <= I893355bf7ee2fbac8f9873385982e6b24128db3c9934e37db7bb8b576a4ac41e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[0] ) begin
                    I7fbf7b7f7a1f0155cb188ee4219620cb35a2fcf98d2687cddfa2508273b70154  <=  ~Ic1d44b04503cdaccd5821f80e822659de6f6e305c3206e603ef6e23dd3dad3ce + 1;
                end else begin
                    I7fbf7b7f7a1f0155cb188ee4219620cb35a2fcf98d2687cddfa2508273b70154  <= Ic1d44b04503cdaccd5821f80e822659de6f6e305c3206e603ef6e23dd3dad3ce ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[0] ) begin
                    Id658b37d70ac8e3a324133f475a77c7948231571aa66ea0dd11b6460fca011a3  <=  ~Ia02e90fa0c6b93819416a3059cf6adaaee9c396532e724c47648f414a16679b6 + 1;
                end else begin
                    Id658b37d70ac8e3a324133f475a77c7948231571aa66ea0dd11b6460fca011a3  <= Ia02e90fa0c6b93819416a3059cf6adaaee9c396532e724c47648f414a16679b6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[0] ) begin
                    Ibe0fac26b5e106fc1753aeb842e8a04067fc91c95e358b1caa58db8192381837  <=  ~I43f540ed8151f48307326f27534afca5105989e179c37e992cc8516996b10bd8 + 1;
                end else begin
                    Ibe0fac26b5e106fc1753aeb842e8a04067fc91c95e358b1caa58db8192381837  <= I43f540ed8151f48307326f27534afca5105989e179c37e992cc8516996b10bd8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[0] ) begin
                    I1a2646b8251f83855c3fe8f6172f36500201ce43b9b5ba2cf0f25fd5d540e89c  <=  ~I3d7d9699881b5d4d42cc19d1489f8116cf6f3eef7781b1fdc8cdedda72233a32 + 1;
                end else begin
                    I1a2646b8251f83855c3fe8f6172f36500201ce43b9b5ba2cf0f25fd5d540e89c  <= I3d7d9699881b5d4d42cc19d1489f8116cf6f3eef7781b1fdc8cdedda72233a32 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[0] ) begin
                    Ib3a2af9bef5f5d8d7228a3b49a5e0d4a37a33117e057078a552588a24d46addc  <=  ~I1b0a3f720c3ed13e66b1c568162495031330a4369a4d0ddf65848c307e1d56e6 + 1;
                end else begin
                    Ib3a2af9bef5f5d8d7228a3b49a5e0d4a37a33117e057078a552588a24d46addc  <= I1b0a3f720c3ed13e66b1c568162495031330a4369a4d0ddf65848c307e1d56e6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[0] ) begin
                    Ic072a2fb2ce65ca734c05e747f12ad094cc5aaf9267dd94dba345b5c7b11dcdc  <=  ~I1927b4579e43362f62245cc1904e0deea9705e4427e3bbaeece21a3e36820df6 + 1;
                end else begin
                    Ic072a2fb2ce65ca734c05e747f12ad094cc5aaf9267dd94dba345b5c7b11dcdc  <= I1927b4579e43362f62245cc1904e0deea9705e4427e3bbaeece21a3e36820df6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[0] ) begin
                    I01d7d3d20ba0eab63d519ae054b6c22c5be4000c846a6a4883ffbbddee37663e  <=  ~Ia341cb94dc5268759917bc49586f20130d999dbbdcd5f1b34e576770d6d063bb + 1;
                end else begin
                    I01d7d3d20ba0eab63d519ae054b6c22c5be4000c846a6a4883ffbbddee37663e  <= Ia341cb94dc5268759917bc49586f20130d999dbbdcd5f1b34e576770d6d063bb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[0] ) begin
                    Id0f930aa222bd91b8a7d5f80a38d84993a63fa1c6aca3d37ed259294e08869d8  <=  ~I34d68a357aa2b44cf3a3b08384498af0e4cc195b0c725a67769d62e36877cb7f + 1;
                end else begin
                    Id0f930aa222bd91b8a7d5f80a38d84993a63fa1c6aca3d37ed259294e08869d8  <= I34d68a357aa2b44cf3a3b08384498af0e4cc195b0c725a67769d62e36877cb7f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[0] ) begin
                    I236cce67d0aea9f9c8d5ea3c39cb598d55f734b44ad6e3972e7f6b91d56001fe  <=  ~I48a2995df1784de9dc4a3b951d711905f920ed0b9fc0e20ee48f8838a3ba6502 + 1;
                end else begin
                    I236cce67d0aea9f9c8d5ea3c39cb598d55f734b44ad6e3972e7f6b91d56001fe  <= I48a2995df1784de9dc4a3b951d711905f920ed0b9fc0e20ee48f8838a3ba6502 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[0] ) begin
                    Ibbbf3f4aa7f74c37a0e8ac8a675ac9a9fec748ac720e6a78e9cf937dd089b8e3  <=  ~I45e3ffea730c76c713d1e61276b644a026af54458af4d3894e44c4416f9e4867 + 1;
                end else begin
                    Ibbbf3f4aa7f74c37a0e8ac8a675ac9a9fec748ac720e6a78e9cf937dd089b8e3  <= I45e3ffea730c76c713d1e61276b644a026af54458af4d3894e44c4416f9e4867 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[0] ) begin
                    Id27dfca888552262f492b81fd23b881938f66eb15f7ab21afb210fc6056fa09f  <=  ~I573b8edf32c67a0863b9e9ecb44ce7154a48ec67472c04821ffcb202bf3b28e4 + 1;
                end else begin
                    Id27dfca888552262f492b81fd23b881938f66eb15f7ab21afb210fc6056fa09f  <= I573b8edf32c67a0863b9e9ecb44ce7154a48ec67472c04821ffcb202bf3b28e4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[0] ) begin
                    I8db02445666e4aa12d7e495ba28ca0eae6ef411094d30330e91eb9eb03b38aa7  <=  ~Ic2544a607bb965371402190fd2fe4afbd85977e8360b5f0091a6f11f885909c8 + 1;
                end else begin
                    I8db02445666e4aa12d7e495ba28ca0eae6ef411094d30330e91eb9eb03b38aa7  <= Ic2544a607bb965371402190fd2fe4afbd85977e8360b5f0091a6f11f885909c8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[0] ) begin
                    I3b1d695a626aefa8e5b146c7f7f26a8da119680783da7afb019209ac9fd719aa  <=  ~I1a641c18ed7edafaa7d5877ae724860b1d54fa6e6890510d1c7febf66944bc55 + 1;
                end else begin
                    I3b1d695a626aefa8e5b146c7f7f26a8da119680783da7afb019209ac9fd719aa  <= I1a641c18ed7edafaa7d5877ae724860b1d54fa6e6890510d1c7febf66944bc55 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[0] ) begin
                    I82bc7aad8e3adf5b7bd03d9fdac6eea60cb800e4502e3af7bdc9d49139563fd0  <=  ~I7301f67cfc0739e38aae8830e112df2193600d9581476251265730522284b6b5 + 1;
                end else begin
                    I82bc7aad8e3adf5b7bd03d9fdac6eea60cb800e4502e3af7bdc9d49139563fd0  <= I7301f67cfc0739e38aae8830e112df2193600d9581476251265730522284b6b5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[0] ) begin
                    I422fb05bbac12ca5df13eb7c0c3fd96a4e819de9669ccd64d40060b5db3f3421  <=  ~I41ff59a42cce4bf7225d8f9296ec89aab75a0ec2dc10f0c341c696fc2461ce3a + 1;
                end else begin
                    I422fb05bbac12ca5df13eb7c0c3fd96a4e819de9669ccd64d40060b5db3f3421  <= I41ff59a42cce4bf7225d8f9296ec89aab75a0ec2dc10f0c341c696fc2461ce3a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[0] ) begin
                    I7200758287b0c7ed92552ced989756e1d49b5418181b9e36421da7e2694ed3a2  <=  ~I799ec6460c042feab5ece45c8877d0614bfea4ebd97b427e1bd00aaba217c1c9 + 1;
                end else begin
                    I7200758287b0c7ed92552ced989756e1d49b5418181b9e36421da7e2694ed3a2  <= I799ec6460c042feab5ece45c8877d0614bfea4ebd97b427e1bd00aaba217c1c9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[0] ) begin
                    If34d8ceb2732716c923a7f250495970948ae431d5f1e0a025618c1070940ec39  <=  ~Ibf5e207961c05c6ea8ee1cc657aa7bf8a0fd7827e4e550b65cb9cc20925f7536 + 1;
                end else begin
                    If34d8ceb2732716c923a7f250495970948ae431d5f1e0a025618c1070940ec39  <= Ibf5e207961c05c6ea8ee1cc657aa7bf8a0fd7827e4e550b65cb9cc20925f7536 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[0] ) begin
                    Ibdd37577b403da9aa72ec3f4707379b1151c0b15edbfc4fd304c4e35c1672da6  <=  ~I1ce1761a25063d6ca639d1aa9094a30899744186121a71229f255eaf3542b80a + 1;
                end else begin
                    Ibdd37577b403da9aa72ec3f4707379b1151c0b15edbfc4fd304c4e35c1672da6  <= I1ce1761a25063d6ca639d1aa9094a30899744186121a71229f255eaf3542b80a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[0] ) begin
                    I6201d3c2d85bffa03f368b5862fba1b2e0ce3735fcc8711cb8107adf16ccdeb9  <=  ~Ifa331e88bb390c67efa83efdb978b28023c3f4a74750928415242eff2a75326a + 1;
                end else begin
                    I6201d3c2d85bffa03f368b5862fba1b2e0ce3735fcc8711cb8107adf16ccdeb9  <= Ifa331e88bb390c67efa83efdb978b28023c3f4a74750928415242eff2a75326a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[0] ) begin
                    I34f861f0a748b0ad1550db8ce40149dc638194b0089cf22e2380a39a49f8c902  <=  ~I7e5dd2b4a968c805518feeef59ac29c86d9c06c30446f8966bff4b169c65962a + 1;
                end else begin
                    I34f861f0a748b0ad1550db8ce40149dc638194b0089cf22e2380a39a49f8c902  <= I7e5dd2b4a968c805518feeef59ac29c86d9c06c30446f8966bff4b169c65962a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[0] ) begin
                    I73ce2860dd9aa9ca2c0d541a6ae1e5069badd35988d922cffb6aef0038cde662  <=  ~I9663885f1f636653b6649709c8859bdf9e407c18311f63a0e6677f6671926884 + 1;
                end else begin
                    I73ce2860dd9aa9ca2c0d541a6ae1e5069badd35988d922cffb6aef0038cde662  <= I9663885f1f636653b6649709c8859bdf9e407c18311f63a0e6677f6671926884 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[0] ) begin
                    I07c37e958136be68b3d658649964c73ca78160582248da1d45eb9ee82c1f679b  <=  ~I9e8163c831756fc1d31bf9bb6e966a5c58738673504240801b73891e606845ac + 1;
                end else begin
                    I07c37e958136be68b3d658649964c73ca78160582248da1d45eb9ee82c1f679b  <= I9e8163c831756fc1d31bf9bb6e966a5c58738673504240801b73891e606845ac ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[0] ) begin
                    I0aafab9f9205eb4a8c16e213e116d949a5c625f7cb2b0f3d124deb80aad2c6c7  <=  ~I211a4aa442cd695ebef8bfdd8734fca64e796eec6eaeae0f7c1c306d89ac50ad + 1;
                end else begin
                    I0aafab9f9205eb4a8c16e213e116d949a5c625f7cb2b0f3d124deb80aad2c6c7  <= I211a4aa442cd695ebef8bfdd8734fca64e796eec6eaeae0f7c1c306d89ac50ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[0] ) begin
                    I96fb06aca6108479f7e21e1835a091a9060c2925cc6320c8ed71a0a0092bdeab  <=  ~I2e3ac37a60fed64971c398ea5f48490f1a8ba9c0fe63583d4996ef4884aa0eea + 1;
                end else begin
                    I96fb06aca6108479f7e21e1835a091a9060c2925cc6320c8ed71a0a0092bdeab  <= I2e3ac37a60fed64971c398ea5f48490f1a8ba9c0fe63583d4996ef4884aa0eea ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[0] ) begin
                    I11c6d693bd6c019722571e1aa6eea0507f351a89cfc6d16f8fc51997981aea81  <=  ~I71f710555439b202404f08c784a66fffed0e12c7dad92ced1b83a6f28245a512 + 1;
                end else begin
                    I11c6d693bd6c019722571e1aa6eea0507f351a89cfc6d16f8fc51997981aea81  <= I71f710555439b202404f08c784a66fffed0e12c7dad92ced1b83a6f28245a512 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[0] ) begin
                    I65b0824920910c82c7d677c2dcf4216e86940b3edc0b3da85d8f65505f58ad48  <=  ~I458d537d6f291b854051834fc85511253dbd0054f1be7bde7ac2696c4e4424ca + 1;
                end else begin
                    I65b0824920910c82c7d677c2dcf4216e86940b3edc0b3da85d8f65505f58ad48  <= I458d537d6f291b854051834fc85511253dbd0054f1be7bde7ac2696c4e4424ca ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[0] ) begin
                    I37084afdf6695d3b8fb0530643c8b03deb2499f4f68ead04e3b5b79aa4467f73  <=  ~I3e27399b8d9e65418758d9dca1b1cfbcb4d908000611b218f4ad2097da556a51 + 1;
                end else begin
                    I37084afdf6695d3b8fb0530643c8b03deb2499f4f68ead04e3b5b79aa4467f73  <= I3e27399b8d9e65418758d9dca1b1cfbcb4d908000611b218f4ad2097da556a51 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[0] ) begin
                    Icc43ea934f0c07465170977b52d2f402fe155ef77f3ca27119fa665a1d918694  <=  ~I38ef2b3fde182cebc6e8265c6e99d08e21e28d55b2eb1b7a161f13e385ac5b72 + 1;
                end else begin
                    Icc43ea934f0c07465170977b52d2f402fe155ef77f3ca27119fa665a1d918694  <= I38ef2b3fde182cebc6e8265c6e99d08e21e28d55b2eb1b7a161f13e385ac5b72 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[0] ) begin
                    I1622b11941b00f6d2ecd90320158533a66501a6ddb78defb4464a937f132c232  <=  ~I0f2d9a8f6ab682ae8c5fb31b30d5c11be65370398f373fda27a64bf6d718193c + 1;
                end else begin
                    I1622b11941b00f6d2ecd90320158533a66501a6ddb78defb4464a937f132c232  <= I0f2d9a8f6ab682ae8c5fb31b30d5c11be65370398f373fda27a64bf6d718193c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[0] ) begin
                    I252a77c3eaec2d6accaee6de3ba5d0b354636e2a2aef4992eca0e2a74eb4d25f  <=  ~Ie504e487c65a8cf270fcb907ff7a6f204c5afe50af53c0b0279719522b595c19 + 1;
                end else begin
                    I252a77c3eaec2d6accaee6de3ba5d0b354636e2a2aef4992eca0e2a74eb4d25f  <= Ie504e487c65a8cf270fcb907ff7a6f204c5afe50af53c0b0279719522b595c19 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[0] ) begin
                    I17dbb17fb2770beac552dafeb238c5e8e7a948c35c7c543508e652cbcda01dee  <=  ~I7306fa7f8f192749aacf00bcfc3ee6266ad06e373f4075503bf8c7daa963f7b6 + 1;
                end else begin
                    I17dbb17fb2770beac552dafeb238c5e8e7a948c35c7c543508e652cbcda01dee  <= I7306fa7f8f192749aacf00bcfc3ee6266ad06e373f4075503bf8c7daa963f7b6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[1] ) begin
                    I96e7a523360a0cc0f3abfea09a566658e5e9f3316c3c412f99fd6340d1b64235  <=  ~Ica9704300b0989fb0bb8dd9ddc1807a4906458c6f7f487fb7d7e214e31458eb8 + 1;
                end else begin
                    I96e7a523360a0cc0f3abfea09a566658e5e9f3316c3c412f99fd6340d1b64235  <= Ica9704300b0989fb0bb8dd9ddc1807a4906458c6f7f487fb7d7e214e31458eb8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[1] ) begin
                    Ibadfd4f0852067e83ba6f0d57699585ae20eb542d1ad8f2cce3bda0d043ff2e0  <=  ~Ic8e52a8db0d0cf4d90f46c2d5b5871d31db974cbd84b5e68f4d872ccb6fb9cf5 + 1;
                end else begin
                    Ibadfd4f0852067e83ba6f0d57699585ae20eb542d1ad8f2cce3bda0d043ff2e0  <= Ic8e52a8db0d0cf4d90f46c2d5b5871d31db974cbd84b5e68f4d872ccb6fb9cf5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[0] ) begin
                    I45ade5cafdcd254cc640ea8725da6961717fd6c50f747242aab6976ace4e8f10  <=  ~I59ef74fe764da43c107f5eb1c48cc198be3cfce3b3c55e0eac3efe7c9af888a0 + 1;
                end else begin
                    I45ade5cafdcd254cc640ea8725da6961717fd6c50f747242aab6976ace4e8f10  <= I59ef74fe764da43c107f5eb1c48cc198be3cfce3b3c55e0eac3efe7c9af888a0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[0] ) begin
                    I597d0e1b64b5d47502804c7ba47fd0c17322bfdbd4d332b11f9742713f76855f  <=  ~Ib33fa9a97b26fc69be1d69ad97dcc345c1701bd9ca2fb0922d724237bd2cf8cd + 1;
                end else begin
                    I597d0e1b64b5d47502804c7ba47fd0c17322bfdbd4d332b11f9742713f76855f  <= Ib33fa9a97b26fc69be1d69ad97dcc345c1701bd9ca2fb0922d724237bd2cf8cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[1] ) begin
                    I8c971b4c1be575fe328c0a4a9ecc5dc75f08d36f65aa58642976d971a6c316d7  <=  ~Ibc1655e6f13d450c6beb85bc81ffd4b765ed49cb361ddcae84e6e635e85513da + 1;
                end else begin
                    I8c971b4c1be575fe328c0a4a9ecc5dc75f08d36f65aa58642976d971a6c316d7  <= Ibc1655e6f13d450c6beb85bc81ffd4b765ed49cb361ddcae84e6e635e85513da ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[0] ) begin
                    I982c94b61dff8249f2f3055f60da6e2c2b0b56c403f151168b28a5a211aa6428  <=  ~I170b2f3df88d573e89dcd7abd2e33192d1e08eb33a333dab67be7795d2371e04 + 1;
                end else begin
                    I982c94b61dff8249f2f3055f60da6e2c2b0b56c403f151168b28a5a211aa6428  <= I170b2f3df88d573e89dcd7abd2e33192d1e08eb33a333dab67be7795d2371e04 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[0] ) begin
                    Ieb5e001b45961175497657da7a0340c2a15b6d8de1b72ad68ac3aa7f96a47af0  <=  ~Ia554b8c5dc66b7db32a935b99a2e41aa84c6c13fa944f2de90eed8c1d462d023 + 1;
                end else begin
                    Ieb5e001b45961175497657da7a0340c2a15b6d8de1b72ad68ac3aa7f96a47af0  <= Ia554b8c5dc66b7db32a935b99a2e41aa84c6c13fa944f2de90eed8c1d462d023 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[1] ) begin
                    I9ab473d34fac3327f03768e14c7bb20056aa8a3dd31520d385552eb6d214f890  <=  ~I60e54e7e8d975cee4bf0823ff91ce212f02e407e9e2064ea4ca882ba4961553f + 1;
                end else begin
                    I9ab473d34fac3327f03768e14c7bb20056aa8a3dd31520d385552eb6d214f890  <= I60e54e7e8d975cee4bf0823ff91ce212f02e407e9e2064ea4ca882ba4961553f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[1] ) begin
                    I4177cb2b0a83442a271f59bf4f758851d5146ee00d76a1177c9a34d4208b7c09  <=  ~I4470cc46d92649aa472f4dce99afb05681b554782384542942fb243099cfc6de + 1;
                end else begin
                    I4177cb2b0a83442a271f59bf4f758851d5146ee00d76a1177c9a34d4208b7c09  <= I4470cc46d92649aa472f4dce99afb05681b554782384542942fb243099cfc6de ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[0] ) begin
                    Ie46448d24890ed6ffa2736abb97331dc3ed219b9324bc0e8453eed6aa2a4806c  <=  ~I9f258a7197af9b66d573a49b5923adec1c8637c53af4c2073805fa31fef73dfe + 1;
                end else begin
                    Ie46448d24890ed6ffa2736abb97331dc3ed219b9324bc0e8453eed6aa2a4806c  <= I9f258a7197af9b66d573a49b5923adec1c8637c53af4c2073805fa31fef73dfe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[1] ) begin
                    Ie000dee1e3953811fe9424588b71a7dbc88f41ec69afd16e17e8fabf141c31ec  <=  ~I52497162427ed0e9f305f509a79ddbdd02f12eebc337f57d63a9e477ce556e44 + 1;
                end else begin
                    Ie000dee1e3953811fe9424588b71a7dbc88f41ec69afd16e17e8fabf141c31ec  <= I52497162427ed0e9f305f509a79ddbdd02f12eebc337f57d63a9e477ce556e44 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[1] ) begin
                    Ia96c921ce4e0590c903d02dc69790c6af52898da90f4766121fa7b31e0ce6190  <=  ~I7d53fc143b190930a55ef8fcf893ea0b45d87abc54330c08bf4b4d5c67d4cbda + 1;
                end else begin
                    Ia96c921ce4e0590c903d02dc69790c6af52898da90f4766121fa7b31e0ce6190  <= I7d53fc143b190930a55ef8fcf893ea0b45d87abc54330c08bf4b4d5c67d4cbda ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[0] ) begin
                    If9628510f239b2275efec7ce187b8eb7360beb042a425934ac81632815361368  <=  ~I7f819482e0a2454a58a949963a2600e43477da52fcac968f397cade6b69be570 + 1;
                end else begin
                    If9628510f239b2275efec7ce187b8eb7360beb042a425934ac81632815361368  <= I7f819482e0a2454a58a949963a2600e43477da52fcac968f397cade6b69be570 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[0] ) begin
                    Iaf205cfa67ea9b2c39d6705da465f081eb75c326c1d80e63e1331a098ca9a4ac  <=  ~I551c9d548f30a033083c22bbd3fb8c0ad11c32fbbf66ccc8d0f6b7a177a49b39 + 1;
                end else begin
                    Iaf205cfa67ea9b2c39d6705da465f081eb75c326c1d80e63e1331a098ca9a4ac  <= I551c9d548f30a033083c22bbd3fb8c0ad11c32fbbf66ccc8d0f6b7a177a49b39 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[1] ) begin
                    Ibadbb4e272ab1105914763e2790898c8e37a553a1b6726e8818431bf5209b369  <=  ~If00a6af912a327873844b41dfbbcb9b7383e07272e5eb09cdf9b4a4a827b4f1f + 1;
                end else begin
                    Ibadbb4e272ab1105914763e2790898c8e37a553a1b6726e8818431bf5209b369  <= If00a6af912a327873844b41dfbbcb9b7383e07272e5eb09cdf9b4a4a827b4f1f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[0] ) begin
                    I6dcc482b16866339b78b922f9a7ec0f4a0ef311c353e6a4e107dfcc351abbb23  <=  ~I770b9333cb3aebf6d60d58661bc3282c1fed64de0824268f9f7aaa2dad91efc7 + 1;
                end else begin
                    I6dcc482b16866339b78b922f9a7ec0f4a0ef311c353e6a4e107dfcc351abbb23  <= I770b9333cb3aebf6d60d58661bc3282c1fed64de0824268f9f7aaa2dad91efc7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[0] ) begin
                    I41a57b30ab1dd9c40a723f99315558a47412465aa3fe967250572e8373aa7180  <=  ~I27a121a528b8c373659d1b04c8b5eaf5856b441ddf1b24331855326f31bfc492 + 1;
                end else begin
                    I41a57b30ab1dd9c40a723f99315558a47412465aa3fe967250572e8373aa7180  <= I27a121a528b8c373659d1b04c8b5eaf5856b441ddf1b24331855326f31bfc492 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[1] ) begin
                    Ia042bc20eb6866de0ab9ca9154f0db63f7d4ad84d553be858a0be88fbb8f7f33  <=  ~I044870873609a6dc7acef74d59eaea493c553cbcc3eff5b580dfd6a8f176d987 + 1;
                end else begin
                    Ia042bc20eb6866de0ab9ca9154f0db63f7d4ad84d553be858a0be88fbb8f7f33  <= I044870873609a6dc7acef74d59eaea493c553cbcc3eff5b580dfd6a8f176d987 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[1] ) begin
                    I782d29ca9e53ffe86cec8809d7d413c9c5ebd9edb6a0d76db2d0c321312d224a  <=  ~I1db3917cd01f808a2a2f4c78ef1ed3328ca804093065a1cfb9e15ef210bb8c93 + 1;
                end else begin
                    I782d29ca9e53ffe86cec8809d7d413c9c5ebd9edb6a0d76db2d0c321312d224a  <= I1db3917cd01f808a2a2f4c78ef1ed3328ca804093065a1cfb9e15ef210bb8c93 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[0] ) begin
                    I9342de9fe82f2273da138f99da619acf144edf1f9c33682fe3b1a09d0121c4d1  <=  ~Idd38249645258d9f8ef1e5cfbda4f15a700ff3b6d78b9c202bfbeca278528f57 + 1;
                end else begin
                    I9342de9fe82f2273da138f99da619acf144edf1f9c33682fe3b1a09d0121c4d1  <= Idd38249645258d9f8ef1e5cfbda4f15a700ff3b6d78b9c202bfbeca278528f57 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[1] ) begin
                    I6a09910e62aa0cf665f69be80c9ad61f2d31115012314b8188cf79fae365626c  <=  ~Ie2757ee84c5d0e87b17c22db78eec37478ff53ed9383587a3afa0e3270afde8f + 1;
                end else begin
                    I6a09910e62aa0cf665f69be80c9ad61f2d31115012314b8188cf79fae365626c  <= Ie2757ee84c5d0e87b17c22db78eec37478ff53ed9383587a3afa0e3270afde8f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[1] ) begin
                    Ifcc25cd8dc442c6720ac0f764b432530aa63681953d8ba16b441892ff5966bfa  <=  ~I85ce012ac5bad111ae4ab945035baf1b2820c82822f28a7b7c314515345af8a3 + 1;
                end else begin
                    Ifcc25cd8dc442c6720ac0f764b432530aa63681953d8ba16b441892ff5966bfa  <= I85ce012ac5bad111ae4ab945035baf1b2820c82822f28a7b7c314515345af8a3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[0] ) begin
                    Icdea1f407aaefacb918babc28247d540a8a52d513d26d7fbb5e81a41797e7555  <=  ~I89db4b6e1da27586c9fb92f89e492af68c0497029c97adbcdd5e3facac07c213 + 1;
                end else begin
                    Icdea1f407aaefacb918babc28247d540a8a52d513d26d7fbb5e81a41797e7555  <= I89db4b6e1da27586c9fb92f89e492af68c0497029c97adbcdd5e3facac07c213 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[0] ) begin
                    I954e0367a6f3af96a7e033da51e7256543d7eabd37191d4b03f3077567cb629f  <=  ~I3bdc9359c749bc85fb3a7fc68446c47edf3565e167d9a28caf4bf5010b95a575 + 1;
                end else begin
                    I954e0367a6f3af96a7e033da51e7256543d7eabd37191d4b03f3077567cb629f  <= I3bdc9359c749bc85fb3a7fc68446c47edf3565e167d9a28caf4bf5010b95a575 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[1] ) begin
                    I78abc91706fec0893eee10a69916f7247b718169155038bdc0bb6f8661ed1c3a  <=  ~I09a731c0252003cf8c9e4848c2e8ecb6a86e0bf4d76ed8fe028e3a609d639aaa + 1;
                end else begin
                    I78abc91706fec0893eee10a69916f7247b718169155038bdc0bb6f8661ed1c3a  <= I09a731c0252003cf8c9e4848c2e8ecb6a86e0bf4d76ed8fe028e3a609d639aaa ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[0] ) begin
                    I30e28a0e32497e3137bb689fdbde46389bc490300e15be88612f28eff07976e6  <=  ~Iae3ca8fe4281bb23b5ed7e87317e7aea52a130420731529f44179ea0274a58f5 + 1;
                end else begin
                    I30e28a0e32497e3137bb689fdbde46389bc490300e15be88612f28eff07976e6  <= Iae3ca8fe4281bb23b5ed7e87317e7aea52a130420731529f44179ea0274a58f5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[0] ) begin
                    I25779b63a47c05d4588d4b33fecaff61647609a62fcc90f0f541c6b30ea9342c  <=  ~I38f8f9e2731f858a15a6f2f3a375d0d29634c0da467767e21318213ae7beee7e + 1;
                end else begin
                    I25779b63a47c05d4588d4b33fecaff61647609a62fcc90f0f541c6b30ea9342c  <= I38f8f9e2731f858a15a6f2f3a375d0d29634c0da467767e21318213ae7beee7e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[1] ) begin
                    I1d91c7e9c2f99df4e0523b7e01b6fa6ea3930382238ccfbc07201b7d3edcc969  <=  ~I01eae75c6d18bb06d82fd21bc1aaf1cb883bed514f5497fbc433fdc42d217535 + 1;
                end else begin
                    I1d91c7e9c2f99df4e0523b7e01b6fa6ea3930382238ccfbc07201b7d3edcc969  <= I01eae75c6d18bb06d82fd21bc1aaf1cb883bed514f5497fbc433fdc42d217535 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[1] ) begin
                    I9095fb177f965807ae5a73a45c76b1c0b6300c6800b17259e5836adea5a78ec8  <=  ~Ie5a56b54b520cb4b1b0e5509ed4b3fa804bfc0be8566ed98b455a29b7148d291 + 1;
                end else begin
                    I9095fb177f965807ae5a73a45c76b1c0b6300c6800b17259e5836adea5a78ec8  <= Ie5a56b54b520cb4b1b0e5509ed4b3fa804bfc0be8566ed98b455a29b7148d291 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[0] ) begin
                    I907aa3f6584035b934017a601019d35f353b3f99c7573bef60fad167f9d9ffe0  <=  ~I0a4b485210baac225fd3f32b36be68140468a6c307f3f91de4416553421e3db5 + 1;
                end else begin
                    I907aa3f6584035b934017a601019d35f353b3f99c7573bef60fad167f9d9ffe0  <= I0a4b485210baac225fd3f32b36be68140468a6c307f3f91de4416553421e3db5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[1] ) begin
                    I58598429d44ad951f91139a213d3b0bdacac6d71f1b9753886dfe1d39d0024ac  <=  ~I172389b084abec531bf617713612fa0d8b27b0967bb62a6514aa873f609bb5b0 + 1;
                end else begin
                    I58598429d44ad951f91139a213d3b0bdacac6d71f1b9753886dfe1d39d0024ac  <= I172389b084abec531bf617713612fa0d8b27b0967bb62a6514aa873f609bb5b0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[1] ) begin
                    Iee510842ece3717ba6eefc3ccd844e97a9718788683d4c7ceaefa6ca0030585b  <=  ~Iff3e149eb4ce60c9f28638248c33ab96208976458886b1735785c2dba298121d + 1;
                end else begin
                    Iee510842ece3717ba6eefc3ccd844e97a9718788683d4c7ceaefa6ca0030585b  <= Iff3e149eb4ce60c9f28638248c33ab96208976458886b1735785c2dba298121d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[0] ) begin
                    If53d34fa90e564a24f6e116baa8a7934ec4c51c5f0bce8160f0f389391792fe9  <=  ~I1bc8f647801308e33369cc5f2652781230a588ae772b1e53992f2124c17ad5d9 + 1;
                end else begin
                    If53d34fa90e564a24f6e116baa8a7934ec4c51c5f0bce8160f0f389391792fe9  <= I1bc8f647801308e33369cc5f2652781230a588ae772b1e53992f2124c17ad5d9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[0] ) begin
                    I979c6bc2b8486315e3db6888ef068b88396857d05a62470d4f3c33833cfde130  <=  ~I4e3be7e07012df2e0a3bc90dcb0b4756a778cfcf9192e3722191ba8be32e7e14 + 1;
                end else begin
                    I979c6bc2b8486315e3db6888ef068b88396857d05a62470d4f3c33833cfde130  <= I4e3be7e07012df2e0a3bc90dcb0b4756a778cfcf9192e3722191ba8be32e7e14 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[1] ) begin
                    I1d9a8ff2514f112838c7e4f568303dfcac3f86d94003ec4f1a40a35b79ee8ef6  <=  ~I5c01e607e3f3ba8c06fa54e0ea9fdf0dea25c19c9eb317e51a670199ad40ea90 + 1;
                end else begin
                    I1d9a8ff2514f112838c7e4f568303dfcac3f86d94003ec4f1a40a35b79ee8ef6  <= I5c01e607e3f3ba8c06fa54e0ea9fdf0dea25c19c9eb317e51a670199ad40ea90 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[0] ) begin
                    I8c2fe0c8cb55f09e4dcdbaa3960acfd815764161f53c6234273dffe4558644cf  <=  ~I38fa842b13449763b8db07a9f91ab3479670dbc6043c1b363df6c93f6d7011b5 + 1;
                end else begin
                    I8c2fe0c8cb55f09e4dcdbaa3960acfd815764161f53c6234273dffe4558644cf  <= I38fa842b13449763b8db07a9f91ab3479670dbc6043c1b363df6c93f6d7011b5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[0] ) begin
                    I469f4965961eacfe3dd0cb82fce4905e19e6695d71bec95956e8209d2ae39ba1  <=  ~Ie52aeb4c0ba45662d7f71f542630151f22c1801244258b9c8c20dcaed7f1472e + 1;
                end else begin
                    I469f4965961eacfe3dd0cb82fce4905e19e6695d71bec95956e8209d2ae39ba1  <= Ie52aeb4c0ba45662d7f71f542630151f22c1801244258b9c8c20dcaed7f1472e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[1] ) begin
                    Iea2dd4d33966d53ae739a16876ac2cf04e1d95374a5af68e59a5703dfef2aa79  <=  ~Ie995e639d0338c10aaafa2dd930d57c74442bbde282aefcedcc9ac3b1eeee565 + 1;
                end else begin
                    Iea2dd4d33966d53ae739a16876ac2cf04e1d95374a5af68e59a5703dfef2aa79  <= Ie995e639d0338c10aaafa2dd930d57c74442bbde282aefcedcc9ac3b1eeee565 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[1] ) begin
                    I68ed84b705e3c00d0fb66182d6eeb93f43999532d713f81fab39a36259e0e7da  <=  ~I3b7705f03e900fd64d1b68f0b4036e5ef40c39722a2e6bc8ea6f22f91fb4b044 + 1;
                end else begin
                    I68ed84b705e3c00d0fb66182d6eeb93f43999532d713f81fab39a36259e0e7da  <= I3b7705f03e900fd64d1b68f0b4036e5ef40c39722a2e6bc8ea6f22f91fb4b044 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[0] ) begin
                    I22c3d90c4ad5f41054f9b3dc7ddae143f567182c7fc695c5cd087f126ccdbcf8  <=  ~I4656f355712fef190fb3697699fda1c25bbe9f7577a4d1a95aab55550fd7bfbf + 1;
                end else begin
                    I22c3d90c4ad5f41054f9b3dc7ddae143f567182c7fc695c5cd087f126ccdbcf8  <= I4656f355712fef190fb3697699fda1c25bbe9f7577a4d1a95aab55550fd7bfbf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[2] ) begin
                    I3d6f6b104bd2ffb35ea6782748bb777ec7eceae47ef2e1d18d37d1677d56cb80  <=  ~Ie53b7792c539fa6f2aac95f09dd4a489c9167cf9d6d749f498ab99380c2e694a + 1;
                end else begin
                    I3d6f6b104bd2ffb35ea6782748bb777ec7eceae47ef2e1d18d37d1677d56cb80  <= Ie53b7792c539fa6f2aac95f09dd4a489c9167cf9d6d749f498ab99380c2e694a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[1] ) begin
                    Iceb8741c9680982b02ba9fa2dd76d3b45155ca5f688b70c41d66f3b3690dce42  <=  ~Ie8270cd60cde73d16c5b65134dd393e02f413312f997a0344223cfe05d27985b + 1;
                end else begin
                    Iceb8741c9680982b02ba9fa2dd76d3b45155ca5f688b70c41d66f3b3690dce42  <= Ie8270cd60cde73d16c5b65134dd393e02f413312f997a0344223cfe05d27985b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[2] ) begin
                    I256cb35fd6d4e6c6e1c1a9b42dcbc307f858e5f9525acee9fa7af42c820664f2  <=  ~I53d82131f37765f57bd586de5a55e92a697f63f20f366913802549f9ce658e68 + 1;
                end else begin
                    I256cb35fd6d4e6c6e1c1a9b42dcbc307f858e5f9525acee9fa7af42c820664f2  <= I53d82131f37765f57bd586de5a55e92a697f63f20f366913802549f9ce658e68 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[1] ) begin
                    If0fe01f34db565bf669e2df82579abb4d3629e8bb001bbf874b9b76f8f780a37  <=  ~I289dc39cab39ac30635179b9cd90bd31489a146c8c026138e1a1f9ef7a0ba30c + 1;
                end else begin
                    If0fe01f34db565bf669e2df82579abb4d3629e8bb001bbf874b9b76f8f780a37  <= I289dc39cab39ac30635179b9cd90bd31489a146c8c026138e1a1f9ef7a0ba30c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[1] ) begin
                    I6d58dbbb9b18e4b347b34e548c70a9bc0d819986fb3a6bcc3ff8a67c1fce9c9f  <=  ~I23d6a001aa9c80161e8b305bf34ef8d675247595457a8326a13fd348a02a1539 + 1;
                end else begin
                    I6d58dbbb9b18e4b347b34e548c70a9bc0d819986fb3a6bcc3ff8a67c1fce9c9f  <= I23d6a001aa9c80161e8b305bf34ef8d675247595457a8326a13fd348a02a1539 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[1] ) begin
                    Ic20328b806ccf89387180fe6d88ba762051c6bc2c7f82494129e8c3600108804  <=  ~I15c69e4ab6a25a44e8cb3ae11dfdf0e1dcf71c2cd63add1ab315e1d8a2d2043f + 1;
                end else begin
                    Ic20328b806ccf89387180fe6d88ba762051c6bc2c7f82494129e8c3600108804  <= I15c69e4ab6a25a44e8cb3ae11dfdf0e1dcf71c2cd63add1ab315e1d8a2d2043f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[1] ) begin
                    I8ab86da421b01a03999daa91e41ae95ff58c6bc38566a3deff72633a5ad1cc18  <=  ~I36dcdce4926fb26d7d1b098549754fdfbc3b61a8947394227deedcb51ef1c374 + 1;
                end else begin
                    I8ab86da421b01a03999daa91e41ae95ff58c6bc38566a3deff72633a5ad1cc18  <= I36dcdce4926fb26d7d1b098549754fdfbc3b61a8947394227deedcb51ef1c374 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[0] ) begin
                    I566a76fd27d46125a614f5e0c72dff06a0c1d836c7fe4a2c4086129386b34dde  <=  ~Ic97aaa16a00e936ef8bd742c1c1c14696a72063ec283fcfd02962ffddc327cb5 + 1;
                end else begin
                    I566a76fd27d46125a614f5e0c72dff06a0c1d836c7fe4a2c4086129386b34dde  <= Ic97aaa16a00e936ef8bd742c1c1c14696a72063ec283fcfd02962ffddc327cb5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[2] ) begin
                    I3cca3cf08c967f80e7e255a590bb9c442abc535cd529f7ff304f25d5519dab04  <=  ~Ia28ac0bd59dbf550e8f75ac42fa8618aef3a8323a0e0cd6bc6dccd79c71fe396 + 1;
                end else begin
                    I3cca3cf08c967f80e7e255a590bb9c442abc535cd529f7ff304f25d5519dab04  <= Ia28ac0bd59dbf550e8f75ac42fa8618aef3a8323a0e0cd6bc6dccd79c71fe396 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[1] ) begin
                    I60014273d45dd5019a1b82bdc0a65e44d9a16368d996c8c9ff312fe27e236171  <=  ~I70f499bcd8ce706da16f5d06d481e5197fda5d63b024d9850a34bdaf8f41c2cd + 1;
                end else begin
                    I60014273d45dd5019a1b82bdc0a65e44d9a16368d996c8c9ff312fe27e236171  <= I70f499bcd8ce706da16f5d06d481e5197fda5d63b024d9850a34bdaf8f41c2cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[2] ) begin
                    I53d3de58d6308b770e4a8884447a5f0b92931c8d83c62c86714b6e539b498894  <=  ~Ie7a936ed864922de2eca56a7a648d209cef422443181f89ebbbd6724f5bd0ee4 + 1;
                end else begin
                    I53d3de58d6308b770e4a8884447a5f0b92931c8d83c62c86714b6e539b498894  <= Ie7a936ed864922de2eca56a7a648d209cef422443181f89ebbbd6724f5bd0ee4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[1] ) begin
                    Ie2e727d2073eda2be7642a6a2937cd3c4e553d8bb6ec56d914231b5bfb12405b  <=  ~Ifa54fad7897ca3a5db0d7fdf35cba73823e245f86c54af8a772f1d30f540247c + 1;
                end else begin
                    Ie2e727d2073eda2be7642a6a2937cd3c4e553d8bb6ec56d914231b5bfb12405b  <= Ifa54fad7897ca3a5db0d7fdf35cba73823e245f86c54af8a772f1d30f540247c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[1] ) begin
                    I42968c25ee2870f891f69991ae3ad8bc1c3acde2f8f4d6c0cacc48f562399c37  <=  ~I8c7c890f6f561a9a81130bf7ef4100851c3d86620903cb6b6d648746c0463b46 + 1;
                end else begin
                    I42968c25ee2870f891f69991ae3ad8bc1c3acde2f8f4d6c0cacc48f562399c37  <= I8c7c890f6f561a9a81130bf7ef4100851c3d86620903cb6b6d648746c0463b46 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[1] ) begin
                    I218ab164221d559f1e8bc2a13f06a7593eb4133134762698eec270be5d4c3906  <=  ~I53795a7f407f9dd9d22f6483bbf9efb36313825abbc84c49e1885b01cb2724ed + 1;
                end else begin
                    I218ab164221d559f1e8bc2a13f06a7593eb4133134762698eec270be5d4c3906  <= I53795a7f407f9dd9d22f6483bbf9efb36313825abbc84c49e1885b01cb2724ed ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[1] ) begin
                    If6cd81d168d83d5f6a7ca18051bbbcea5c7a9e017cfffcf72f31f73275c3a4d4  <=  ~I9d28182f6270a0cad620a562c047b449c03bc2036e855d1842707337fbf007eb + 1;
                end else begin
                    If6cd81d168d83d5f6a7ca18051bbbcea5c7a9e017cfffcf72f31f73275c3a4d4  <= I9d28182f6270a0cad620a562c047b449c03bc2036e855d1842707337fbf007eb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[0] ) begin
                    I08240dfbc0f698324c1ffdb8e769016bb8b947fb0b8dbb72839375cdb4cc47e1  <=  ~I2837d4f41e5abdb0abe8c9282938afdd85015263ad60e9a187ee91944f18bd1a + 1;
                end else begin
                    I08240dfbc0f698324c1ffdb8e769016bb8b947fb0b8dbb72839375cdb4cc47e1  <= I2837d4f41e5abdb0abe8c9282938afdd85015263ad60e9a187ee91944f18bd1a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[2] ) begin
                    Ic4839247bb24d460ee6d963d31fc390e8d9d679cd73f058d94ec34a18ceb39c0  <=  ~I832e0057c56a4b0624a8ba7fc95565ff1322ef3b377d21b243c1fa69a9b83982 + 1;
                end else begin
                    Ic4839247bb24d460ee6d963d31fc390e8d9d679cd73f058d94ec34a18ceb39c0  <= I832e0057c56a4b0624a8ba7fc95565ff1322ef3b377d21b243c1fa69a9b83982 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[1] ) begin
                    Ib53bac100fd49f57a5185ff4ad973dfe8eaef6de1937bb32d9246dae9459442b  <=  ~I81243c0fe8b8a3ab03ea4a07b48ae230b9783bc2b49006705893387b2eb0353b + 1;
                end else begin
                    Ib53bac100fd49f57a5185ff4ad973dfe8eaef6de1937bb32d9246dae9459442b  <= I81243c0fe8b8a3ab03ea4a07b48ae230b9783bc2b49006705893387b2eb0353b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[2] ) begin
                    Ife27bd449bf6acad3f06d6e337bfc29c612ba6b3f06927e6f9699ab24d1e836e  <=  ~I53e079434705c9ad3bf3e5cdf3f1d09bd1b0f7742fab2145a089e823e5c28f30 + 1;
                end else begin
                    Ife27bd449bf6acad3f06d6e337bfc29c612ba6b3f06927e6f9699ab24d1e836e  <= I53e079434705c9ad3bf3e5cdf3f1d09bd1b0f7742fab2145a089e823e5c28f30 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[1] ) begin
                    I7d0cbdb63988e88f9f3f69b35029cb2078b97b6cc9008644b2721eda7fb6cfad  <=  ~I77f3f1abf296aafc631f7b3d8bec79228071d4097f2083f70dfee8fa6ca52ba9 + 1;
                end else begin
                    I7d0cbdb63988e88f9f3f69b35029cb2078b97b6cc9008644b2721eda7fb6cfad  <= I77f3f1abf296aafc631f7b3d8bec79228071d4097f2083f70dfee8fa6ca52ba9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[1] ) begin
                    I05bd9a1d7818f4945ddc448149dee571e80dca8b6eba7ab79b17b6f84d3f35f4  <=  ~I1704967bdd23aca028c7fd652f9a0efcc55a31662c9f9b65911b7c1241205d9c + 1;
                end else begin
                    I05bd9a1d7818f4945ddc448149dee571e80dca8b6eba7ab79b17b6f84d3f35f4  <= I1704967bdd23aca028c7fd652f9a0efcc55a31662c9f9b65911b7c1241205d9c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[1] ) begin
                    Ie17e17c22c7215d0482ba310638db13a96c0943216f9ebaf53c0c29c69971b23  <=  ~Ia2313572dea3f44e7ec31d1474ed481064164548d3de394b69a6e99f60561388 + 1;
                end else begin
                    Ie17e17c22c7215d0482ba310638db13a96c0943216f9ebaf53c0c29c69971b23  <= Ia2313572dea3f44e7ec31d1474ed481064164548d3de394b69a6e99f60561388 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[1] ) begin
                    I7ae7cc2f052d37b650c0abeccd841b1b18abb4049c976fbdbab72ea579a5d206  <=  ~Icb8aee17be074ffae08bde14b025127c77773cdf482aa5fade629781c3488e18 + 1;
                end else begin
                    I7ae7cc2f052d37b650c0abeccd841b1b18abb4049c976fbdbab72ea579a5d206  <= Icb8aee17be074ffae08bde14b025127c77773cdf482aa5fade629781c3488e18 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[0] ) begin
                    I989259874d3f12b373358db47fed6245f192edac9e7df00531ea7ba75c360d4c  <=  ~I4b2da3ec326ef0ce2bd1ef54c04f06bb0c9c7fe6f0736613537206d5f5568ff9 + 1;
                end else begin
                    I989259874d3f12b373358db47fed6245f192edac9e7df00531ea7ba75c360d4c  <= I4b2da3ec326ef0ce2bd1ef54c04f06bb0c9c7fe6f0736613537206d5f5568ff9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[2] ) begin
                    Ie873b138e19cd7f7e8afa8bd8f8c4610b65d0fcd647e76d880d25f6fe36c54ef  <=  ~I475e873205aaae01975a2852b3d3d99aeb7ec9aa17759595012bf55fea91ff81 + 1;
                end else begin
                    Ie873b138e19cd7f7e8afa8bd8f8c4610b65d0fcd647e76d880d25f6fe36c54ef  <= I475e873205aaae01975a2852b3d3d99aeb7ec9aa17759595012bf55fea91ff81 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[1] ) begin
                    I4f56f225d6fa40e0469f803c2f72ca27e9c45768ad2af9af9ad10e529e249aa0  <=  ~I9d7892388f5775db1b77de0b60b10ed4f40c44774e1ca7ffc723e5fad503c487 + 1;
                end else begin
                    I4f56f225d6fa40e0469f803c2f72ca27e9c45768ad2af9af9ad10e529e249aa0  <= I9d7892388f5775db1b77de0b60b10ed4f40c44774e1ca7ffc723e5fad503c487 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[2] ) begin
                    Idf239af48228dc01198fdd7240b8282cf247cbc6969403dd994aeac0e5f81898  <=  ~Ib459acc97fee8ddd325d7d8b18d5c339a3c1e03c919c750f88070ec8a4f8a0ad + 1;
                end else begin
                    Idf239af48228dc01198fdd7240b8282cf247cbc6969403dd994aeac0e5f81898  <= Ib459acc97fee8ddd325d7d8b18d5c339a3c1e03c919c750f88070ec8a4f8a0ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[1] ) begin
                    I83ec3e2a8ec621acd2afe475255e144f2158e1941ec685a346b75fc471b9cb76  <=  ~I25711c9c95cd06f19d25d01854fdb8290f4759c9133d1a0c9e88548b886050a1 + 1;
                end else begin
                    I83ec3e2a8ec621acd2afe475255e144f2158e1941ec685a346b75fc471b9cb76  <= I25711c9c95cd06f19d25d01854fdb8290f4759c9133d1a0c9e88548b886050a1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[1] ) begin
                    I6e148041c3612c795f1eb1513a9eba29e0509f02f94971fed189dd9f03d54a4c  <=  ~If9e2ce38db8f4cb30a3748fc7ee1244c98a4ef3c6dc840123405c585f6a867b7 + 1;
                end else begin
                    I6e148041c3612c795f1eb1513a9eba29e0509f02f94971fed189dd9f03d54a4c  <= If9e2ce38db8f4cb30a3748fc7ee1244c98a4ef3c6dc840123405c585f6a867b7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[1] ) begin
                    I5fa628cdc28fdeb96014a4d2c2d06b092136cf2a14a0420bd5d3861b83687413  <=  ~I6b1a6a399505ffa0312c9c79ecca8d63de6c5a1c9f6c0590296cb316c22d114f + 1;
                end else begin
                    I5fa628cdc28fdeb96014a4d2c2d06b092136cf2a14a0420bd5d3861b83687413  <= I6b1a6a399505ffa0312c9c79ecca8d63de6c5a1c9f6c0590296cb316c22d114f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[1] ) begin
                    I533d6897ed500a803f6f6468e36a2a922495b3effbeb405b47ffb7a5f4d82c89  <=  ~I5454f64581fced198aa8ed832feea4c5a3de221d45b8eb42ae5820d82e540931 + 1;
                end else begin
                    I533d6897ed500a803f6f6468e36a2a922495b3effbeb405b47ffb7a5f4d82c89  <= I5454f64581fced198aa8ed832feea4c5a3de221d45b8eb42ae5820d82e540931 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[0] ) begin
                    I06186aec49594899011a9d7bce163a3a43ec094d7c92033df033594ed5eb43ac  <=  ~Ie2235e43965f0eebff14c5c279ef56fc3e4055cc263c20f8d993756e7a5d9b2d + 1;
                end else begin
                    I06186aec49594899011a9d7bce163a3a43ec094d7c92033df033594ed5eb43ac  <= Ie2235e43965f0eebff14c5c279ef56fc3e4055cc263c20f8d993756e7a5d9b2d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[2] ) begin
                    I7ce5fe43a760b5a43815388233952e1bfe5d8b5a7c002f26ae2d462129aad434  <=  ~I72979b4880af333f9e67500779c23973ada097a3cd1e2d4dff0eed1c570f299f + 1;
                end else begin
                    I7ce5fe43a760b5a43815388233952e1bfe5d8b5a7c002f26ae2d462129aad434  <= I72979b4880af333f9e67500779c23973ada097a3cd1e2d4dff0eed1c570f299f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[1] ) begin
                    I8e23f89e84e219d5351bdfd4aab58f61c1cb310cc731164c6e0dd2eac37b07af  <=  ~I4d0c6d6a69f818fe0856050283b987099cd8c7f3c8c22fdc825a01734c4642bc + 1;
                end else begin
                    I8e23f89e84e219d5351bdfd4aab58f61c1cb310cc731164c6e0dd2eac37b07af  <= I4d0c6d6a69f818fe0856050283b987099cd8c7f3c8c22fdc825a01734c4642bc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[2] ) begin
                    Iea2bd90043dd35ae24830a90ed10d12869de66637ab0237a1ad459fa916b57af  <=  ~I811e21f3227b2bc3bd72e9b312edf9bf8e88261543c6bdb1bb09607f49b8206d + 1;
                end else begin
                    Iea2bd90043dd35ae24830a90ed10d12869de66637ab0237a1ad459fa916b57af  <= I811e21f3227b2bc3bd72e9b312edf9bf8e88261543c6bdb1bb09607f49b8206d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[1] ) begin
                    If2b1e365b8ee6d4afa8536f5c2f5c80d31e86ab6729b26795614d75a6a18ef42  <=  ~I4e06a2f339c14dfd77c1d58f78598240d08a7fc156a785a8a3fcae2d2d6d0549 + 1;
                end else begin
                    If2b1e365b8ee6d4afa8536f5c2f5c80d31e86ab6729b26795614d75a6a18ef42  <= I4e06a2f339c14dfd77c1d58f78598240d08a7fc156a785a8a3fcae2d2d6d0549 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[2] ) begin
                    I83c8ad082be8fe1a71adac4f41a3bd7019d2df299d19f8e5a293367e49b04fa5  <=  ~I167bb55e57f960522bce657a28f3a58bb6d82aec339cd46a3e8c4136ee023474 + 1;
                end else begin
                    I83c8ad082be8fe1a71adac4f41a3bd7019d2df299d19f8e5a293367e49b04fa5  <= I167bb55e57f960522bce657a28f3a58bb6d82aec339cd46a3e8c4136ee023474 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[1] ) begin
                    I0b525cae7fe005cf25a07cb0b1486152d726fc74aa55f03480f10af97379953b  <=  ~Ifde56fe010824d9eea62caa160db5bde8de47e31630cd6a8c5e0572df0fa0709 + 1;
                end else begin
                    I0b525cae7fe005cf25a07cb0b1486152d726fc74aa55f03480f10af97379953b  <= Ifde56fe010824d9eea62caa160db5bde8de47e31630cd6a8c5e0572df0fa0709 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[2] ) begin
                    I17eff5960d8d41f0832a48fe9a3ae0dfeef1bfc44b73eff506fe1d3813398d15  <=  ~I1b81ea9b142b222ca4b90724e3c4facaba82a4dea5c9b05c66032b06a459706e + 1;
                end else begin
                    I17eff5960d8d41f0832a48fe9a3ae0dfeef1bfc44b73eff506fe1d3813398d15  <= I1b81ea9b142b222ca4b90724e3c4facaba82a4dea5c9b05c66032b06a459706e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[2] ) begin
                    Iedf1b21de2a0eb04c4a64f9eb34e2b0b3a152d90b1938b61ca45c880eab16ab6  <=  ~I3e9361e7d30732f3e689391f56f9007c32c2368c9eb9d85b933f798babb0da68 + 1;
                end else begin
                    Iedf1b21de2a0eb04c4a64f9eb34e2b0b3a152d90b1938b61ca45c880eab16ab6  <= I3e9361e7d30732f3e689391f56f9007c32c2368c9eb9d85b933f798babb0da68 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[2] ) begin
                    I11855780f53e8711f8eca9370af31f472dffd126c02cfce8154a959f33c68af6  <=  ~I1774935be7ae799801f3b949e3a99707c4b32e7b1538e9f63cd8b940295ea6b1 + 1;
                end else begin
                    I11855780f53e8711f8eca9370af31f472dffd126c02cfce8154a959f33c68af6  <= I1774935be7ae799801f3b949e3a99707c4b32e7b1538e9f63cd8b940295ea6b1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[1] ) begin
                    Ic754ed4f2d29b948b422876f371df4f89b86976e25183ce1b9f664e1a9b19f56  <=  ~Ia4f0bde88d8ea45e325a92c25209a97269d31e2e3999ffe83696236b611de74d + 1;
                end else begin
                    Ic754ed4f2d29b948b422876f371df4f89b86976e25183ce1b9f664e1a9b19f56  <= Ia4f0bde88d8ea45e325a92c25209a97269d31e2e3999ffe83696236b611de74d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[2] ) begin
                    I634dc6f7c843c6e4c63ce6a21b9cd7a386600d1155c0696988403fc1ab790217  <=  ~I30378eb921b9521d10fa2953f99f0f362b986bac12404a78a5f50619fe3b55fd + 1;
                end else begin
                    I634dc6f7c843c6e4c63ce6a21b9cd7a386600d1155c0696988403fc1ab790217  <= I30378eb921b9521d10fa2953f99f0f362b986bac12404a78a5f50619fe3b55fd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[1] ) begin
                    I169d92aaa7eb4f8516e38745955b91d8f6e0ff43cb212186293bb78884282978  <=  ~I972ff0b38d85487454c289292e792035f568f072c33914f87e1f9c981da34370 + 1;
                end else begin
                    I169d92aaa7eb4f8516e38745955b91d8f6e0ff43cb212186293bb78884282978  <= I972ff0b38d85487454c289292e792035f568f072c33914f87e1f9c981da34370 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[2] ) begin
                    I25600d0eb62c066eda0baba4269851387918088406d117377eb8bcc2e080e426  <=  ~I22ad40f4d98f11e2fc7b9a8d56e44092f6e319c4edb2a67c5d9dcacb6a038846 + 1;
                end else begin
                    I25600d0eb62c066eda0baba4269851387918088406d117377eb8bcc2e080e426  <= I22ad40f4d98f11e2fc7b9a8d56e44092f6e319c4edb2a67c5d9dcacb6a038846 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[1] ) begin
                    Icad68e9babee274d9a5b79cf432d9e2a1938e06f51aeb564af6936972b3f8e54  <=  ~If52bfa5da5e6508360b34b20a9607809dc732ad7d40860c8677bb6983d8c30a2 + 1;
                end else begin
                    Icad68e9babee274d9a5b79cf432d9e2a1938e06f51aeb564af6936972b3f8e54  <= If52bfa5da5e6508360b34b20a9607809dc732ad7d40860c8677bb6983d8c30a2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[2] ) begin
                    I09e6d011dacfba2800f9ade6a495076a67e4acc6a944fd649a7c382422e8fa6a  <=  ~I2e9200c7443fa92d38415a8988c0a7ae2366612db06cfc84d9de4faf53d7d1c4 + 1;
                end else begin
                    I09e6d011dacfba2800f9ade6a495076a67e4acc6a944fd649a7c382422e8fa6a  <= I2e9200c7443fa92d38415a8988c0a7ae2366612db06cfc84d9de4faf53d7d1c4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[1] ) begin
                    Idc64cee034c1ee132335ae593844b2c46e3f1b1b2cda8699940df311735a32a0  <=  ~If23a3c0642ef8cb4b2d375a21de5253ad97342b92d29b8b7417bbd9ad0fb2fd5 + 1;
                end else begin
                    Idc64cee034c1ee132335ae593844b2c46e3f1b1b2cda8699940df311735a32a0  <= If23a3c0642ef8cb4b2d375a21de5253ad97342b92d29b8b7417bbd9ad0fb2fd5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[2] ) begin
                    I2f687e6270528a72aa2f9f9cc0a5a6368f8eef358270329cc40b56abc0e4a35e  <=  ~I8b801d7872264ef55cc09008ded93c39bcf86fcd83e472ebc91d27c953520017 + 1;
                end else begin
                    I2f687e6270528a72aa2f9f9cc0a5a6368f8eef358270329cc40b56abc0e4a35e  <= I8b801d7872264ef55cc09008ded93c39bcf86fcd83e472ebc91d27c953520017 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[2] ) begin
                    I5b4ba308b0fc2946fb11b66aa5c24c7b5cb2a21955116b97f3790de65cd2a064  <=  ~I727fdffb518b29e800d3761e94d33c96bf32b4006f248d8eeeb18a035a7c8abe + 1;
                end else begin
                    I5b4ba308b0fc2946fb11b66aa5c24c7b5cb2a21955116b97f3790de65cd2a064  <= I727fdffb518b29e800d3761e94d33c96bf32b4006f248d8eeeb18a035a7c8abe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[2] ) begin
                    I4135dbaf658fb73b41800cd275824d1c9f410ab1b6e555b6c4c8df12f96c5861  <=  ~I4b5a25e13e61b54b754dbb201add03176d432d0c31f3ee1a4086797eec57cbd4 + 1;
                end else begin
                    I4135dbaf658fb73b41800cd275824d1c9f410ab1b6e555b6c4c8df12f96c5861  <= I4b5a25e13e61b54b754dbb201add03176d432d0c31f3ee1a4086797eec57cbd4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[1] ) begin
                    Ia9ea47bb0829c979af002fb7aa0e22072671c2876bcdf79365ff2b3691172149  <=  ~If4413af8c4f8f3dd1f90f00fb5067c95a240f9e3ba7271b134cfda0a1fad603b + 1;
                end else begin
                    Ia9ea47bb0829c979af002fb7aa0e22072671c2876bcdf79365ff2b3691172149  <= If4413af8c4f8f3dd1f90f00fb5067c95a240f9e3ba7271b134cfda0a1fad603b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[2] ) begin
                    Iac9f4a2fa823ae63e73b655020376580991cd4b2b3123204a757afeefe35a10f  <=  ~I0640e35183fc639f884fbb98626d0d54556ba20b2a709c1b4eedad0d3e27ad12 + 1;
                end else begin
                    Iac9f4a2fa823ae63e73b655020376580991cd4b2b3123204a757afeefe35a10f  <= I0640e35183fc639f884fbb98626d0d54556ba20b2a709c1b4eedad0d3e27ad12 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[1] ) begin
                    I737ae96fe290087c8ae686b90b2ac94df2185f7ad8b4252a6ec850278ba5ea9d  <=  ~I79f29e0d9e4930c0e8eab1a5fa373778c2663402943ae843e94dc1d3ac60192a + 1;
                end else begin
                    I737ae96fe290087c8ae686b90b2ac94df2185f7ad8b4252a6ec850278ba5ea9d  <= I79f29e0d9e4930c0e8eab1a5fa373778c2663402943ae843e94dc1d3ac60192a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[2] ) begin
                    I61f7e06790f5516eba113bb79388fb515faa1b3a3bf06598a07f534ce2845618  <=  ~If41e7a25c141c9a83ddd7dbf5bcbb72f579ba7d25231b25ab91ecdd1b8c50af0 + 1;
                end else begin
                    I61f7e06790f5516eba113bb79388fb515faa1b3a3bf06598a07f534ce2845618  <= If41e7a25c141c9a83ddd7dbf5bcbb72f579ba7d25231b25ab91ecdd1b8c50af0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[1] ) begin
                    I16ffb13aa3dfd9da5da39d9b2246d5ab46fd0fdb7c02781abf4d8bd754bbbdf3  <=  ~Iabb9a156ffea98c56dcbde6d29fd606deeb21debc4aa2629e41c035547d5a589 + 1;
                end else begin
                    I16ffb13aa3dfd9da5da39d9b2246d5ab46fd0fdb7c02781abf4d8bd754bbbdf3  <= Iabb9a156ffea98c56dcbde6d29fd606deeb21debc4aa2629e41c035547d5a589 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[2] ) begin
                    I308f551a8479d066b2a4b473206e8f407082cf83b37a376e6b0e1454f7ea2635  <=  ~I496dabb1a4608940824606478478a3050517d422cfb20c53c37523f34aa08a45 + 1;
                end else begin
                    I308f551a8479d066b2a4b473206e8f407082cf83b37a376e6b0e1454f7ea2635  <= I496dabb1a4608940824606478478a3050517d422cfb20c53c37523f34aa08a45 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[1] ) begin
                    I710a57e6c5c8e228325430ba2a5fc32ed9da101d76ccf1d8c9f3397859b39ef3  <=  ~I8bf71b880aa8654933f2008a17308e8366b6f6f22f52091e06364bd10004b891 + 1;
                end else begin
                    I710a57e6c5c8e228325430ba2a5fc32ed9da101d76ccf1d8c9f3397859b39ef3  <= I8bf71b880aa8654933f2008a17308e8366b6f6f22f52091e06364bd10004b891 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[2] ) begin
                    I82772b528a8c156f2932a23a720f8446f3062e9605839897b4652bb2936fca1d  <=  ~I1748e381924bfb743c1257d7830da580af261ef967ffdc1adfafee17c67693aa + 1;
                end else begin
                    I82772b528a8c156f2932a23a720f8446f3062e9605839897b4652bb2936fca1d  <= I1748e381924bfb743c1257d7830da580af261ef967ffdc1adfafee17c67693aa ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[2] ) begin
                    I7c1e9623dc53c8aa8611b46c0375994510a97c4d49d0b091964cbe4671acf1d6  <=  ~I7412e7d6cab6a1cdead2bfb425b79f89328cf155ce5e3b7e8593a4abc457d4aa + 1;
                end else begin
                    I7c1e9623dc53c8aa8611b46c0375994510a97c4d49d0b091964cbe4671acf1d6  <= I7412e7d6cab6a1cdead2bfb425b79f89328cf155ce5e3b7e8593a4abc457d4aa ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[2] ) begin
                    Ie44aa17133d02266160c8fd6f75716f8bc4a3775356cd1ef0f495b13145ba864  <=  ~I39fc2e50c10ec72f5df6ea43b36d62fae7c1c3cbf6f54e921133adc9d8ca884f + 1;
                end else begin
                    Ie44aa17133d02266160c8fd6f75716f8bc4a3775356cd1ef0f495b13145ba864  <= I39fc2e50c10ec72f5df6ea43b36d62fae7c1c3cbf6f54e921133adc9d8ca884f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[1] ) begin
                    I2ef69d9eec4f925b598115d569d2d85a4545871f2ac62635f9b072ba718b595f  <=  ~Ic3be1c01d32bc2fd127d4c4b371fc566b3977bf6f5ecaf4fb7f662f7bdcb36ae + 1;
                end else begin
                    I2ef69d9eec4f925b598115d569d2d85a4545871f2ac62635f9b072ba718b595f  <= Ic3be1c01d32bc2fd127d4c4b371fc566b3977bf6f5ecaf4fb7f662f7bdcb36ae ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[2] ) begin
                    If16869134ec7e59b567e29a1125f0d27eff7a3c612240e25462e2ee84a7e0104  <=  ~Ic9bd71f61271b1ff2f37d36580487d70287b498a51770475819cbfe50d3e48e6 + 1;
                end else begin
                    If16869134ec7e59b567e29a1125f0d27eff7a3c612240e25462e2ee84a7e0104  <= Ic9bd71f61271b1ff2f37d36580487d70287b498a51770475819cbfe50d3e48e6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[1] ) begin
                    I59a4b1b33d114a1b5bdd708e1f856f4bf729c6b86a4064967ca1faf779189164  <=  ~I5217a6046ea279ff9f6f40af49af30f0cdeb374e8c2543da9bb27ce89b08044a + 1;
                end else begin
                    I59a4b1b33d114a1b5bdd708e1f856f4bf729c6b86a4064967ca1faf779189164  <= I5217a6046ea279ff9f6f40af49af30f0cdeb374e8c2543da9bb27ce89b08044a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[2] ) begin
                    I1aadd9b378df1ab58a1b1af097539d1407636833d9c2d8b08c8f70be326fe199  <=  ~Id8c201e2467b255d627059eb66fab4ef48d0c235488dc0f7eb7c350a1d39467e + 1;
                end else begin
                    I1aadd9b378df1ab58a1b1af097539d1407636833d9c2d8b08c8f70be326fe199  <= Id8c201e2467b255d627059eb66fab4ef48d0c235488dc0f7eb7c350a1d39467e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[1] ) begin
                    I1e6d7d9769dc32e1e014951538f1cd1014e9d07b675e6369e88ad5a6fd400787  <=  ~I89de4a293c5da110f92bc9aa9b6ecc790b2fb3e1d282a6373d5ddaff63ef6518 + 1;
                end else begin
                    I1e6d7d9769dc32e1e014951538f1cd1014e9d07b675e6369e88ad5a6fd400787  <= I89de4a293c5da110f92bc9aa9b6ecc790b2fb3e1d282a6373d5ddaff63ef6518 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[2] ) begin
                    Ia428f915c49f84567006696ba3f5c783035325755b4fefcf74d65aaae1f3d3c9  <=  ~I66a3806824b2190f9af7e907d1b4e068fa12560233a9a67bcfc8835373d6d78e + 1;
                end else begin
                    Ia428f915c49f84567006696ba3f5c783035325755b4fefcf74d65aaae1f3d3c9  <= I66a3806824b2190f9af7e907d1b4e068fa12560233a9a67bcfc8835373d6d78e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[1] ) begin
                    I8c8bc477ddc4000dde6459d7cbc4ba665fd4ecd97242d9f9fe97ca6825bb033b  <=  ~Ia7af92f6f7d9e7629ea5a0dc73f90acb4cb2dd8694485491a528df10a2b00aea + 1;
                end else begin
                    I8c8bc477ddc4000dde6459d7cbc4ba665fd4ecd97242d9f9fe97ca6825bb033b  <= Ia7af92f6f7d9e7629ea5a0dc73f90acb4cb2dd8694485491a528df10a2b00aea ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[2] ) begin
                    I44103a07ffcd818c0d9280b96ba08c32f96edc83a981ec9748ed3d6e9c061d62  <=  ~Ia0e8b0cadc0431f58baf6bd1e0fc4ea9babaadf97f47eea75ce07e41cd0e8822 + 1;
                end else begin
                    I44103a07ffcd818c0d9280b96ba08c32f96edc83a981ec9748ed3d6e9c061d62  <= Ia0e8b0cadc0431f58baf6bd1e0fc4ea9babaadf97f47eea75ce07e41cd0e8822 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[2] ) begin
                    Ic0a386f5301913434a3d6aaea1d56d6acb3484fababb7b8831d09563bd8842cb  <=  ~I5c3df19631206eafab24135f4eff9ad9449c874e02c4fa9770d4fc4ede66b3f4 + 1;
                end else begin
                    Ic0a386f5301913434a3d6aaea1d56d6acb3484fababb7b8831d09563bd8842cb  <= I5c3df19631206eafab24135f4eff9ad9449c874e02c4fa9770d4fc4ede66b3f4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[2] ) begin
                    If258ff7e66143201e30b3fd451e1b8e2ec9e46596c2653ec836617c093f28018  <=  ~I74ae8440b495f97712924217bb791b022bbfc59b228632b7f96649f2a2fa053e + 1;
                end else begin
                    If258ff7e66143201e30b3fd451e1b8e2ec9e46596c2653ec836617c093f28018  <= I74ae8440b495f97712924217bb791b022bbfc59b228632b7f96649f2a2fa053e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[1] ) begin
                    Icd8ef17fc44642a3c86a1cb62727eb607e3a4e6d0b021406b9b710ea5c96c06f  <=  ~Ia9c79734a6daa19386ecd68dad6da50274ac40a694cfd496dc40736cb4b33da7 + 1;
                end else begin
                    Icd8ef17fc44642a3c86a1cb62727eb607e3a4e6d0b021406b9b710ea5c96c06f  <= Ia9c79734a6daa19386ecd68dad6da50274ac40a694cfd496dc40736cb4b33da7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[3] ) begin
                    I23ef4f4232fa0d8813a25ddca38a2745fb660c05dbe9ddc2cc33c47d45b3fecf  <=  ~I8d71dedf25220f16c883b67bc750a6e3c8886a6238f13693a22b41345296b0b5 + 1;
                end else begin
                    I23ef4f4232fa0d8813a25ddca38a2745fb660c05dbe9ddc2cc33c47d45b3fecf  <= I8d71dedf25220f16c883b67bc750a6e3c8886a6238f13693a22b41345296b0b5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[3] ) begin
                    Ifb57457918458a6aa9c5df68dbb83243fbc49b3b7037575f43749dfe1bef373a  <=  ~Ieaea96e9413e940b5858f87f12dd18ef7c88b6e84caea900505a50fe657e21e4 + 1;
                end else begin
                    Ifb57457918458a6aa9c5df68dbb83243fbc49b3b7037575f43749dfe1bef373a  <= Ieaea96e9413e940b5858f87f12dd18ef7c88b6e84caea900505a50fe657e21e4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[2] ) begin
                    I9d1a378e4d5703b65f197cb76a1982cc10e0c17654eabcf10d9df091086d8acd  <=  ~Ic8d159cee07bee92aa9171ca69177796c91fa7542a63970a29d785b3cac2f30c + 1;
                end else begin
                    I9d1a378e4d5703b65f197cb76a1982cc10e0c17654eabcf10d9df091086d8acd  <= Ic8d159cee07bee92aa9171ca69177796c91fa7542a63970a29d785b3cac2f30c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c != Iea53e5522afe762dd4185f0262512abbb94b905893974c13e954df5553942b1d[0] ) begin
                    I65cb4f1288affe61a7cd9981878d8519db25d724cecbb80eb3932ccedafcd5bb  <=  ~I4aee30afbdf3dfb74a29ea9bc15aa1b0d200331984b528fade3be76c3249e3f3 + 1;
                end else begin
                    I65cb4f1288affe61a7cd9981878d8519db25d724cecbb80eb3932ccedafcd5bb  <= I4aee30afbdf3dfb74a29ea9bc15aa1b0d200331984b528fade3be76c3249e3f3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[3] ) begin
                    I8ab1772a3bc752331b0bf62069643cadb48bc13bbb06ad3eddc68ac603d73654  <=  ~Ib48fdf999d6a37fee27e903a4581bf51bd4307f83a7a18c3d7fd5ff5e8490a4f + 1;
                end else begin
                    I8ab1772a3bc752331b0bf62069643cadb48bc13bbb06ad3eddc68ac603d73654  <= Ib48fdf999d6a37fee27e903a4581bf51bd4307f83a7a18c3d7fd5ff5e8490a4f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[3] ) begin
                    I8d95c0be0c84d3ee590f8e77065a6ef224e0a75b50aeadea980f9ef4b8d25001  <=  ~Ie581e7d5885d31995c15b699ff1c7f397dd32496d88a5a4c77d1c5bcda532212 + 1;
                end else begin
                    I8d95c0be0c84d3ee590f8e77065a6ef224e0a75b50aeadea980f9ef4b8d25001  <= Ie581e7d5885d31995c15b699ff1c7f397dd32496d88a5a4c77d1c5bcda532212 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[2] ) begin
                    I5df828301af902c72794032c0e55d8e7548c9b2277b2edc77f53796ff8e04804  <=  ~I317cbed94b414a879715617065e78d4ac271816f7f331e5545ba55a46bcd9a5b + 1;
                end else begin
                    I5df828301af902c72794032c0e55d8e7548c9b2277b2edc77f53796ff8e04804  <= I317cbed94b414a879715617065e78d4ac271816f7f331e5545ba55a46bcd9a5b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a != If481e9fd41cf8181d432f397381b8376d9da7ddfba17b52e65e301e74c3b9b0d[0] ) begin
                    I577e642ba232b9a606abfddc4d84ce4354744e2f953da3b285e417dbfc5aef16  <=  ~I76b80ce969069fa14c6d7022d6c072434dfaed48bb2b30aae77035d134019afb + 1;
                end else begin
                    I577e642ba232b9a606abfddc4d84ce4354744e2f953da3b285e417dbfc5aef16  <= I76b80ce969069fa14c6d7022d6c072434dfaed48bb2b30aae77035d134019afb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[3] ) begin
                    Id5055b759fe480d476c4bf08c420a5dafe9e65cb03c6d6991c1d225af0a51d7b  <=  ~I732d56627c4f920af6fac9e623551f6c4c0e5e970b37e4d2f3b0dbc0d2491e29 + 1;
                end else begin
                    Id5055b759fe480d476c4bf08c420a5dafe9e65cb03c6d6991c1d225af0a51d7b  <= I732d56627c4f920af6fac9e623551f6c4c0e5e970b37e4d2f3b0dbc0d2491e29 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[3] ) begin
                    I3a2c9aabb8b064f82bd6f6571bdebdd704abb7526f4977a7b98613f883fdc62a  <=  ~I7c758d1653b4abf515df4c565803d4d5130fad01c8b46a5d447571d0fde55bb8 + 1;
                end else begin
                    I3a2c9aabb8b064f82bd6f6571bdebdd704abb7526f4977a7b98613f883fdc62a  <= I7c758d1653b4abf515df4c565803d4d5130fad01c8b46a5d447571d0fde55bb8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[2] ) begin
                    I0705e6f1954b14f35dd7fa8a64370c2f9e6e39b6e265857e72946815d1f994fe  <=  ~If8ee177b4825244aa2459f76ce3cfe5435b03e72d750c440474a42fee5009643 + 1;
                end else begin
                    I0705e6f1954b14f35dd7fa8a64370c2f9e6e39b6e265857e72946815d1f994fe  <= If8ee177b4825244aa2459f76ce3cfe5435b03e72d750c440474a42fee5009643 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df != If2e4ac195be838db9dd7b062319aba299887896862f1a340013226fa025b18fc[0] ) begin
                    Ic68515eee7d422be9cf8950e48b81d743d5491851d5a117d1f9b70d1d9b55060  <=  ~Ibbffe343259cc28309085b16cf40fb046a0a7c9d5dcef49182ab8ba0a9acbb2a + 1;
                end else begin
                    Ic68515eee7d422be9cf8950e48b81d743d5491851d5a117d1f9b70d1d9b55060  <= Ibbffe343259cc28309085b16cf40fb046a0a7c9d5dcef49182ab8ba0a9acbb2a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[3] ) begin
                    I42d1b7202048c81ca3a8bba0dbbce65501cb7a519fde37085c68d01db7edd635  <=  ~I6ab2cbc5eeb87f6f79360ad8b27bcdf5daad4c85f829eaa00ed855099653be55 + 1;
                end else begin
                    I42d1b7202048c81ca3a8bba0dbbce65501cb7a519fde37085c68d01db7edd635  <= I6ab2cbc5eeb87f6f79360ad8b27bcdf5daad4c85f829eaa00ed855099653be55 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[3] ) begin
                    Ieedfb1902d1f76f95f5f971b578c2440fa5de47dd78e9dc70c35698f813048cb  <=  ~Ib928fe4e8b8da0fa26516833082019238c839091b1fb32c244e57a2aac417273 + 1;
                end else begin
                    Ieedfb1902d1f76f95f5f971b578c2440fa5de47dd78e9dc70c35698f813048cb  <= Ib928fe4e8b8da0fa26516833082019238c839091b1fb32c244e57a2aac417273 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[2] ) begin
                    I3780e5266741d9a9435818f002588f4c44ae518b77a30ede57a3823e1e1e5867  <=  ~Ib59d2666a9c62eea256e01a7e240af2a1c11a86a51058e6ed4034007a881acf1 + 1;
                end else begin
                    I3780e5266741d9a9435818f002588f4c44ae518b77a30ede57a3823e1e1e5867  <= Ib59d2666a9c62eea256e01a7e240af2a1c11a86a51058e6ed4034007a881acf1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a != I40914301545dfe0b6673f76e0dc0d1ab3968ca3b18fe8f4ff63d5623c31bafa7[0] ) begin
                    I0ca47358f982879bb85bd78f6bc19192a5ed8c62214073342b37b040aea331b2  <=  ~I0eccf85cb5b32056038d4f13293549f535d994925067f49a8f1abb6253ed45be + 1;
                end else begin
                    I0ca47358f982879bb85bd78f6bc19192a5ed8c62214073342b37b040aea331b2  <= I0eccf85cb5b32056038d4f13293549f535d994925067f49a8f1abb6253ed45be ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[4] ) begin
                    Id5e78e4ed6db0562ed51d1da1f34242f54def8255088c3a1ccf0221ee8fa153f  <=  ~I5c11c8d23929c41fd11d326b4535976b5e6ad33e2969128e4ec4ccfb0897a22c + 1;
                end else begin
                    Id5e78e4ed6db0562ed51d1da1f34242f54def8255088c3a1ccf0221ee8fa153f  <= I5c11c8d23929c41fd11d326b4535976b5e6ad33e2969128e4ec4ccfb0897a22c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[4] ) begin
                    I88272c473a90efa576a83d0c277090f5814599e5aa192b878cde74215909c46b  <=  ~I7c9db5ef7c22e9722e1811495675725bc9367c52f47417ac0127b2ece6c2b6d5 + 1;
                end else begin
                    I88272c473a90efa576a83d0c277090f5814599e5aa192b878cde74215909c46b  <= I7c9db5ef7c22e9722e1811495675725bc9367c52f47417ac0127b2ece6c2b6d5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[2] ) begin
                    I9a15ed1b2fa413056071c97b4f003717902f38d29805752222c45cbb2cf58109  <=  ~I3d113258d0831ee2590c286fb25bc418e5c1d0033cfa04428717bc3782db11a5 + 1;
                end else begin
                    I9a15ed1b2fa413056071c97b4f003717902f38d29805752222c45cbb2cf58109  <= I3d113258d0831ee2590c286fb25bc418e5c1d0033cfa04428717bc3782db11a5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[2] ) begin
                    I1c7699448a10638886eaa021495d4c7cc378fe1e9b0aafccda001c15484b9419  <=  ~I37fbc80705b247541af9b0468d3bb960bd4b8c1908084a570dc6435714c0f2eb + 1;
                end else begin
                    I1c7699448a10638886eaa021495d4c7cc378fe1e9b0aafccda001c15484b9419  <= I37fbc80705b247541af9b0468d3bb960bd4b8c1908084a570dc6435714c0f2eb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[3] ) begin
                    Iba503643311c9dc3366b9bb843dcc1ee2f0243c4cf78004a660fca224b36c5f2  <=  ~I04ca88712e988bdef397bb8c4e680b6709f92094d54013e6d786aa459174baf5 + 1;
                end else begin
                    Iba503643311c9dc3366b9bb843dcc1ee2f0243c4cf78004a660fca224b36c5f2  <= I04ca88712e988bdef397bb8c4e680b6709f92094d54013e6d786aa459174baf5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 != Idf30e1a70a723113d32f621f0375dd85270da2f7386cff5ef4ff88cfca78b848[0] ) begin
                    I1606027ef88387f2150285b55cef89212359f49ab1a49fb71e457a3dba0c438a  <=  ~Ie8303e1d3cd1305166144c2a9c72da17dc5ff4c6afdb56ea458d2c017a90fcac + 1;
                end else begin
                    I1606027ef88387f2150285b55cef89212359f49ab1a49fb71e457a3dba0c438a  <= Ie8303e1d3cd1305166144c2a9c72da17dc5ff4c6afdb56ea458d2c017a90fcac ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[4] ) begin
                    I4bce49360270b653e45b914c493ca8e5b74beb0b6b85838bb3b54f1f39389fe3  <=  ~I9c8296a684c3ac2e51841b13d88cf64656b4d2f7ac1625a77e0cbed908eb5f8a + 1;
                end else begin
                    I4bce49360270b653e45b914c493ca8e5b74beb0b6b85838bb3b54f1f39389fe3  <= I9c8296a684c3ac2e51841b13d88cf64656b4d2f7ac1625a77e0cbed908eb5f8a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[4] ) begin
                    I91589fd8a2ab91f079bb41631c44926b2c6f83b82448d758d97578c314d0b76c  <=  ~I70b00c7b7fd70b24b225260cda2515d3d5df30d630e9fab4b9f85d810f441649 + 1;
                end else begin
                    I91589fd8a2ab91f079bb41631c44926b2c6f83b82448d758d97578c314d0b76c  <= I70b00c7b7fd70b24b225260cda2515d3d5df30d630e9fab4b9f85d810f441649 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[2] ) begin
                    Iac4172f940fcbc93db2047b26fece588f3fa63ef255ef404beb5e6ea016b2ba3  <=  ~I891eaf9692501bbe1df2bd2f2470be83664f12d9e6211b5523bd7500a1e9fc70 + 1;
                end else begin
                    Iac4172f940fcbc93db2047b26fece588f3fa63ef255ef404beb5e6ea016b2ba3  <= I891eaf9692501bbe1df2bd2f2470be83664f12d9e6211b5523bd7500a1e9fc70 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[2] ) begin
                    I2cb87b14b006ce6a36ee5439eb18a4287c5b9ae79748faee259c0435d0dac81c  <=  ~I807e8a0a095e42d08f8682b77d262989f5440738b49f26eda30b3e70efc7a8e3 + 1;
                end else begin
                    I2cb87b14b006ce6a36ee5439eb18a4287c5b9ae79748faee259c0435d0dac81c  <= I807e8a0a095e42d08f8682b77d262989f5440738b49f26eda30b3e70efc7a8e3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[3] ) begin
                    Id595e96924941a80a6ade8778fcbcef39b07a62fa1d7350fe50182fdae302556  <=  ~I24a328d80a0dd14fa15ad6101cafcef8008c5846474fcd62cfde858dd3d75461 + 1;
                end else begin
                    Id595e96924941a80a6ade8778fcbcef39b07a62fa1d7350fe50182fdae302556  <= I24a328d80a0dd14fa15ad6101cafcef8008c5846474fcd62cfde858dd3d75461 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc != Ic246bc24fb918b7c4a32727a332df57bfb205adc05150ae8d944a77cbdc62822[0] ) begin
                    Ic09f51154140ef91861243d7b35f05961565b368264d44c8fd5d0f85bd0fa213  <=  ~I8273973db378daf42a5ba6dc50c960e8433a2dcb5d17c30f95be6bf89ec0f0b8 + 1;
                end else begin
                    Ic09f51154140ef91861243d7b35f05961565b368264d44c8fd5d0f85bd0fa213  <= I8273973db378daf42a5ba6dc50c960e8433a2dcb5d17c30f95be6bf89ec0f0b8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[4] ) begin
                    I93e543ef3d58bc8bd48a279299dadae1d7f4528c3d09d7106b969e15565d3a15  <=  ~I7ecba0b25a70555c9243a99717462e9f43cacafcbb2ce9b03d34054858620493 + 1;
                end else begin
                    I93e543ef3d58bc8bd48a279299dadae1d7f4528c3d09d7106b969e15565d3a15  <= I7ecba0b25a70555c9243a99717462e9f43cacafcbb2ce9b03d34054858620493 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[4] ) begin
                    I28940d6e8fc5937055f8f50c0d65ac9fd892bdc9f0f2a571808f930c8ad21717  <=  ~Ied4b1e4e915dc6bf15ce0f505d7ac9fa6c5b8cbcc5831cdf270791ea45402c8c + 1;
                end else begin
                    I28940d6e8fc5937055f8f50c0d65ac9fd892bdc9f0f2a571808f930c8ad21717  <= Ied4b1e4e915dc6bf15ce0f505d7ac9fa6c5b8cbcc5831cdf270791ea45402c8c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[2] ) begin
                    I50e7a3df23a8147b9a87cb5e38d44bce7613b2a717d1e3a8bda1171f9522997f  <=  ~I2b2b4121708eceb760e2854c76289daff432118cee2479045dcbd8ebe358e3cc + 1;
                end else begin
                    I50e7a3df23a8147b9a87cb5e38d44bce7613b2a717d1e3a8bda1171f9522997f  <= I2b2b4121708eceb760e2854c76289daff432118cee2479045dcbd8ebe358e3cc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[2] ) begin
                    I54da11ab334a3942047eb5953935aedd00ef1a24bb5361fba51504632ae61831  <=  ~I8eba7f46df1f21311e46e2657b38d61800060add0c96dccfa9c45fae66711d7d + 1;
                end else begin
                    I54da11ab334a3942047eb5953935aedd00ef1a24bb5361fba51504632ae61831  <= I8eba7f46df1f21311e46e2657b38d61800060add0c96dccfa9c45fae66711d7d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[3] ) begin
                    I3f9e2f1be98a5d14a8b79b252e9b5a2b3a09304f27a3526a4a66b365b682787c  <=  ~I587e2742d73f804efba3b90efacfca020ee8a5e13c2a490ec60ac494be39a275 + 1;
                end else begin
                    I3f9e2f1be98a5d14a8b79b252e9b5a2b3a09304f27a3526a4a66b365b682787c  <= I587e2742d73f804efba3b90efacfca020ee8a5e13c2a490ec60ac494be39a275 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 != I6cac9957a16e7cfa8a125b40d8ce42cb7f502078a791b177d9bbe9589b612426[0] ) begin
                    Ie28425115106f4b2405fad6fb2994a76e64dfa60e7bc165f46ae67411932a1cf  <=  ~Ic4766de4b982a051c7546be035a94bb07bc822061d5bd46d9a4070d026b7a593 + 1;
                end else begin
                    Ie28425115106f4b2405fad6fb2994a76e64dfa60e7bc165f46ae67411932a1cf  <= Ic4766de4b982a051c7546be035a94bb07bc822061d5bd46d9a4070d026b7a593 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[4] ) begin
                    I07bdf8f629cfc9c094023be167a717880dc3a42099b01bffb431036521cd6019  <=  ~I5ce28b3e49d61224902a9c1f675a4032351731bd0d14cf3bcab007b30d7e5c22 + 1;
                end else begin
                    I07bdf8f629cfc9c094023be167a717880dc3a42099b01bffb431036521cd6019  <= I5ce28b3e49d61224902a9c1f675a4032351731bd0d14cf3bcab007b30d7e5c22 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[4] ) begin
                    I52f4d169be660862052b60924958cc9a0eb99b1454608fc48d47192452f8b390  <=  ~I07afa69acae532add7b503ba1bf357b95ab120399bc63d32e65af6f61a369f15 + 1;
                end else begin
                    I52f4d169be660862052b60924958cc9a0eb99b1454608fc48d47192452f8b390  <= I07afa69acae532add7b503ba1bf357b95ab120399bc63d32e65af6f61a369f15 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[2] ) begin
                    I15b5266ec781a5ae11540d23bf8b1a0b2eb45d94ab6f367a872885ff3207d5a9  <=  ~I4c0f888abd9ba96ae660c5a3f6e9c627c5775611d7a2956fa3049c5574fde7df + 1;
                end else begin
                    I15b5266ec781a5ae11540d23bf8b1a0b2eb45d94ab6f367a872885ff3207d5a9  <= I4c0f888abd9ba96ae660c5a3f6e9c627c5775611d7a2956fa3049c5574fde7df ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[2] ) begin
                    I3df4fc0f2f099890a34d7b376328da6460d429e2516a5f8fd1aee5a8fee835df  <=  ~I4bb74c7a5d5fa7f8a3bcc33e4aac51ace977350ac258b3af687b215c37407b49 + 1;
                end else begin
                    I3df4fc0f2f099890a34d7b376328da6460d429e2516a5f8fd1aee5a8fee835df  <= I4bb74c7a5d5fa7f8a3bcc33e4aac51ace977350ac258b3af687b215c37407b49 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[3] ) begin
                    I360ab21cba3dfd419f0ca83f85d9633b918c3d24a00214399b0465d7106466ad  <=  ~Ia781a129677ad67c301dedf105bd58147a815283dd2c06d65ca7ada0aca7cc7e + 1;
                end else begin
                    I360ab21cba3dfd419f0ca83f85d9633b918c3d24a00214399b0465d7106466ad  <= Ia781a129677ad67c301dedf105bd58147a815283dd2c06d65ca7ada0aca7cc7e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 != Iee4ad1e7709a56d53cd8b97f587f1f791fb88bf278fcfef32a29fa05247ca13d[0] ) begin
                    I64862889bfd7d2a15503bc07af594be59cbaa8758863f78311d6f15ecadcc99f  <=  ~Ieff7f5ac404485dc7719d026c898a08cddf9eac3289347c09da180a04400da13 + 1;
                end else begin
                    I64862889bfd7d2a15503bc07af594be59cbaa8758863f78311d6f15ecadcc99f  <= Ieff7f5ac404485dc7719d026c898a08cddf9eac3289347c09da180a04400da13 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[5] ) begin
                    I17cdc222663e370d6ef2539ad03c45a7949d9606583c17568a24c528a3e8c12f  <=  ~Idbea312fceb0d3b89f626dc27620dc564adf927f2587857f0c80926c0f323433 + 1;
                end else begin
                    I17cdc222663e370d6ef2539ad03c45a7949d9606583c17568a24c528a3e8c12f  <= Idbea312fceb0d3b89f626dc27620dc564adf927f2587857f0c80926c0f323433 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[3] ) begin
                    I3d6bb14416567aa7b8883b3d1778b55c251a22ed42b09bb3cbae6a5210cf11f0  <=  ~Id1537778668b48b3115e7b1a3cde430a348b515e592a110c520b33226ecf7f47 + 1;
                end else begin
                    I3d6bb14416567aa7b8883b3d1778b55c251a22ed42b09bb3cbae6a5210cf11f0  <= Id1537778668b48b3115e7b1a3cde430a348b515e592a110c520b33226ecf7f47 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[3] ) begin
                    Ide2ca364c5742f786e5408980fbe12322ebcc2920fd99ed322112d3623d9e372  <=  ~I4d749601335050fe4f61b7b9280c1f83ae58f99216ee191f039f6b94b185e74c + 1;
                end else begin
                    Ide2ca364c5742f786e5408980fbe12322ebcc2920fd99ed322112d3623d9e372  <= I4d749601335050fe4f61b7b9280c1f83ae58f99216ee191f039f6b94b185e74c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[3] ) begin
                    Ibe3e6de02f0c30287dd89b07be5254ff70d9683389574d02f1423e792bd2d534  <=  ~I2a445ed5096a1929dc2ef74b28f3243c9e05c70b4e0aed9baedfe94c28d8e4ad + 1;
                end else begin
                    Ibe3e6de02f0c30287dd89b07be5254ff70d9683389574d02f1423e792bd2d534  <= I2a445ed5096a1929dc2ef74b28f3243c9e05c70b4e0aed9baedfe94c28d8e4ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[4] ) begin
                    I2c061ca6ba4299d676b5c6f1e1cc920bc1104e7ac730d207949b952d1a98300f  <=  ~Iae58883a74ef0111e20be8cc9df222d4e0e213d390b08244a5361328ba38895f + 1;
                end else begin
                    I2c061ca6ba4299d676b5c6f1e1cc920bc1104e7ac730d207949b952d1a98300f  <= Iae58883a74ef0111e20be8cc9df222d4e0e213d390b08244a5361328ba38895f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 != I16a4499c48e5c24fd8a6d49ec3bf63c20c85f440c0c897cdb840e9f28fa2e68a[0] ) begin
                    Ied4424f3e85f3fb92f4e40bc63909f4e77698a18a1d0ee651e54e4de06ee330f  <=  ~Ibd5a78278d93327ec1527d2329cb8bdc601611fa5ee53fc37e64259d6bc217a2 + 1;
                end else begin
                    Ied4424f3e85f3fb92f4e40bc63909f4e77698a18a1d0ee651e54e4de06ee330f  <= Ibd5a78278d93327ec1527d2329cb8bdc601611fa5ee53fc37e64259d6bc217a2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[5] ) begin
                    Ibb4ff9ffdb2771ff640bf958798f8447a0dbcf15ed0ef9f82068826ec621de77  <=  ~Id1f021d678d21318bd8881474b337f0b540c16dc97a33c4fc3abc12bb662f4a5 + 1;
                end else begin
                    Ibb4ff9ffdb2771ff640bf958798f8447a0dbcf15ed0ef9f82068826ec621de77  <= Id1f021d678d21318bd8881474b337f0b540c16dc97a33c4fc3abc12bb662f4a5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[3] ) begin
                    I5c1a09aa19ef4bb254881dd92543acf840270aa36ad4e0f5f63a6182a4c93a1d  <=  ~Id4d52f3a7303153d65a86d328d1e7e5dcdd602d284aba3e104ee0528d9b1d465 + 1;
                end else begin
                    I5c1a09aa19ef4bb254881dd92543acf840270aa36ad4e0f5f63a6182a4c93a1d  <= Id4d52f3a7303153d65a86d328d1e7e5dcdd602d284aba3e104ee0528d9b1d465 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[3] ) begin
                    Ib1b15c9e15e963cc4f2e9caa1b6b132e338947224b705b51ebe710d7e0f661d7  <=  ~I608fc1c1a500a0fd76e9a326afc6c5a26d1cd78f1b150d970f5ca74d1d7a3193 + 1;
                end else begin
                    Ib1b15c9e15e963cc4f2e9caa1b6b132e338947224b705b51ebe710d7e0f661d7  <= I608fc1c1a500a0fd76e9a326afc6c5a26d1cd78f1b150d970f5ca74d1d7a3193 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[3] ) begin
                    I005ecc3a38317079c7bc5008817e11017c33671f77364ad9a07d0eff1e0ebf0b  <=  ~I7b2d4fe3f2c703eace8068da2810bc7bc190900ec3959bfc4a396e72ef5a8200 + 1;
                end else begin
                    I005ecc3a38317079c7bc5008817e11017c33671f77364ad9a07d0eff1e0ebf0b  <= I7b2d4fe3f2c703eace8068da2810bc7bc190900ec3959bfc4a396e72ef5a8200 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[4] ) begin
                    I05806fb5d45e4d6f569c12116644b625b7ba071eb052ab97525f06fca03dd88b  <=  ~I72d8c9fea747adec725ada83bdebc85126870df2cd2cb9f88d2d043635bfdd84 + 1;
                end else begin
                    I05806fb5d45e4d6f569c12116644b625b7ba071eb052ab97525f06fca03dd88b  <= I72d8c9fea747adec725ada83bdebc85126870df2cd2cb9f88d2d043635bfdd84 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 != Ibed209db0bc502e3fceb4ab86ac20a2ebf87c43391a546d592e5aa32709aa8bd[0] ) begin
                    I6c850d46af2f31f4e3d31c3fd2b2d9c7471ccf817b452a4fa2602485f5e7f164  <=  ~I4f237165ee7800d1fd20968d90afd5a858b8ae73675c1a03b67be17159247ffa + 1;
                end else begin
                    I6c850d46af2f31f4e3d31c3fd2b2d9c7471ccf817b452a4fa2602485f5e7f164  <= I4f237165ee7800d1fd20968d90afd5a858b8ae73675c1a03b67be17159247ffa ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[5] ) begin
                    Ib6ff050679c6366efde7b9809fcf42051f107c18863bcea79d41b5fee0603e9c  <=  ~I333abb8de54c2cdc50519fe091024d9862592e0191ef4acb0b6e1b7c45701234 + 1;
                end else begin
                    Ib6ff050679c6366efde7b9809fcf42051f107c18863bcea79d41b5fee0603e9c  <= I333abb8de54c2cdc50519fe091024d9862592e0191ef4acb0b6e1b7c45701234 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[3] ) begin
                    I6a10084ceb62d383dbc5871a208fc087b23de418b2c780813ae950bf4e594c96  <=  ~I6ef7e70fed5f181598201b2c2c0002f1251010c752be38c1f229c337e4a66428 + 1;
                end else begin
                    I6a10084ceb62d383dbc5871a208fc087b23de418b2c780813ae950bf4e594c96  <= I6ef7e70fed5f181598201b2c2c0002f1251010c752be38c1f229c337e4a66428 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[3] ) begin
                    I45b03b0185f9efbc11c707a64fda9203cc82ec2fbaee7ff34610c74d7cc1132b  <=  ~I75665f397a59da51376855f9b737164887c48da916cdadc4b4d1605f3d8e4071 + 1;
                end else begin
                    I45b03b0185f9efbc11c707a64fda9203cc82ec2fbaee7ff34610c74d7cc1132b  <= I75665f397a59da51376855f9b737164887c48da916cdadc4b4d1605f3d8e4071 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[3] ) begin
                    I1b5d096081c0190c0ce6a674de1afee9ccd766a9cfab0637a0aec33199061bbf  <=  ~Ie81e5c2a20cacfd646fdc8795e265386030f32624e917b5877a38d9790ed93be + 1;
                end else begin
                    I1b5d096081c0190c0ce6a674de1afee9ccd766a9cfab0637a0aec33199061bbf  <= Ie81e5c2a20cacfd646fdc8795e265386030f32624e917b5877a38d9790ed93be ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[4] ) begin
                    Iefbb3d08b0b2fc51d2f6b60b25b8143f3f88a705e770396e2f6d050632ded97e  <=  ~I9760a21471e149d0c56a22ba9a49f377439bba25562cdba484b355531562bd05 + 1;
                end else begin
                    Iefbb3d08b0b2fc51d2f6b60b25b8143f3f88a705e770396e2f6d050632ded97e  <= I9760a21471e149d0c56a22ba9a49f377439bba25562cdba484b355531562bd05 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 != I05dc9e8db597a2123632b2934d864ae64cab5192401d8f66ebebd95618590ba2[0] ) begin
                    I1a1a9f7ee74e17c4a0d7064ca9fae938002b1b685f3cb6309569081b0d971aed  <=  ~Ie9ad099032e87edfcc146b2b8fc401eb78cd1c370d99a7d87b96cffcb2bace7f + 1;
                end else begin
                    I1a1a9f7ee74e17c4a0d7064ca9fae938002b1b685f3cb6309569081b0d971aed  <= Ie9ad099032e87edfcc146b2b8fc401eb78cd1c370d99a7d87b96cffcb2bace7f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[5] ) begin
                    Ifaa925832248fd0e2f5841096d9618c2fdaa3c63a3130b57f493782f96473088  <=  ~I42d22931f7defa6032679880bb907c668d62e4c65343d359f7ee0679bb098ef2 + 1;
                end else begin
                    Ifaa925832248fd0e2f5841096d9618c2fdaa3c63a3130b57f493782f96473088  <= I42d22931f7defa6032679880bb907c668d62e4c65343d359f7ee0679bb098ef2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[3] ) begin
                    I0e9a7c6c53b89ca2685615c270e8ef3d3f51fad8619953972e1037edfe633834  <=  ~I5d35fcce50496260be81878d7799638cbce05d2afe98817fe9c53a675ee5f98d + 1;
                end else begin
                    I0e9a7c6c53b89ca2685615c270e8ef3d3f51fad8619953972e1037edfe633834  <= I5d35fcce50496260be81878d7799638cbce05d2afe98817fe9c53a675ee5f98d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[3] ) begin
                    Ife00518e7b24a5de694b56a32211898b3c23d2dbd2df91a4197216c23fb5aa7b  <=  ~I0876112eaaac7d4bd5dda75039d334a15e6d500f29e0c471e8d6dd0ba6cf70e9 + 1;
                end else begin
                    Ife00518e7b24a5de694b56a32211898b3c23d2dbd2df91a4197216c23fb5aa7b  <= I0876112eaaac7d4bd5dda75039d334a15e6d500f29e0c471e8d6dd0ba6cf70e9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[3] ) begin
                    Ia8a4fca33add1c3c58b04eafe9d023751882f409c5d2905f77aae3fef8c2b008  <=  ~I612926c7fd5a7811c91d55336a1ea5a427e4c28826227d05d2e08d501bb032d0 + 1;
                end else begin
                    Ia8a4fca33add1c3c58b04eafe9d023751882f409c5d2905f77aae3fef8c2b008  <= I612926c7fd5a7811c91d55336a1ea5a427e4c28826227d05d2e08d501bb032d0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[4] ) begin
                    I134dfd9d579ba8b2d72bf1c47119a086fcfb6b7d591cc2c5558e451f57636d0c  <=  ~I4075a88832d68ad5005c73387153538516b97eb30d8d1bfc9f3d205cf338e042 + 1;
                end else begin
                    I134dfd9d579ba8b2d72bf1c47119a086fcfb6b7d591cc2c5558e451f57636d0c  <= I4075a88832d68ad5005c73387153538516b97eb30d8d1bfc9f3d205cf338e042 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d != Ib309786164a7d646c17533008b3aaf0fd86eda3c5ee167efc2080ef5b26a9ddf[0] ) begin
                    Ib5929b32be13a8436b74dadded1f26d3742e1424b6025d1eacda112bf4749a15  <=  ~I4471c46046bb6606ad97bff8b36a4a9c1643c861791e8b3bf97a41e8cb385220 + 1;
                end else begin
                    Ib5929b32be13a8436b74dadded1f26d3742e1424b6025d1eacda112bf4749a15  <= I4471c46046bb6606ad97bff8b36a4a9c1643c861791e8b3bf97a41e8cb385220 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[5] ) begin
                    Ia3e877a9f66cb7582b125e56b7c3f79601eb8e700f54e14f967a4d9df9b5725d  <=  ~Iee30715a934f261b8e1fb4814e196f3307e095ec0dbfcb10ac1fcaa1d1d16372 + 1;
                end else begin
                    Ia3e877a9f66cb7582b125e56b7c3f79601eb8e700f54e14f967a4d9df9b5725d  <= Iee30715a934f261b8e1fb4814e196f3307e095ec0dbfcb10ac1fcaa1d1d16372 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[4] ) begin
                    Ib99b447a19aa10415461faaa8d8026b0073582bd078930f2cdf0f531259d9c50  <=  ~I8b323499e4c61f57b164a287da64b2f1c933376dc7ec202d666ce57ccffc139f + 1;
                end else begin
                    Ib99b447a19aa10415461faaa8d8026b0073582bd078930f2cdf0f531259d9c50  <= I8b323499e4c61f57b164a287da64b2f1c933376dc7ec202d666ce57ccffc139f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[4] ) begin
                    Ica9ef16b19711ccdfe32e34eed347b590635f1ba7983272eb02f980f80642254  <=  ~Ic936076da3dcc6a7f335b0d3b428e8b01cfeb9240df6dd50bcfb2188cc37ae8c + 1;
                end else begin
                    Ica9ef16b19711ccdfe32e34eed347b590635f1ba7983272eb02f980f80642254  <= Ic936076da3dcc6a7f335b0d3b428e8b01cfeb9240df6dd50bcfb2188cc37ae8c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[5] ) begin
                    Ib2630bec8f9f78489ca6cfe0bf25746b720aa422b9d529d67d6dde2d045d9c3c  <=  ~I1cbbfb485fecaa90d26f81a89b89c0d778558fbc218268369c32c33117c33468 + 1;
                end else begin
                    Ib2630bec8f9f78489ca6cfe0bf25746b720aa422b9d529d67d6dde2d045d9c3c  <= I1cbbfb485fecaa90d26f81a89b89c0d778558fbc218268369c32c33117c33468 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[2] ) begin
                    Id7310932ca8964fd49adc052220c04855b028e29fb7a48521a36e2dbe1d6d5f4  <=  ~I5bd88b9b16b4fbeeecae426d343179b982f46fe09abc37e1db23e03a43157b89 + 1;
                end else begin
                    Id7310932ca8964fd49adc052220c04855b028e29fb7a48521a36e2dbe1d6d5f4  <= I5bd88b9b16b4fbeeecae426d343179b982f46fe09abc37e1db23e03a43157b89 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 != Id9bbd0f5c16ba0ffae6a0e5304e1726b97df06f06feaccbb1bbcaf0e01be3823[0] ) begin
                    Ibcb7809e1db6cb82ba62be017c5b8685cb6f988f85a0d29ce2459f6ac80498dd  <=  ~Ia5fcf505c93f7902d4ed6f1877bf51599e910bbcc6002e122623c389e72e2600 + 1;
                end else begin
                    Ibcb7809e1db6cb82ba62be017c5b8685cb6f988f85a0d29ce2459f6ac80498dd  <= Ia5fcf505c93f7902d4ed6f1877bf51599e910bbcc6002e122623c389e72e2600 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[5] ) begin
                    Ic20b5a20229313d70c01a5f53e13e96095c1d8695144668e66efdc81efdd8374  <=  ~Ib2ed8f97504f1f2331d11107b05d538282eba6248d7d8fc3c9ccbb4a0cfd7e70 + 1;
                end else begin
                    Ic20b5a20229313d70c01a5f53e13e96095c1d8695144668e66efdc81efdd8374  <= Ib2ed8f97504f1f2331d11107b05d538282eba6248d7d8fc3c9ccbb4a0cfd7e70 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[4] ) begin
                    I54b0a17c9919d856bb3ed7cbbd8e42fd4ffa33ce8c32d45e4be1e28b71426ee5  <=  ~Ia2d0125fd752a306fa45115b7d888f2eb705d6f14d3e5d4f5191024ed7b1f746 + 1;
                end else begin
                    I54b0a17c9919d856bb3ed7cbbd8e42fd4ffa33ce8c32d45e4be1e28b71426ee5  <= Ia2d0125fd752a306fa45115b7d888f2eb705d6f14d3e5d4f5191024ed7b1f746 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[4] ) begin
                    I6024b75d70e3da7df4e532e712df56a8bed06352ba0a545ec355f59473929d41  <=  ~If45da818944a7fc1d4baf55234b4a8299f0513f6db7e1e8cd87e7b57f72eb817 + 1;
                end else begin
                    I6024b75d70e3da7df4e532e712df56a8bed06352ba0a545ec355f59473929d41  <= If45da818944a7fc1d4baf55234b4a8299f0513f6db7e1e8cd87e7b57f72eb817 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[5] ) begin
                    I71c3a88492c33461f93d43680f11eae8ef3e9402a4b931c5d31f959a2f8c147e  <=  ~I18d435d55c2e6ef05cdc85c7c5f1fc2e74307ca98333e485f5fcb8eb038dc3f1 + 1;
                end else begin
                    I71c3a88492c33461f93d43680f11eae8ef3e9402a4b931c5d31f959a2f8c147e  <= I18d435d55c2e6ef05cdc85c7c5f1fc2e74307ca98333e485f5fcb8eb038dc3f1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[2] ) begin
                    I58df4f7ee4282cdb7bb80c9f1d907ff37590b1db22994f3a07b521132ab80087  <=  ~I6b9155f4e226a633f272039c862d58cbce7e31a597a37e1be49eb81b0b72cf47 + 1;
                end else begin
                    I58df4f7ee4282cdb7bb80c9f1d907ff37590b1db22994f3a07b521132ab80087  <= I6b9155f4e226a633f272039c862d58cbce7e31a597a37e1be49eb81b0b72cf47 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d != I4294b001f220e009c2a65fbf8b36ce1d8961c317ae8ded31cbe5aa288191e009[0] ) begin
                    Idb971d0017094cf8b28e639623f85e6e5fc2c03a1da1e19a1ef87b959fe8e1cf  <=  ~Ie7dce49639675176aa767ea6d5b2171e0c72deebe4e007b620860a1f8b177060 + 1;
                end else begin
                    Idb971d0017094cf8b28e639623f85e6e5fc2c03a1da1e19a1ef87b959fe8e1cf  <= Ie7dce49639675176aa767ea6d5b2171e0c72deebe4e007b620860a1f8b177060 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[5] ) begin
                    Ifbf3cda7e0639ad343a64c5b3d2f45017f1d280bf72c96520cbf272104c90ad9  <=  ~I8043c8446ed3aac742a14c3df20420bdd5f0e6561e15c32f4045e2ce8b6f3330 + 1;
                end else begin
                    Ifbf3cda7e0639ad343a64c5b3d2f45017f1d280bf72c96520cbf272104c90ad9  <= I8043c8446ed3aac742a14c3df20420bdd5f0e6561e15c32f4045e2ce8b6f3330 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[4] ) begin
                    I9afcfde9391d485e865b08f9b8ff69cc2ecaace5f5e26e27b7e1775b625722c0  <=  ~Ieb807bb8e9746d06de25556b579e51494e760b3a4312caa4862cbf2776acbccb + 1;
                end else begin
                    I9afcfde9391d485e865b08f9b8ff69cc2ecaace5f5e26e27b7e1775b625722c0  <= Ieb807bb8e9746d06de25556b579e51494e760b3a4312caa4862cbf2776acbccb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[4] ) begin
                    Id364040d3b9f1ebf34ae3fdf7465d955b49d7a2f4709219f76229766d6df98a4  <=  ~Ie1f84176002d4791b93729913c6021f1ffd76c58ad11593dc088cbcf2e4bc4c9 + 1;
                end else begin
                    Id364040d3b9f1ebf34ae3fdf7465d955b49d7a2f4709219f76229766d6df98a4  <= Ie1f84176002d4791b93729913c6021f1ffd76c58ad11593dc088cbcf2e4bc4c9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[5] ) begin
                    I5f4870fc880aac0f84130a26e3cd493954ea49eb3804dd17a91b2ba1cea599f3  <=  ~If56795023544f4a2942b0910b389ee77a220fffaf45786cb20c1806f3d76f76a + 1;
                end else begin
                    I5f4870fc880aac0f84130a26e3cd493954ea49eb3804dd17a91b2ba1cea599f3  <= If56795023544f4a2942b0910b389ee77a220fffaf45786cb20c1806f3d76f76a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[2] ) begin
                    If8cefdab8d831c3db83e1ef615ca534f34c58b9903520c7741cafbc84e28d207  <=  ~Ic9d92acd0f4cc0aa5cf4bc5a5f14bb848cb4267dd6aec78011f70039bf4f7c8c + 1;
                end else begin
                    If8cefdab8d831c3db83e1ef615ca534f34c58b9903520c7741cafbc84e28d207  <= Ic9d92acd0f4cc0aa5cf4bc5a5f14bb848cb4267dd6aec78011f70039bf4f7c8c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 != Id1fe66d1340965020f513e73a4f77d18f4703c194c3954d40a7f1bc37fc1342b[0] ) begin
                    I89373d12365deb440d5337a2586fcdab81347ca28ff6f261a12e35a235bd23c6  <=  ~I83b87ecce5b21302ac79a58afdd995b617634440666c2a50df5ba1868c7f81c2 + 1;
                end else begin
                    I89373d12365deb440d5337a2586fcdab81347ca28ff6f261a12e35a235bd23c6  <= I83b87ecce5b21302ac79a58afdd995b617634440666c2a50df5ba1868c7f81c2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[5] ) begin
                    Iade009d6c5b9e00f5459c53b0c254dda356081e6965366db7b7ac42a992e3ae7  <=  ~Ida44179080ae7121a94fa6ddc8d15e57d73d73f15c2007f200eb205bd6c0c63f + 1;
                end else begin
                    Iade009d6c5b9e00f5459c53b0c254dda356081e6965366db7b7ac42a992e3ae7  <= Ida44179080ae7121a94fa6ddc8d15e57d73d73f15c2007f200eb205bd6c0c63f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[4] ) begin
                    I63f5ecb10fc3ed9bd8bf79403afed8ab1a70600ceb1e755de0d44af98495ea88  <=  ~I0708b20a51af5c02051540c2de37aeeca5959bd958280e953a9cdf18c324d905 + 1;
                end else begin
                    I63f5ecb10fc3ed9bd8bf79403afed8ab1a70600ceb1e755de0d44af98495ea88  <= I0708b20a51af5c02051540c2de37aeeca5959bd958280e953a9cdf18c324d905 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[4] ) begin
                    I3097f16921e899a99f2a2b013a3f6d339ac9672fa5e17655ceba4de2d506e151  <=  ~I25510ca31a420de3078e0615a3a9f602e7a6f8698e6a79cb0d2688aa63f8e7cd + 1;
                end else begin
                    I3097f16921e899a99f2a2b013a3f6d339ac9672fa5e17655ceba4de2d506e151  <= I25510ca31a420de3078e0615a3a9f602e7a6f8698e6a79cb0d2688aa63f8e7cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[5] ) begin
                    Ief44fc6df0864dd0766877e0d673847250f53ab137cd9029916ab7149446f9c2  <=  ~Ief493235efee1fdb4705ae4a1a0244c57346ff2b56b269552c6b5d64595056ca + 1;
                end else begin
                    Ief44fc6df0864dd0766877e0d673847250f53ab137cd9029916ab7149446f9c2  <= Ief493235efee1fdb4705ae4a1a0244c57346ff2b56b269552c6b5d64595056ca ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[2] ) begin
                    I2a3d1a32b282fd624497621815c6ff85c904f5f3fb50f18cf345c5a5d7a557ef  <=  ~I0a5ffd7c103836e4867f6819fab3096c582f2ce1db2c303bfebf50104b7d496b + 1;
                end else begin
                    I2a3d1a32b282fd624497621815c6ff85c904f5f3fb50f18cf345c5a5d7a557ef  <= I0a5ffd7c103836e4867f6819fab3096c582f2ce1db2c303bfebf50104b7d496b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 != Ie95c9af987f352eca30c8546d306af7cdada8d2a8037200d303e6afbd5a4f448[0] ) begin
                    Ib8f9b76d6cf7a74f0d437f634ce888096a0d6d81d66dc6c60b62a60006b661e9  <=  ~Ife97a26fdf22e53aaf139436dd732d1fc8cd6cb4957269b6d0666495a0873c4f + 1;
                end else begin
                    Ib8f9b76d6cf7a74f0d437f634ce888096a0d6d81d66dc6c60b62a60006b661e9  <= Ife97a26fdf22e53aaf139436dd732d1fc8cd6cb4957269b6d0666495a0873c4f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[6] ) begin
                    I2c22aed0ed8abb0cb8906a35a4d44cfd7cc68b2924e474680a2eb6cf7caf5582  <=  ~I2bb55e3fbb0c342fd0434fbb00b85eae3c5f4075979e290f3d22673c392e3a60 + 1;
                end else begin
                    I2c22aed0ed8abb0cb8906a35a4d44cfd7cc68b2924e474680a2eb6cf7caf5582  <= I2bb55e3fbb0c342fd0434fbb00b85eae3c5f4075979e290f3d22673c392e3a60 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[6] ) begin
                    I53e90d4a2bbfaffcf92f2e9fd80c491e61990aa575337df13d24211a558315a0  <=  ~I7dbeb05d89d3fea39368b48237973c682e796d24aba3438109147cc316b96ba2 + 1;
                end else begin
                    I53e90d4a2bbfaffcf92f2e9fd80c491e61990aa575337df13d24211a558315a0  <= I7dbeb05d89d3fea39368b48237973c682e796d24aba3438109147cc316b96ba2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[2] ) begin
                    I5c0776e9826af1a98810296a7cb86adde5b1b41c434e6040bc6a5a30172d1bf7  <=  ~I6e863b3eb7ba8e7ad90945ec76c695330de32ae32b69ae2a03091d1ef0142670 + 1;
                end else begin
                    I5c0776e9826af1a98810296a7cb86adde5b1b41c434e6040bc6a5a30172d1bf7  <= I6e863b3eb7ba8e7ad90945ec76c695330de32ae32b69ae2a03091d1ef0142670 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2 != Id34d005cdd89bf304f95101c6fbfdd40d6c0b1742b5f3bee3bf043bf88c3d063[0] ) begin
                    Ie55394a5e3d49de60fbc4f33b3f9813b885da2049376036c935e8cd7c85010d7  <=  ~Ib13a4de6ca8fc3856fdeaa543ff8aae727f62ebff652acce5e23c6c121ee740a + 1;
                end else begin
                    Ie55394a5e3d49de60fbc4f33b3f9813b885da2049376036c935e8cd7c85010d7  <= Ib13a4de6ca8fc3856fdeaa543ff8aae727f62ebff652acce5e23c6c121ee740a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[6] ) begin
                    I65e452247faa2c9d6b01dcbbebd5e8c31884c88e70dc8ec76d55aac7e77e2d46  <=  ~I22692863c63315b86c8a72a902c88573f4af6aa3b1691f68ed588a38ac77f7c2 + 1;
                end else begin
                    I65e452247faa2c9d6b01dcbbebd5e8c31884c88e70dc8ec76d55aac7e77e2d46  <= I22692863c63315b86c8a72a902c88573f4af6aa3b1691f68ed588a38ac77f7c2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[6] ) begin
                    I4aabce2cc01e829bb9c3d6a984cf2b5bf9230cf3913db788c47a932ddf71b869  <=  ~I2f18a4d6ae6bbfa53e26a0aa169b1cd1c40ff544f7fd42b9ac493729ffa90ce3 + 1;
                end else begin
                    I4aabce2cc01e829bb9c3d6a984cf2b5bf9230cf3913db788c47a932ddf71b869  <= I2f18a4d6ae6bbfa53e26a0aa169b1cd1c40ff544f7fd42b9ac493729ffa90ce3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[2] ) begin
                    Ib8d3655f6360b2b189b79353d38c9c9989af811109144d45af0f8b68a3276149  <=  ~I5c4daf848487e7de6d8f95704179a300218ae460e56dbe71d33805739ea61144 + 1;
                end else begin
                    Ib8d3655f6360b2b189b79353d38c9c9989af811109144d45af0f8b68a3276149  <= I5c4daf848487e7de6d8f95704179a300218ae460e56dbe71d33805739ea61144 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a != I79d61ad4114817a49b1dc8e9314d9e3be9758d861974ead362ff0ac862d1d77f[0] ) begin
                    Ia6240db37d8e82731a264e5e3eeabb88e632dc6445647a26b4abdb142ff44c03  <=  ~I94386cfbe9c6f26a678c961cdb0f15d314fc3e6bd04edc61d5596107adc68969 + 1;
                end else begin
                    Ia6240db37d8e82731a264e5e3eeabb88e632dc6445647a26b4abdb142ff44c03  <= I94386cfbe9c6f26a678c961cdb0f15d314fc3e6bd04edc61d5596107adc68969 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[6] ) begin
                    Ia4691d32d9e84827a250e0b3d6ea8142c24c9df4ade01c19583e6cfca06cd990  <=  ~Icbf8ff1f03b79fbbdd3d73ba2d399ba98a814ca4db6f6541ce67d8e5558d0eb8 + 1;
                end else begin
                    Ia4691d32d9e84827a250e0b3d6ea8142c24c9df4ade01c19583e6cfca06cd990  <= Icbf8ff1f03b79fbbdd3d73ba2d399ba98a814ca4db6f6541ce67d8e5558d0eb8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[6] ) begin
                    I52dd625c97050874c15b1980a389843c4a7a890d73f6efb003c4324c029772aa  <=  ~Ia69053f259b67f0fd728ca4fcd2bd39802adb86be01404890b17989eb74240db + 1;
                end else begin
                    I52dd625c97050874c15b1980a389843c4a7a890d73f6efb003c4324c029772aa  <= Ia69053f259b67f0fd728ca4fcd2bd39802adb86be01404890b17989eb74240db ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[2] ) begin
                    I20ddfee724da47731a2062b2732598b429c42f7d22bcfb300dc084de362a2bdb  <=  ~Id372f6f6b6b8b583699e8af0deba407a85b166caf3110f896594d222f0114cb8 + 1;
                end else begin
                    I20ddfee724da47731a2062b2732598b429c42f7d22bcfb300dc084de362a2bdb  <= Id372f6f6b6b8b583699e8af0deba407a85b166caf3110f896594d222f0114cb8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de != Icfe1fffea36cf64044389903be9550fe283d4dbb7f1b47aff2005e70765a6045[0] ) begin
                    I4dfaddc409bf6d3698f255e55590182c2c8c067e0766311322460720dbd0967d  <=  ~Id9b0a59eec0b8ceb485b7dafbff07051b5bd44c8b9ee4c3fda3773cef4450e78 + 1;
                end else begin
                    I4dfaddc409bf6d3698f255e55590182c2c8c067e0766311322460720dbd0967d  <= Id9b0a59eec0b8ceb485b7dafbff07051b5bd44c8b9ee4c3fda3773cef4450e78 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[6] ) begin
                    Iba81256fd46cc69f1367fc6ed7b712d2695e099c52b476f9b39f0a13404dceaa  <=  ~Ic0563f05659ac941778904304c02575d9c9f2125ee05515ffd05749e20880d90 + 1;
                end else begin
                    Iba81256fd46cc69f1367fc6ed7b712d2695e099c52b476f9b39f0a13404dceaa  <= Ic0563f05659ac941778904304c02575d9c9f2125ee05515ffd05749e20880d90 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[6] ) begin
                    Ie278ca9a470ffe4ac78bc335aec472b66707cf02bd91256aff2e7c73b5d2c6b6  <=  ~I81590f464fadabf1667af046de2f41172c36389854de1ad410e32cbe3b719ced + 1;
                end else begin
                    Ie278ca9a470ffe4ac78bc335aec472b66707cf02bd91256aff2e7c73b5d2c6b6  <= I81590f464fadabf1667af046de2f41172c36389854de1ad410e32cbe3b719ced ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[2] ) begin
                    Ie2c7966ff2c1e84a7ae016f31b0f8b9ca7aa42eec03467c7e3dda37dc34f070c  <=  ~Ib2f85bbcac9533694e4da81d1e86313ed14510ac8a37929a6158c888ba9cdb0c + 1;
                end else begin
                    Ie2c7966ff2c1e84a7ae016f31b0f8b9ca7aa42eec03467c7e3dda37dc34f070c  <= Ib2f85bbcac9533694e4da81d1e86313ed14510ac8a37929a6158c888ba9cdb0c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb != Ib08cf17b2065d04f587d1a8231ec1e4bbb6b2b15819de8a7efe18b477515ccf8[0] ) begin
                    I1dd3e1e1e78d9e24a54fc937e7a25fc0e2514eabd1c1cc662d81ba73aa44680b  <=  ~I6128d022628a70641f03bc8d1508dc00be5665cbb426ab6b2befa774ad124efc + 1;
                end else begin
                    I1dd3e1e1e78d9e24a54fc937e7a25fc0e2514eabd1c1cc662d81ba73aa44680b  <= I6128d022628a70641f03bc8d1508dc00be5665cbb426ab6b2befa774ad124efc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[7] ) begin
                    Ic9dc8459f6cd65f223a6386c82f754469ef74fbab59ded4fd1370fb69136c847  <=  ~I9eb8c67587f031f7dd6668286278ec62c632eebd218d4b5fca188e6447de8cff + 1;
                end else begin
                    Ic9dc8459f6cd65f223a6386c82f754469ef74fbab59ded4fd1370fb69136c847  <= I9eb8c67587f031f7dd6668286278ec62c632eebd218d4b5fca188e6447de8cff ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 != I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[3] ) begin
                    I1c886223618a03ba9e18de68462ddcc522338cd26d24b5e126da9da1df1339f4  <=  ~I930d8c08531d026f47ecb265d741cbd6a41286e3898d547ec9770fe114da36a2 + 1;
                end else begin
                    I1c886223618a03ba9e18de68462ddcc522338cd26d24b5e126da9da1df1339f4  <= I930d8c08531d026f47ecb265d741cbd6a41286e3898d547ec9770fe114da36a2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[3] ) begin
                    Ief38674752576e92e90fbe2a7abcfc952274123875a95657dd42c910133cccde  <=  ~I7401c9a97f13630805f89ca9767771302df865505689963bf68db913a151a1bd + 1;
                end else begin
                    Ief38674752576e92e90fbe2a7abcfc952274123875a95657dd42c910133cccde  <= I7401c9a97f13630805f89ca9767771302df865505689963bf68db913a151a1bd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[6] ) begin
                    Ic57569daaae5eb0e66117615c8c6043b5f76b114b5c34b0df50445f66a22849e  <=  ~I0533ded3a5c68b582fb4785c33ad5742da4947c904b1a52e05c80a3645f3fef1 + 1;
                end else begin
                    Ic57569daaae5eb0e66117615c8c6043b5f76b114b5c34b0df50445f66a22849e  <= I0533ded3a5c68b582fb4785c33ad5742da4947c904b1a52e05c80a3645f3fef1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 != I21832b7270210e1bb6a23930ad9ced36d3da201d80310263e26eb96bebd23612[0] ) begin
                    I80d4a0cc8b63f2ce0dcb344da5a47c95cc28b5f93d5bc6b77e9b875cdd58db99  <=  ~I2616f37126555e344d3b2f904a46af3f8a5fcfd59fcbf0677377f16cd59f3be5 + 1;
                end else begin
                    I80d4a0cc8b63f2ce0dcb344da5a47c95cc28b5f93d5bc6b77e9b875cdd58db99  <= I2616f37126555e344d3b2f904a46af3f8a5fcfd59fcbf0677377f16cd59f3be5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[7] ) begin
                    I11bf8ca77f64484279bd3f36febe1c6869fb79b4585a800449a0e5c683c6aa18  <=  ~Ia049b06c7b1e457c3ee5643e87fc729a409f2fa943275ce5dda083fb1253c2eb + 1;
                end else begin
                    I11bf8ca77f64484279bd3f36febe1c6869fb79b4585a800449a0e5c683c6aa18  <= Ia049b06c7b1e457c3ee5643e87fc729a409f2fa943275ce5dda083fb1253c2eb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 != I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[3] ) begin
                    I1b02edd5d00090446500b1dbf66a7e674de978c068b81ff0b0fb7abb9ffb1654  <=  ~I6d785370057273f67048d3cda9ebfb0c8bc43fc5f34af47935e45302ed66e021 + 1;
                end else begin
                    I1b02edd5d00090446500b1dbf66a7e674de978c068b81ff0b0fb7abb9ffb1654  <= I6d785370057273f67048d3cda9ebfb0c8bc43fc5f34af47935e45302ed66e021 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[3] ) begin
                    Idaf1699bc7916d99a2a5ce0174383c189dca6d7537734b19dc379bd634d0d209  <=  ~If668ac9edc8047d257ed4f162d07f8f326c0c3ffed244595bc249275f04f02b0 + 1;
                end else begin
                    Idaf1699bc7916d99a2a5ce0174383c189dca6d7537734b19dc379bd634d0d209  <= If668ac9edc8047d257ed4f162d07f8f326c0c3ffed244595bc249275f04f02b0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[6] ) begin
                    I7a7bbb1d7d9b77199c0b29fda08f8a63112052ffb0a502a05586ced336e13c62  <=  ~I8ecda1185b64bb196b1281095a7e3bf01377e6fbc7ec9cb20a3700f458944fa9 + 1;
                end else begin
                    I7a7bbb1d7d9b77199c0b29fda08f8a63112052ffb0a502a05586ced336e13c62  <= I8ecda1185b64bb196b1281095a7e3bf01377e6fbc7ec9cb20a3700f458944fa9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 != I5dcc76c47f3c9129431152fa6f7047be203fc556198b45db15a9991647bb8c85[0] ) begin
                    Iec19b0b63d20ea69dbcb23411a298bb6e833ee523fdf082f9343a695891a990f  <=  ~I4b6ef863f3c19600f1325225dfeba21b5e9333dff55ddcf9f0cd8e8ec3581a32 + 1;
                end else begin
                    Iec19b0b63d20ea69dbcb23411a298bb6e833ee523fdf082f9343a695891a990f  <= I4b6ef863f3c19600f1325225dfeba21b5e9333dff55ddcf9f0cd8e8ec3581a32 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[7] ) begin
                    I5ef535b2e573d96fd518cbd837132928a2a0c6a25d4eb3c360f1cc0aed89656c  <=  ~I2cfed4bfd244233c8d85a9ebd9edd2c03f3bbbeddb7c7a32de444794e9c44e17 + 1;
                end else begin
                    I5ef535b2e573d96fd518cbd837132928a2a0c6a25d4eb3c360f1cc0aed89656c  <= I2cfed4bfd244233c8d85a9ebd9edd2c03f3bbbeddb7c7a32de444794e9c44e17 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 != I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[3] ) begin
                    I661bc8acd80497efe43e3d6fd92bc4107b1ca63eaf162cff5695b35f8d4a7e26  <=  ~If7e91102c5105c0ecfc871fce4bfb86900fbfc837d6f06f3229d362d20e51ae0 + 1;
                end else begin
                    I661bc8acd80497efe43e3d6fd92bc4107b1ca63eaf162cff5695b35f8d4a7e26  <= If7e91102c5105c0ecfc871fce4bfb86900fbfc837d6f06f3229d362d20e51ae0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[3] ) begin
                    Id160a3b60a3c7a3ad93044461ade9ccf0b7a627efa4b1bba84a2ea0d4fbdb551  <=  ~I7643b1d4690f708c2c0d93adf0c5ac9ef99fe85eedc024e505edc74208d0f94f + 1;
                end else begin
                    Id160a3b60a3c7a3ad93044461ade9ccf0b7a627efa4b1bba84a2ea0d4fbdb551  <= I7643b1d4690f708c2c0d93adf0c5ac9ef99fe85eedc024e505edc74208d0f94f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[6] ) begin
                    I918037e81d2f9c05c6a8b94c64724b1d0ec8afafe5666df433fee3e296171f54  <=  ~I78f713264010c545a0147149b2fa2efaa92985405649e4c4313a0832e8222787 + 1;
                end else begin
                    I918037e81d2f9c05c6a8b94c64724b1d0ec8afafe5666df433fee3e296171f54  <= I78f713264010c545a0147149b2fa2efaa92985405649e4c4313a0832e8222787 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 != I450f5b0f5d2b96636ae010048040ebd744fc4ca164cd764bb33615741ecaa62f[0] ) begin
                    Ib612f39370c6527c5f6eedb0eb5e7676212642673e940402586e823ddcbfb4c6  <=  ~I6fc297df8d4527160ce05230a017f3710f7c026c6b11d64babe81959156f3462 + 1;
                end else begin
                    Ib612f39370c6527c5f6eedb0eb5e7676212642673e940402586e823ddcbfb4c6  <= I6fc297df8d4527160ce05230a017f3710f7c026c6b11d64babe81959156f3462 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[7] ) begin
                    Ie57b3acbbf1d1593e02ad38bc0e07bb84db2655f9282adb3ac5edc311e882641  <=  ~Ie3e13531d22eb604e4a351dce5ee5512894170b3dd6f87962756c534438688ea + 1;
                end else begin
                    Ie57b3acbbf1d1593e02ad38bc0e07bb84db2655f9282adb3ac5edc311e882641  <= Ie3e13531d22eb604e4a351dce5ee5512894170b3dd6f87962756c534438688ea ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 != I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[3] ) begin
                    Idb259e613b71ccde839570ff2e7f21a9cb7bf676ffd4aadfb08d6a963bea9640  <=  ~I10312c661b621655f99ef4c729f81bfd1c6aabf28b2f3372264d69d6d177d475 + 1;
                end else begin
                    Idb259e613b71ccde839570ff2e7f21a9cb7bf676ffd4aadfb08d6a963bea9640  <= I10312c661b621655f99ef4c729f81bfd1c6aabf28b2f3372264d69d6d177d475 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[3] ) begin
                    I39b8420e976cbdf011232d83446a5cb92c2ba58577792c9c61dd71358205e936  <=  ~Ic4b994b93547d46c87ce7cd1fff323144f9de0ff6e79ef0ce9ecc1db89340e6b + 1;
                end else begin
                    I39b8420e976cbdf011232d83446a5cb92c2ba58577792c9c61dd71358205e936  <= Ic4b994b93547d46c87ce7cd1fff323144f9de0ff6e79ef0ce9ecc1db89340e6b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[6] ) begin
                    I353e1673347daf260e61fbba813cd14f83c52ce3f6e5168c0fa6308d41e93590  <=  ~I38340f75bcbf775a9e070a528d926355b818091cd8e5c1792450d2713ae436bc + 1;
                end else begin
                    I353e1673347daf260e61fbba813cd14f83c52ce3f6e5168c0fa6308d41e93590  <= I38340f75bcbf775a9e070a528d926355b818091cd8e5c1792450d2713ae436bc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 != I35d64df6881fde0d4836aa408258db7cc1bfb2f066abf8c9345670b78c466b9e[0] ) begin
                    Ifa501efa24e47050960fb3c383458a20f54abcbc5ca45bbe2d15a037670cd5cd  <=  ~Iad0e03f141449cf08d3cfdfcd976e4b5a8401179533f5aa4f8216198b749a4e1 + 1;
                end else begin
                    Ifa501efa24e47050960fb3c383458a20f54abcbc5ca45bbe2d15a037670cd5cd  <= Iad0e03f141449cf08d3cfdfcd976e4b5a8401179533f5aa4f8216198b749a4e1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[7] ) begin
                    Ib0641eb8fe554f69ebb57e8e900f995c07bddadffd25c01781ba234b87af4a94  <=  ~Ibc82061cbb8fc5b88d39b5b714381ff331de2b2877376cb96a32d6742f3cac6d + 1;
                end else begin
                    Ib0641eb8fe554f69ebb57e8e900f995c07bddadffd25c01781ba234b87af4a94  <= Ibc82061cbb8fc5b88d39b5b714381ff331de2b2877376cb96a32d6742f3cac6d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[8] ) begin
                    Ic486b9953b158eae95a2d8914f8144e669e056675946d245c8239bfc249a16ac  <=  ~I49af7bf73e330c26c437d8f0447a930c63d4677498d07a28ff9b2b25860258d0 + 1;
                end else begin
                    Ic486b9953b158eae95a2d8914f8144e669e056675946d245c8239bfc249a16ac  <= I49af7bf73e330c26c437d8f0447a930c63d4677498d07a28ff9b2b25860258d0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[3] ) begin
                    If270910122bcee1c18cc592dba9b38c026f792d8d1472400a09edee9d7633e22  <=  ~I5e977efb6007fb448a0cd05362289e5bbace24ff868e4fb623ba54135e53fc82 + 1;
                end else begin
                    If270910122bcee1c18cc592dba9b38c026f792d8d1472400a09edee9d7633e22  <= I5e977efb6007fb448a0cd05362289e5bbace24ff868e4fb623ba54135e53fc82 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[5] ) begin
                    Ia79355adc994f77e150b93a3e38c8bd6f0a5848a212ac64559cf1210ee0d11d7  <=  ~I98233f63b47681b1d8b5e3decd1ab8ad783734a17e2b27c88234f00b23fa30cb + 1;
                end else begin
                    Ia79355adc994f77e150b93a3e38c8bd6f0a5848a212ac64559cf1210ee0d11d7  <= I98233f63b47681b1d8b5e3decd1ab8ad783734a17e2b27c88234f00b23fa30cb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 != I11944fb91fa1b1d5f076cc36db77f0f8434f0edbb1236c7a9bcb45f79432ea9f[0] ) begin
                    I8f088dd043a22011add21694f90df62fe1d2f6670cc72cfee805c9fb49756c77  <=  ~I58660674a5ad4c7022a05e5cfcd03fdc7161e65e8050cc59ae6fefc404b6b310 + 1;
                end else begin
                    I8f088dd043a22011add21694f90df62fe1d2f6670cc72cfee805c9fb49756c77  <= I58660674a5ad4c7022a05e5cfcd03fdc7161e65e8050cc59ae6fefc404b6b310 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[7] ) begin
                    I3a1380b85cc7f797ff92d02b7081d1ec3ba069aac74162ca059c399daa10690d  <=  ~I9612c348b28222bc7559977c8bd902d73267c977bfbe179506c88be746830331 + 1;
                end else begin
                    I3a1380b85cc7f797ff92d02b7081d1ec3ba069aac74162ca059c399daa10690d  <= I9612c348b28222bc7559977c8bd902d73267c977bfbe179506c88be746830331 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[8] ) begin
                    I632095e999af63661b01bfe8bad0078cfc2e74217253d3971230968c235bc526  <=  ~Ifea5f415406637bbe581d11e57aaab23cecc2dc1957f45152f03d3006334d24c + 1;
                end else begin
                    I632095e999af63661b01bfe8bad0078cfc2e74217253d3971230968c235bc526  <= Ifea5f415406637bbe581d11e57aaab23cecc2dc1957f45152f03d3006334d24c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[3] ) begin
                    Idc29625b375c44e890e371217aaa25d5fda337ba8177fcceca881adc72292a3b  <=  ~Ie56c2e96de8be01add59d3005f52661524c2193f6bd0fae2a759d4afe9607388 + 1;
                end else begin
                    Idc29625b375c44e890e371217aaa25d5fda337ba8177fcceca881adc72292a3b  <= Ie56c2e96de8be01add59d3005f52661524c2193f6bd0fae2a759d4afe9607388 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[5] ) begin
                    I7cd9dadb64725f4217f1330c893724a7537a616ef41d9dc49fd2794125e0dc3d  <=  ~I1744ca88c13acb5d2afa42ffe0ee5823eab5e32cbcf3248db4faffd6fe9e2537 + 1;
                end else begin
                    I7cd9dadb64725f4217f1330c893724a7537a616ef41d9dc49fd2794125e0dc3d  <= I1744ca88c13acb5d2afa42ffe0ee5823eab5e32cbcf3248db4faffd6fe9e2537 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 != I49642204473312df5a3bcab2692aa7558f44f21416226675a4ec10b0543cc5e9[0] ) begin
                    Id86d515c6d081de87b9ed3c3521ab079e93ee082d8a0b396d44b3b70cac06b9b  <=  ~I2646e32dd3a69da746d970611fa0a89f96286df22ebdcef1ab746d70c4db4331 + 1;
                end else begin
                    Id86d515c6d081de87b9ed3c3521ab079e93ee082d8a0b396d44b3b70cac06b9b  <= I2646e32dd3a69da746d970611fa0a89f96286df22ebdcef1ab746d70c4db4331 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[7] ) begin
                    I608b794037b45c46a29ea01e378b63a1f267c4b489b0866fe2f6090936fa9d44  <=  ~I4c7da80c76f8d8ad9ed1199810aaa919460f955b2745ae54cdea9276ad5e2491 + 1;
                end else begin
                    I608b794037b45c46a29ea01e378b63a1f267c4b489b0866fe2f6090936fa9d44  <= I4c7da80c76f8d8ad9ed1199810aaa919460f955b2745ae54cdea9276ad5e2491 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[8] ) begin
                    Ib22de4dadb6e63ea49c52cd8bc86dadfd7b73a002dd8e726a9cf1b7b299a8c46  <=  ~I1e411a908fa94c50629647023bf56aaf275299c8c49933fe67ccf00d3ed68d7b + 1;
                end else begin
                    Ib22de4dadb6e63ea49c52cd8bc86dadfd7b73a002dd8e726a9cf1b7b299a8c46  <= I1e411a908fa94c50629647023bf56aaf275299c8c49933fe67ccf00d3ed68d7b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[3] ) begin
                    I76599c709cdbb3f3cfe4071b96fb7dcdf8e072fe85ad5c8e7bbabd4f6182303a  <=  ~Ia06978f4049096a298ffcdf526e89060e8f27418076fa351962ec6f407576753 + 1;
                end else begin
                    I76599c709cdbb3f3cfe4071b96fb7dcdf8e072fe85ad5c8e7bbabd4f6182303a  <= Ia06978f4049096a298ffcdf526e89060e8f27418076fa351962ec6f407576753 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[5] ) begin
                    If0d62663c8a08719b83a27c76fa62525eb14d452d4ff0f33e94c67f58d7c86f9  <=  ~I93695abbc93c5e195bbc5a1fee05aa7ceb4c58b273ed67ec6f28538aef0843e4 + 1;
                end else begin
                    If0d62663c8a08719b83a27c76fa62525eb14d452d4ff0f33e94c67f58d7c86f9  <= I93695abbc93c5e195bbc5a1fee05aa7ceb4c58b273ed67ec6f28538aef0843e4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a != I24e0d361a2679430549932a968d7cc25f980275fea5554e3453ed0a652d31caa[0] ) begin
                    I4f94812066080b656de1a2807f5f669b2a81085bfc0470f9868bf5945856b451  <=  ~I81b17367c5766001911129ae2370c1dc7b3509565fe78fa6e552b7ef936da360 + 1;
                end else begin
                    I4f94812066080b656de1a2807f5f669b2a81085bfc0470f9868bf5945856b451  <= I81b17367c5766001911129ae2370c1dc7b3509565fe78fa6e552b7ef936da360 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[7] ) begin
                    I31ca3705bdc7e063c61023d93193b3ced40cf440afd817d0d730f6c8d37f8b92  <=  ~I189d5a40f26a8b2893b53242a4ec7613797831a4a2192289df09283c7da753d8 + 1;
                end else begin
                    I31ca3705bdc7e063c61023d93193b3ced40cf440afd817d0d730f6c8d37f8b92  <= I189d5a40f26a8b2893b53242a4ec7613797831a4a2192289df09283c7da753d8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[8] ) begin
                    I255a6c7b69c31d60711a86b1f0da51040ab60c48952002406e028a200a835049  <=  ~I15429bf02bcaf6ac17ed02efb1e65c5c37254aedb9ef6181c2731c3f7e2a829d + 1;
                end else begin
                    I255a6c7b69c31d60711a86b1f0da51040ab60c48952002406e028a200a835049  <= I15429bf02bcaf6ac17ed02efb1e65c5c37254aedb9ef6181c2731c3f7e2a829d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[3] ) begin
                    I58c6fbcd5f77398c3514e6a850bb69d9f57880a387f10132aa63079c0a1f4857  <=  ~I1807ee521c06cb799faa136864a31c00869398289b0e3b185e702f42cb0e7412 + 1;
                end else begin
                    I58c6fbcd5f77398c3514e6a850bb69d9f57880a387f10132aa63079c0a1f4857  <= I1807ee521c06cb799faa136864a31c00869398289b0e3b185e702f42cb0e7412 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[5] ) begin
                    I9331a9d6610ae5cb77aa3d477fce0c0ad7378a884c86c4872a1573f2d8a90d8c  <=  ~Id4ff3dcea8b6c38c5288cac263296941b841255967f2f58fa97a49fadb2fd2c8 + 1;
                end else begin
                    I9331a9d6610ae5cb77aa3d477fce0c0ad7378a884c86c4872a1573f2d8a90d8c  <= Id4ff3dcea8b6c38c5288cac263296941b841255967f2f58fa97a49fadb2fd2c8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 != I386015f8daacd2ac9cfed376d3418b56ac13f075a43dde939e4056c29565a926[0] ) begin
                    Ia92baf4463c96e210b460ea02d7775353edc6d475d7a315b594b9798cfd17900  <=  ~I3856054a7ed02c524f8816bd8ba22a48935b393ced40e98c693416364ff512b3 + 1;
                end else begin
                    Ia92baf4463c96e210b460ea02d7775353edc6d475d7a315b594b9798cfd17900  <= I3856054a7ed02c524f8816bd8ba22a48935b393ced40e98c693416364ff512b3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[8] ) begin
                    Iee9c2c6a9b8e84402eb1e0de611c1cb8ae1e802226f2c07833bafaba74f1ac15  <=  ~I358ca9d90eebc0e19c434a7d1070a69b3c20b4f8152adcc45c0b73e8cf2c9902 + 1;
                end else begin
                    Iee9c2c6a9b8e84402eb1e0de611c1cb8ae1e802226f2c07833bafaba74f1ac15  <= I358ca9d90eebc0e19c434a7d1070a69b3c20b4f8152adcc45c0b73e8cf2c9902 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[6] ) begin
                    I48d9ec419ebe83e2a5a8281e7beac36acc9e554b86b154736dc51ff940f5348d  <=  ~I1e60aaae452f97c016f3f3929c33637509d02988bea72048f7901a440232a85a + 1;
                end else begin
                    I48d9ec419ebe83e2a5a8281e7beac36acc9e554b86b154736dc51ff940f5348d  <= I1e60aaae452f97c016f3f3929c33637509d02988bea72048f7901a440232a85a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[4] ) begin
                    If145a331c8a8abde8c26d2571cc8b38e1eaf2768a4658d350cb602bf8614a521  <=  ~I312753748b2d173f2dde21bfad8dcf880f5fae94cd73fea4dbedb01c43c99b43 + 1;
                end else begin
                    If145a331c8a8abde8c26d2571cc8b38e1eaf2768a4658d350cb602bf8614a521  <= I312753748b2d173f2dde21bfad8dcf880f5fae94cd73fea4dbedb01c43c99b43 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[3] ) begin
                    Ibae8222f76059e8f61dff938a64e23080eb668880ac50ecbb50de852472a22ad  <=  ~I6f210ff43165afc5b4c3a9a22dab74940c409a5fbdf9c47b9eaa68fa08918f23 + 1;
                end else begin
                    Ibae8222f76059e8f61dff938a64e23080eb668880ac50ecbb50de852472a22ad  <= I6f210ff43165afc5b4c3a9a22dab74940c409a5fbdf9c47b9eaa68fa08918f23 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 != I32832b039ae7e6f4b1e38cfdf680e5044e383b921a76189054511ebe5b8c0d7c[0] ) begin
                    I9d4c230c86454c5c5f9ec98917ffc8d23fd19105ef93ba860ac2650bcf43ba4d  <=  ~I3422d7c29697052f1d70152dce7d92858081099a7bd19bcb2a48add3d660ef12 + 1;
                end else begin
                    I9d4c230c86454c5c5f9ec98917ffc8d23fd19105ef93ba860ac2650bcf43ba4d  <= I3422d7c29697052f1d70152dce7d92858081099a7bd19bcb2a48add3d660ef12 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[8] ) begin
                    I14919dedf2b4d4caae8efa1726435d1946f48e1e9b1052133bebe8affeb3556d  <=  ~I90ed9972249e176fb13ac19818b591acc7f7048588409d394fbbb79ac26b3519 + 1;
                end else begin
                    I14919dedf2b4d4caae8efa1726435d1946f48e1e9b1052133bebe8affeb3556d  <= I90ed9972249e176fb13ac19818b591acc7f7048588409d394fbbb79ac26b3519 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[6] ) begin
                    I1b68e82cfc8606d3a9325ff2da047f345e2f34b44eb428bf2a3bdcf42a6e869e  <=  ~Iee565a93d37ce096492969d59077dd347ffeabe00c447298bd22adb6f66926dc + 1;
                end else begin
                    I1b68e82cfc8606d3a9325ff2da047f345e2f34b44eb428bf2a3bdcf42a6e869e  <= Iee565a93d37ce096492969d59077dd347ffeabe00c447298bd22adb6f66926dc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[4] ) begin
                    I9cd4ac82c1e6f2dab27efa85314df34a40d8747959eba18330bd424a38debece  <=  ~I8ef1e4ffe1fdc795a0b74f93f87b834e26e14a3a6cf78496df39c9cbdc70a819 + 1;
                end else begin
                    I9cd4ac82c1e6f2dab27efa85314df34a40d8747959eba18330bd424a38debece  <= I8ef1e4ffe1fdc795a0b74f93f87b834e26e14a3a6cf78496df39c9cbdc70a819 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[3] ) begin
                    Iadfdcb3c0764107a2b0deaaf039babe6a08f1018f3718f5539718ed6a5aa962d  <=  ~I7bcdd7375cc16a2a91d81c5608f9953d21293d5121600dc475a15b190967b143 + 1;
                end else begin
                    Iadfdcb3c0764107a2b0deaaf039babe6a08f1018f3718f5539718ed6a5aa962d  <= I7bcdd7375cc16a2a91d81c5608f9953d21293d5121600dc475a15b190967b143 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 != I09fff9b84a38f3d19685f9627d01a7183cf65d72110802f11e8da0e01194bf88[0] ) begin
                    Ia4a28d520896fadbeabee4130dcf862a9542852d87be480b1df2b67817f0ce65  <=  ~I75bab5d1e71ba5ad182fb01cfa39d37572ab33f5f848dd0775e3358154e4644f + 1;
                end else begin
                    Ia4a28d520896fadbeabee4130dcf862a9542852d87be480b1df2b67817f0ce65  <= I75bab5d1e71ba5ad182fb01cfa39d37572ab33f5f848dd0775e3358154e4644f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[8] ) begin
                    Ic48347f5264e8e479996a8dba0171a108b602be1e1d24b2fcb43cd2bdb82f61d  <=  ~I7f17ac4c0a37a850db6a1d3c1a5b2483c0f3afd684853df30d66933c8c593d03 + 1;
                end else begin
                    Ic48347f5264e8e479996a8dba0171a108b602be1e1d24b2fcb43cd2bdb82f61d  <= I7f17ac4c0a37a850db6a1d3c1a5b2483c0f3afd684853df30d66933c8c593d03 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[6] ) begin
                    Ibdd77bf8b31352e365f7e6440a57247a8ba62e667b000c1347165bb39f3c7c2b  <=  ~I6f8e6ce3128ce55b822fddcc664d0340c940bc85adbb5c93acff37548e3018fe + 1;
                end else begin
                    Ibdd77bf8b31352e365f7e6440a57247a8ba62e667b000c1347165bb39f3c7c2b  <= I6f8e6ce3128ce55b822fddcc664d0340c940bc85adbb5c93acff37548e3018fe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[4] ) begin
                    Iad8ee4f6cd13a9f415cd3519de0179a66cfc993a840b3101cee554b55c0e7e7a  <=  ~I3234faedbd9c50f29c09060c3f7ad76e44648841500b09c499875ea77aad9537 + 1;
                end else begin
                    Iad8ee4f6cd13a9f415cd3519de0179a66cfc993a840b3101cee554b55c0e7e7a  <= I3234faedbd9c50f29c09060c3f7ad76e44648841500b09c499875ea77aad9537 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[3] ) begin
                    I00e5abb30adb527f6b32257212dc21f9797e9793ebbcc10feae9e524188539d2  <=  ~I74189716f0b6628c0d75d54cd0815cd8fa65b9047c3f51c5218fa0ba7b7fc47f + 1;
                end else begin
                    I00e5abb30adb527f6b32257212dc21f9797e9793ebbcc10feae9e524188539d2  <= I74189716f0b6628c0d75d54cd0815cd8fa65b9047c3f51c5218fa0ba7b7fc47f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 != Ib82c65f09934744abbba984b6e375bd69ce7231a5085bb00ba4e673cfd3aba38[0] ) begin
                    Ide9498000905141bb106efc7e2184bd460d0e59a2270b10d42f981cf3bd514cb  <=  ~Icaffca7436caceaf13fa42e9e496c7b149d5931e08057ec92a73fbeb9e610648 + 1;
                end else begin
                    Ide9498000905141bb106efc7e2184bd460d0e59a2270b10d42f981cf3bd514cb  <= Icaffca7436caceaf13fa42e9e496c7b149d5931e08057ec92a73fbeb9e610648 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[8] ) begin
                    I789461a909fa4abaf3840dfca4f63bfa63fdab389e149fddb7d8ae2b876dc912  <=  ~I13009f7de199aa969d82e233d26476e44aa1bfbb7d8a4fbfa0fe4f1f1e7579ff + 1;
                end else begin
                    I789461a909fa4abaf3840dfca4f63bfa63fdab389e149fddb7d8ae2b876dc912  <= I13009f7de199aa969d82e233d26476e44aa1bfbb7d8a4fbfa0fe4f1f1e7579ff ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[6] ) begin
                    Ifedfb1db4b16b86149f5eb8b0adf06499331d423c368c0077c738a190a1814f0  <=  ~I8c7ca4914849b513537d3688dc1b76461348ca06e80e489afb60a2a082e905bd + 1;
                end else begin
                    Ifedfb1db4b16b86149f5eb8b0adf06499331d423c368c0077c738a190a1814f0  <= I8c7ca4914849b513537d3688dc1b76461348ca06e80e489afb60a2a082e905bd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[4] ) begin
                    Ib63856036797d30e60f13453da509ace15e3324c25bdfdea5aa495d592e2006a  <=  ~I9117209a7cbd232356943389578d67bb7d6c217e7e40bdbb904fb46fb00e9385 + 1;
                end else begin
                    Ib63856036797d30e60f13453da509ace15e3324c25bdfdea5aa495d592e2006a  <= I9117209a7cbd232356943389578d67bb7d6c217e7e40bdbb904fb46fb00e9385 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[3] ) begin
                    Ibb57ab5a5468d08c8b299ee67b535b83995e94d6223d0c6d93dba8580906e319  <=  ~I0f16d6ab2d87cb715b071b05ad14fc6be271b1d7966b71c80795894643e6fc91 + 1;
                end else begin
                    Ibb57ab5a5468d08c8b299ee67b535b83995e94d6223d0c6d93dba8580906e319  <= I0f16d6ab2d87cb715b071b05ad14fc6be271b1d7966b71c80795894643e6fc91 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa != I8ec5727130bf67c04580aa1b5b46cdf964db65750f2fc9ce55025b1c117b2bef[0] ) begin
                    Ie9a6b0e499ede3f80403e8f9c795ef4e93108ee8db755e12fb931259f1699712  <=  ~I9fe8ab2f590451df0986a4f7a74194c27699bdfae0f182440f4c1875633cfcf3 + 1;
                end else begin
                    Ie9a6b0e499ede3f80403e8f9c795ef4e93108ee8db755e12fb931259f1699712  <= I9fe8ab2f590451df0986a4f7a74194c27699bdfae0f182440f4c1875633cfcf3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[9] ) begin
                    Id6c8c2ebab66fb903f108466c8d15060ed1328fe9a979858569c39069bf050c7  <=  ~I57876d51522e735eff337a69dc597cdcbb100bb3d3e0e541aad4428637f34e26 + 1;
                end else begin
                    Id6c8c2ebab66fb903f108466c8d15060ed1328fe9a979858569c39069bf050c7  <= I57876d51522e735eff337a69dc597cdcbb100bb3d3e0e541aad4428637f34e26 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec != I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[3] ) begin
                    I6687de5f8cb258492154a67fd3a3d5ee88d97a4db1c6c273ad158d5205ae3b48  <=  ~I9fc6ec0055cf4788a1f382e41d1bd50b2ee07f2cdacf368e2075fdeef55f53b5 + 1;
                end else begin
                    I6687de5f8cb258492154a67fd3a3d5ee88d97a4db1c6c273ad158d5205ae3b48  <= I9fc6ec0055cf4788a1f382e41d1bd50b2ee07f2cdacf368e2075fdeef55f53b5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[7] ) begin
                    Idf77a6217d51b2439f71afbf5956a52a241f2bf8722f54cb166d83c3b45f6721  <=  ~Ib2ce92509ff0447a434264639ad96df47b161136cea1535b3e802c0c4ebc32e8 + 1;
                end else begin
                    Idf77a6217d51b2439f71afbf5956a52a241f2bf8722f54cb166d83c3b45f6721  <= Ib2ce92509ff0447a434264639ad96df47b161136cea1535b3e802c0c4ebc32e8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec != I862dddc300df692e8bbf4ca45a24d840e51ac1e975631cf4ebb8337ceefc2eb1[0] ) begin
                    I362132341c8e8a464a2bc93e7cc5b1d9d7804dd93965614dc340b48fad5c92da  <=  ~I20b66d31e195a0db14cc87da1f6d8810b5f1056c2250bd5cfcb02fb4edc9dd0e + 1;
                end else begin
                    I362132341c8e8a464a2bc93e7cc5b1d9d7804dd93965614dc340b48fad5c92da  <= I20b66d31e195a0db14cc87da1f6d8810b5f1056c2250bd5cfcb02fb4edc9dd0e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[9] ) begin
                    I24bc395a7644f2a2d7702656737c32662f8c2e8a7e2b2d4c1bca200dcdf49219  <=  ~Ie7595f637907686de85c9038415609949a80fee8bbb0c4e9f3873225ae6c56bc + 1;
                end else begin
                    I24bc395a7644f2a2d7702656737c32662f8c2e8a7e2b2d4c1bca200dcdf49219  <= Ie7595f637907686de85c9038415609949a80fee8bbb0c4e9f3873225ae6c56bc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef != I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[3] ) begin
                    I67183da8c2763243a285b7cd41d838337f98eb6e59feaaa0a9150bcd6c29877b  <=  ~I6d41031fb10896690dda6067df08ad914896baaa5f83c46b4051cd5a02f3baef + 1;
                end else begin
                    I67183da8c2763243a285b7cd41d838337f98eb6e59feaaa0a9150bcd6c29877b  <= I6d41031fb10896690dda6067df08ad914896baaa5f83c46b4051cd5a02f3baef ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[7] ) begin
                    I5cbbcfd1cfc35b3e78d01b29831195106ebd9ba5907f44dee6761c2b047c4a60  <=  ~Idc6c8bd2a37e01dec18007c8fa763941f7016bf299e3cebbbbee3066d4bf8c7b + 1;
                end else begin
                    I5cbbcfd1cfc35b3e78d01b29831195106ebd9ba5907f44dee6761c2b047c4a60  <= Idc6c8bd2a37e01dec18007c8fa763941f7016bf299e3cebbbbee3066d4bf8c7b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef != Id08a37df0c5095196e2d760938c4d0b7e8716c25b55d9a9656d86c2c473f9c2f[0] ) begin
                    I4b3c222863418745872c878545e419ee8f9c531f2cba89d28f0787992b0be8ed  <=  ~Iac1565ee006c23dca041f0aaff4dd7023b8a22cb72c9f206170be661a66d4732 + 1;
                end else begin
                    I4b3c222863418745872c878545e419ee8f9c531f2cba89d28f0787992b0be8ed  <= Iac1565ee006c23dca041f0aaff4dd7023b8a22cb72c9f206170be661a66d4732 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[9] ) begin
                    Id89c8a47964d1e4aa4bb9e96a79092cf7fb55eee5808d6323ecbdecf8926adcd  <=  ~I7318d295676d4cc0682f246020963a6411be5cfc2fa525dd7af0f2e651b4f9f8 + 1;
                end else begin
                    Id89c8a47964d1e4aa4bb9e96a79092cf7fb55eee5808d6323ecbdecf8926adcd  <= I7318d295676d4cc0682f246020963a6411be5cfc2fa525dd7af0f2e651b4f9f8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d != Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[3] ) begin
                    I1e8142c7ece070c02ed90211fbeb423bc2a4ab19fae011793be99c68ff103705  <=  ~I596ee6206f54965079551ffb23aa3c1948f6fbcd48659c4e30b205dd06de79f6 + 1;
                end else begin
                    I1e8142c7ece070c02ed90211fbeb423bc2a4ab19fae011793be99c68ff103705  <= I596ee6206f54965079551ffb23aa3c1948f6fbcd48659c4e30b205dd06de79f6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[7] ) begin
                    Ie1657c5216d7c6e743a23819c08b7c7f2fc8a56793e1bc67fa5c5f3b37976641  <=  ~I7c8c24bd3806dbea5552d386a7363828eb5a822bb292fa0c14ba407a1937d11d + 1;
                end else begin
                    Ie1657c5216d7c6e743a23819c08b7c7f2fc8a56793e1bc67fa5c5f3b37976641  <= I7c8c24bd3806dbea5552d386a7363828eb5a822bb292fa0c14ba407a1937d11d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d != I40204cd18eb803f82fc3ef933553c6ec41331f6d4a15538c287b8f57adebb89e[0] ) begin
                    Ie39e570f1b5dd9f1ae893af78d81e458d077fcde2aeaba432209269b79785582  <=  ~Ib7690a963a38d899184e89d3e51ac5cd99cc0ea9b2fca1c2e36e51ea65b893ac + 1;
                end else begin
                    Ie39e570f1b5dd9f1ae893af78d81e458d077fcde2aeaba432209269b79785582  <= Ib7690a963a38d899184e89d3e51ac5cd99cc0ea9b2fca1c2e36e51ea65b893ac ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[9] ) begin
                    I6a66a98136fb7fe52fd830d869dc53a3855a545aedc1d16927f76bc12e319060  <=  ~Ie55d9e9e5c4a66363393994597d9138fccd6c11a2a6c939768b63d9cf933ae1a + 1;
                end else begin
                    I6a66a98136fb7fe52fd830d869dc53a3855a545aedc1d16927f76bc12e319060  <= Ie55d9e9e5c4a66363393994597d9138fccd6c11a2a6c939768b63d9cf933ae1a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00 != Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[3] ) begin
                    Ie130bec82505842b184f5dd86865ab095110bc65e59662767e152f427dd7462c  <=  ~Id2a5a1513f2b8c1f000f58640c3650ae03d4d56205a8cbd04742be5b91c8c594 + 1;
                end else begin
                    Ie130bec82505842b184f5dd86865ab095110bc65e59662767e152f427dd7462c  <= Id2a5a1513f2b8c1f000f58640c3650ae03d4d56205a8cbd04742be5b91c8c594 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[7] ) begin
                    I136f70cfdde5473f8944efa2b1093ed76f82dd06a341413ee2a56054ebef5fd2  <=  ~I9a2e9ef69e2c24fdb342d3334d2b71a1bebf10ffe1518dc5f3ebd5ff34dc719a + 1;
                end else begin
                    I136f70cfdde5473f8944efa2b1093ed76f82dd06a341413ee2a56054ebef5fd2  <= I9a2e9ef69e2c24fdb342d3334d2b71a1bebf10ffe1518dc5f3ebd5ff34dc719a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00 != I677f733f4e801d99dc2fd1987683a7ac6c8609d84da6c95b8a7056ce07845665[0] ) begin
                    I50ebc7f8f7cf324814b5885b2b18c90bf5007d8030744263d6e66880d836eea0  <=  ~I8052be48c5148738c00fa7e5be66ac6898d51e7fca2e5905ef028d897d47b236 + 1;
                end else begin
                    I50ebc7f8f7cf324814b5885b2b18c90bf5007d8030744263d6e66880d836eea0  <= I8052be48c5148738c00fa7e5be66ac6898d51e7fca2e5905ef028d897d47b236 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[9] ) begin
                    I443435c78145236b927711299e8bedd0d29a743e3784ac22f70b2284b6be11c1  <=  ~Ifc4766e0c1913ae910a794a3de1155638a9352251d646b270e3aba4eac09aa31 + 1;
                end else begin
                    I443435c78145236b927711299e8bedd0d29a743e3784ac22f70b2284b6be11c1  <= Ifc4766e0c1913ae910a794a3de1155638a9352251d646b270e3aba4eac09aa31 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[10] ) begin
                    Ifea15bb5031583fe42f92f554866179105e46b1eac3c6b691958a998c26ac2da  <=  ~I2322db4da4e5112d362e202ee964c08830d852a01c92f802c1c8bc2978ba25e6 + 1;
                end else begin
                    Ifea15bb5031583fe42f92f554866179105e46b1eac3c6b691958a998c26ac2da  <= I2322db4da4e5112d362e202ee964c08830d852a01c92f802c1c8bc2978ba25e6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b != I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[4] ) begin
                    I2c865426b0f044469b391bbc13f977fdd19dc89c908574ba289388e382d55cbc  <=  ~If29e3e5b3c3425bf0fd40a98d32046f215032a8ae181688dff1c4a253b0460ef + 1;
                end else begin
                    I2c865426b0f044469b391bbc13f977fdd19dc89c908574ba289388e382d55cbc  <= If29e3e5b3c3425bf0fd40a98d32046f215032a8ae181688dff1c4a253b0460ef ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[4] ) begin
                    I9349cba960e03e6068aa27e997993b0c466e040a1ee9e6053536d3346c84214f  <=  ~I51e9d69995015664cbb95900d25d26d386de1f49fa7b7d612964802060fd7a8b + 1;
                end else begin
                    I9349cba960e03e6068aa27e997993b0c466e040a1ee9e6053536d3346c84214f  <= I51e9d69995015664cbb95900d25d26d386de1f49fa7b7d612964802060fd7a8b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b != Ifeb10787a88bae5943b616e3bf751faff5e7eea80e45e24d60a760f4d6b0154c[0] ) begin
                    I326b57b49d3fcfe654c4cb9ebcd6edc0ad7969e3b531f498e3c31270a5c4aa70  <=  ~I2af69278f44ee2d81c64b9447b85bd09d2ce2a8dc86bacb9a175b33f72d4f851 + 1;
                end else begin
                    I326b57b49d3fcfe654c4cb9ebcd6edc0ad7969e3b531f498e3c31270a5c4aa70  <= I2af69278f44ee2d81c64b9447b85bd09d2ce2a8dc86bacb9a175b33f72d4f851 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[9] ) begin
                    I852a201bdaecd968b6f9c9b6bd64dc8035a17fb92ffc806a690781666354b069  <=  ~Ib82fbfc182e6598a7a8dbae45ea083d2922e3f10e781ac40e1c89f79097f1f23 + 1;
                end else begin
                    I852a201bdaecd968b6f9c9b6bd64dc8035a17fb92ffc806a690781666354b069  <= Ib82fbfc182e6598a7a8dbae45ea083d2922e3f10e781ac40e1c89f79097f1f23 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[10] ) begin
                    I385f4177f3a22b6fa4a6352d164c7d54c94b980806080c51d00a65f030966110  <=  ~Ie3180a2d7f37d66f9895c1de89329e69ef7e88d0808fce147b25636e639efdd5 + 1;
                end else begin
                    I385f4177f3a22b6fa4a6352d164c7d54c94b980806080c51d00a65f030966110  <= Ie3180a2d7f37d66f9895c1de89329e69ef7e88d0808fce147b25636e639efdd5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 != I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[4] ) begin
                    Ic72f2f8a61b8ecf8960d476bcf8fbbfd4389e932377679286e7182cc12c418c8  <=  ~Ifb545544cfc26097f08bb8236d489536608fd3ef900015de2da0a8a5dfcd44ef + 1;
                end else begin
                    Ic72f2f8a61b8ecf8960d476bcf8fbbfd4389e932377679286e7182cc12c418c8  <= Ifb545544cfc26097f08bb8236d489536608fd3ef900015de2da0a8a5dfcd44ef ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[4] ) begin
                    I6fdc128e94d85f0f7f884ee1ff44fdb6de2ad5b93d83c3e36ae235afcd3d23c0  <=  ~I90ba4bf676fa4d1eb6132a37c0b4a580ef39ac1cc44d6111b84d6c7b907922b2 + 1;
                end else begin
                    I6fdc128e94d85f0f7f884ee1ff44fdb6de2ad5b93d83c3e36ae235afcd3d23c0  <= I90ba4bf676fa4d1eb6132a37c0b4a580ef39ac1cc44d6111b84d6c7b907922b2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 != Iecc97eedc286cd1c3d301e35036e81a10d164d59da9252a92ca5f355a828367b[0] ) begin
                    Id3898be2185f86831f58bd16651edee3d1bb21fa07b33a1928740ab496404178  <=  ~Ie66d53b4bed43cf8037cd1937f7562e7bdd6cac54cfc8313572b853088528a0f + 1;
                end else begin
                    Id3898be2185f86831f58bd16651edee3d1bb21fa07b33a1928740ab496404178  <= Ie66d53b4bed43cf8037cd1937f7562e7bdd6cac54cfc8313572b853088528a0f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[9] ) begin
                    Ib62b5b3c80d193b97bd6b5c0d5678e424026381949c3f24546d367df930cbcae  <=  ~Id812808edf2372138b1569ea1a2ae0583ef70eaad98a941b8394d5d9efeb44c5 + 1;
                end else begin
                    Ib62b5b3c80d193b97bd6b5c0d5678e424026381949c3f24546d367df930cbcae  <= Id812808edf2372138b1569ea1a2ae0583ef70eaad98a941b8394d5d9efeb44c5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[10] ) begin
                    Ia84166c5479fb08b9d5bafbf3446230d231e77cb1a3034b53477e2f0632ca74a  <=  ~I6b9daca681053a70322aec979459e65099a78668854de86dd3f51ad58c5dced5 + 1;
                end else begin
                    Ia84166c5479fb08b9d5bafbf3446230d231e77cb1a3034b53477e2f0632ca74a  <= I6b9daca681053a70322aec979459e65099a78668854de86dd3f51ad58c5dced5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 != I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[4] ) begin
                    Ie9b1b4412060f1e9acccc1f3ff897bce33f24fea3bfc91266f9e42c1f38aaaad  <=  ~Ieafce3772abd32b8004981fe3f3d102d629075a15b6dfff65169984219911dd9 + 1;
                end else begin
                    Ie9b1b4412060f1e9acccc1f3ff897bce33f24fea3bfc91266f9e42c1f38aaaad  <= Ieafce3772abd32b8004981fe3f3d102d629075a15b6dfff65169984219911dd9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[4] ) begin
                    I09673e64aaf6f35dbf4aae16ffba969d08a800d32ab25413bfcdbd540d7b01f3  <=  ~I279bb276ee61f29e0c143251191c161862c9d95cf0bf3a3fdcb6b3d6acaee983 + 1;
                end else begin
                    I09673e64aaf6f35dbf4aae16ffba969d08a800d32ab25413bfcdbd540d7b01f3  <= I279bb276ee61f29e0c143251191c161862c9d95cf0bf3a3fdcb6b3d6acaee983 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 != Ia9a21e6f22a6cc828e041980ab142b418938a92bf8e868216402a46b8c614a19[0] ) begin
                    I2aa77512781cba636ab96a5d09527e1ac34623ea2bb6c6a8d742bbcf6eff499a  <=  ~Ife98dd3babdd2b2db4edbc673874d3f8f184f531c9d96b1a89b68ba60a9a57d1 + 1;
                end else begin
                    I2aa77512781cba636ab96a5d09527e1ac34623ea2bb6c6a8d742bbcf6eff499a  <= Ife98dd3babdd2b2db4edbc673874d3f8f184f531c9d96b1a89b68ba60a9a57d1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[9] ) begin
                    I6ff3298d93471156b56cfbbea17c8dc0405bfe8654e9f830bb33bc6c9a649b3e  <=  ~I038f11e434287c1e184cece6178f4ce26889bc2ea583aba8889b8953306e2e60 + 1;
                end else begin
                    I6ff3298d93471156b56cfbbea17c8dc0405bfe8654e9f830bb33bc6c9a649b3e  <= I038f11e434287c1e184cece6178f4ce26889bc2ea583aba8889b8953306e2e60 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[10] ) begin
                    Id1e80f29821e7ae727d759f44b21e84843025c938468caf7c8adfba52f1cae43  <=  ~I25c61073e64c8149ae96f3157045d317349321841e21a3d69b3baf3bd70bbd03 + 1;
                end else begin
                    Id1e80f29821e7ae727d759f44b21e84843025c938468caf7c8adfba52f1cae43  <= I25c61073e64c8149ae96f3157045d317349321841e21a3d69b3baf3bd70bbd03 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 != I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[4] ) begin
                    Iac242fc0dcf37a86cc334319d77aaae46dd223017f2a6489c4e33314eabc9874  <=  ~Id156956a3b93d6a741a81c5a94e057e054ad7d4467a54a691bbd147afb30ead7 + 1;
                end else begin
                    Iac242fc0dcf37a86cc334319d77aaae46dd223017f2a6489c4e33314eabc9874  <= Id156956a3b93d6a741a81c5a94e057e054ad7d4467a54a691bbd147afb30ead7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[4] ) begin
                    Ia2417744c8f15898d5d951e15cdf8c03d932cdac6acd27e32045e0fbfbfe4f30  <=  ~Ie4eea240addf4997dde0e268e6404bea936a04629cd4d244a101a6a38e6ec03e + 1;
                end else begin
                    Ia2417744c8f15898d5d951e15cdf8c03d932cdac6acd27e32045e0fbfbfe4f30  <= Ie4eea240addf4997dde0e268e6404bea936a04629cd4d244a101a6a38e6ec03e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 != I355f4f82732333ae56692d1c7ee89b368d938d9ce1d5f806be7e46482c10e19c[0] ) begin
                    I225543794992ac9aa68ac3eeea38d41077ab5512b9f3b95fbd65a839294088e9  <=  ~I536f7bfebdfdbdfef2f9b530022a63e1a70a1ef0b344d7f34ef956bed72fc94b + 1;
                end else begin
                    I225543794992ac9aa68ac3eeea38d41077ab5512b9f3b95fbd65a839294088e9  <= I536f7bfebdfdbdfef2f9b530022a63e1a70a1ef0b344d7f34ef956bed72fc94b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[11] ) begin
                    Ibcf016cc83d0fcc2c731aa53147c199b32b3dc7a9f1a255e1a0e31615077205f  <=  ~I53a83ec9af418aeb6869bf9db2b0ce128564fcf62d2a16506906303025076ca3 + 1;
                end else begin
                    Ibcf016cc83d0fcc2c731aa53147c199b32b3dc7a9f1a255e1a0e31615077205f  <= I53a83ec9af418aeb6869bf9db2b0ce128564fcf62d2a16506906303025076ca3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[4] ) begin
                    I6e88f83ef5bc5f950a4bcb904ffede2603201e72e362aedb8db04412f7bc2bd5  <=  ~I4644d5f1dfb72ca4669b26a415cb9aeb54051fe8d28a6461d696f00bdf6c930a + 1;
                end else begin
                    I6e88f83ef5bc5f950a4bcb904ffede2603201e72e362aedb8db04412f7bc2bd5  <= I4644d5f1dfb72ca4669b26a415cb9aeb54051fe8d28a6461d696f00bdf6c930a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[8] ) begin
                    I6dc5ebe003a649f0e4106dc27f25387651d43259f0ddafad10411795ee48b40c  <=  ~Ie02a7d9471f0915572b8db6797d0ea1f2fa380d96a4e02a5783e584800e6676b + 1;
                end else begin
                    I6dc5ebe003a649f0e4106dc27f25387651d43259f0ddafad10411795ee48b40c  <= Ie02a7d9471f0915572b8db6797d0ea1f2fa380d96a4e02a5783e584800e6676b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[5] ) begin
                    I3ae1a42457a669272eeff1bc293c80c67239ef6b725a09eacb82b06ec84edd65  <=  ~I0f39af323e102d03f5089838b2b6576c03169135defb533f54e57d8450f1130e + 1;
                end else begin
                    I3ae1a42457a669272eeff1bc293c80c67239ef6b725a09eacb82b06ec84edd65  <= I0f39af323e102d03f5089838b2b6576c03169135defb533f54e57d8450f1130e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba != I9b2ce64b97ca55921bacb9b6aa4cdc8da5c1e33db4215a2470b7cfab3693576c[0] ) begin
                    Idd1dac44a6f35d558d400160a087fe7628ef80ad72c3962df2b3a3809b89bcdd  <=  ~Iaaee3c7078bf1bcda85bade0d66984c675177a0f1c66c58f47e3775916797a57 + 1;
                end else begin
                    Idd1dac44a6f35d558d400160a087fe7628ef80ad72c3962df2b3a3809b89bcdd  <= Iaaee3c7078bf1bcda85bade0d66984c675177a0f1c66c58f47e3775916797a57 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[11] ) begin
                    I544bba815490c8592dda0fd85cb612828256c09ba1431bc2632b74cc9cd2aa29  <=  ~Ifcc101725d905f243fff4a458ab8da67311d5563911d69daad960072e1927054 + 1;
                end else begin
                    I544bba815490c8592dda0fd85cb612828256c09ba1431bc2632b74cc9cd2aa29  <= Ifcc101725d905f243fff4a458ab8da67311d5563911d69daad960072e1927054 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[4] ) begin
                    I0d9bc57dbbebd429ee5a5e5dabc1cd0bd9f4de95a920346b9e61cee83969ba0f  <=  ~If5e789a890f931a53acd095741f7a5936f15da9e0007b159a3a3762ec13223f8 + 1;
                end else begin
                    I0d9bc57dbbebd429ee5a5e5dabc1cd0bd9f4de95a920346b9e61cee83969ba0f  <= If5e789a890f931a53acd095741f7a5936f15da9e0007b159a3a3762ec13223f8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[8] ) begin
                    Icac36c9706c9e063b771faf556f6699e280687be228aebf6ce71f5ae775a9754  <=  ~Ic7fa79c98c1eda80a19d8475857fb44ab41c53596b0b59806fa776d4c4ad02f4 + 1;
                end else begin
                    Icac36c9706c9e063b771faf556f6699e280687be228aebf6ce71f5ae775a9754  <= Ic7fa79c98c1eda80a19d8475857fb44ab41c53596b0b59806fa776d4c4ad02f4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[5] ) begin
                    I6d70d8c6d44eb58daff53226cbb59eb647b6dec6bed37021a64e16ac5318d484  <=  ~I6c1edf3d3971f7ab6f93e50a9500cd37fa3bb42d75c70d236f514e4c15a61f2b + 1;
                end else begin
                    I6d70d8c6d44eb58daff53226cbb59eb647b6dec6bed37021a64e16ac5318d484  <= I6c1edf3d3971f7ab6f93e50a9500cd37fa3bb42d75c70d236f514e4c15a61f2b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 != I2d78ac4a4125ec25a02df6484c0ae640a37f915383b72f33b91e87cdf376fdf7[0] ) begin
                    Ic039114ea8ac4120b09973c79fdc044251fc66bdeb18a498dd6ed7265cdfba2a  <=  ~Ic3234b24482f57a12d4db307382a5591bd66ceb0dd4bb120eadc7ab2770d003d + 1;
                end else begin
                    Ic039114ea8ac4120b09973c79fdc044251fc66bdeb18a498dd6ed7265cdfba2a  <= Ic3234b24482f57a12d4db307382a5591bd66ceb0dd4bb120eadc7ab2770d003d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[11] ) begin
                    I7530c712ec14c8fe97d1699177ef642847c5c1ce6185d1eab39b8416b562b454  <=  ~Icaa9abc6adde275d5c5011fc8cf6ead11032cc1bfc286b3a392ec507e4ff0d4c + 1;
                end else begin
                    I7530c712ec14c8fe97d1699177ef642847c5c1ce6185d1eab39b8416b562b454  <= Icaa9abc6adde275d5c5011fc8cf6ead11032cc1bfc286b3a392ec507e4ff0d4c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[4] ) begin
                    Ia9d25b6cb880b9a00c9bb27bdb80c08988eee46afccbd578659eb98301fbb8a8  <=  ~Ifc444a5134bbeeda6005a847d5ce4e180e6c809776e32d1ac709c3827d1d84b4 + 1;
                end else begin
                    Ia9d25b6cb880b9a00c9bb27bdb80c08988eee46afccbd578659eb98301fbb8a8  <= Ifc444a5134bbeeda6005a847d5ce4e180e6c809776e32d1ac709c3827d1d84b4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[8] ) begin
                    Ic02dae50f30bea04d63949eadbcf892ce936efc5373a6185668a20311dd59f4f  <=  ~I41fff62fe024b1bc1071aae30dd931c1dabf2e12d0d1cdc295bbbbd946d63358 + 1;
                end else begin
                    Ic02dae50f30bea04d63949eadbcf892ce936efc5373a6185668a20311dd59f4f  <= I41fff62fe024b1bc1071aae30dd931c1dabf2e12d0d1cdc295bbbbd946d63358 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[5] ) begin
                    I19797110801d39a7970e6d8665215c967071ad9a1bad12c33401b44f595772b7  <=  ~I8ef6ca3a27d76c9635bc942fcfb21cae619dc5b7bc842952e2a29f7f2915e62b + 1;
                end else begin
                    I19797110801d39a7970e6d8665215c967071ad9a1bad12c33401b44f595772b7  <= I8ef6ca3a27d76c9635bc942fcfb21cae619dc5b7bc842952e2a29f7f2915e62b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb != Id727bdc545af53e8f89be0ac5627d0c0c0f0bd7d75030bcb41f198a4fe9c7d64[0] ) begin
                    I21b3fa431ddc4bc8eacfb17a90fdac2bb32e4d0f4d0118715642c37601a1f883  <=  ~I1ec8e7e460c616e3d6459dd35f82ebcebdc1bd7f9680c38489e292be831ada10 + 1;
                end else begin
                    I21b3fa431ddc4bc8eacfb17a90fdac2bb32e4d0f4d0118715642c37601a1f883  <= I1ec8e7e460c616e3d6459dd35f82ebcebdc1bd7f9680c38489e292be831ada10 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[11] ) begin
                    I8b2c2b27add863ad56639a306f803b656ee8f91170e649d29aedc5321181f857  <=  ~I3c396eafe78ef3a7c94cae71c86a808a9fc88960e7519256fb1c0b54bc865334 + 1;
                end else begin
                    I8b2c2b27add863ad56639a306f803b656ee8f91170e649d29aedc5321181f857  <= I3c396eafe78ef3a7c94cae71c86a808a9fc88960e7519256fb1c0b54bc865334 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[4] ) begin
                    I1517acf28729695d689aced1c7eb358d9acfc4453fedf95a76fc22c972550c63  <=  ~I78382168abd43ba48f24ad5e574782b47afeeffe0632ae5b4aeff07ebedabf4f + 1;
                end else begin
                    I1517acf28729695d689aced1c7eb358d9acfc4453fedf95a76fc22c972550c63  <= I78382168abd43ba48f24ad5e574782b47afeeffe0632ae5b4aeff07ebedabf4f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[8] ) begin
                    I8ea9b55580c15fa584fb934e010debd92e2e893630de456e85036d583921011b  <=  ~I55de212bade4801bfd54acbc885f19f7f43fc63874f6a531f8289cccb06c81a2 + 1;
                end else begin
                    I8ea9b55580c15fa584fb934e010debd92e2e893630de456e85036d583921011b  <= I55de212bade4801bfd54acbc885f19f7f43fc63874f6a531f8289cccb06c81a2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[5] ) begin
                    I2790277776fa84c3edba2332cf538f8ea3a40c1b06cece7463a3b4757b1fe213  <=  ~Ia4c73e87649527da20616919420137fa4c1c8cfb4c85f4728a8441109168c6ad + 1;
                end else begin
                    I2790277776fa84c3edba2332cf538f8ea3a40c1b06cece7463a3b4757b1fe213  <= Ia4c73e87649527da20616919420137fa4c1c8cfb4c85f4728a8441109168c6ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 != I7661c17a1c73dbca82a6d3bfba2ab85ebb0131c1e513f093e1b0aec54907595d[0] ) begin
                    I1c6d953c9a0e96d328cc4b515867b2ac21d2947a85e96be19f38e67a8b15001c  <=  ~I04eb84d9339dab27e5615403aad9f09e40f6b123c73c8c8fd6c27f8e91ed4af6 + 1;
                end else begin
                    I1c6d953c9a0e96d328cc4b515867b2ac21d2947a85e96be19f38e67a8b15001c  <= I04eb84d9339dab27e5615403aad9f09e40f6b123c73c8c8fd6c27f8e91ed4af6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[10] ) begin
                    I4a86387a3136768ab52d320fae7fe63c7c74bb5541d18889faa263c71b2bfce6  <=  ~I49fac311626d99832accfdbaf5db0e3da11e0d89693c843295ada1310a5d8f84 + 1;
                end else begin
                    I4a86387a3136768ab52d320fae7fe63c7c74bb5541d18889faa263c71b2bfce6  <= I49fac311626d99832accfdbaf5db0e3da11e0d89693c843295ada1310a5d8f84 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[4] ) begin
                    Ia42e25bf722566321268c83de181d196619f062381c7fdb381ab5f6aeba6589b  <=  ~Ic15cf2e839052d47aa87202bae190c69e5410914d9e00120099307d6f7a663c5 + 1;
                end else begin
                    Ia42e25bf722566321268c83de181d196619f062381c7fdb381ab5f6aeba6589b  <= Ic15cf2e839052d47aa87202bae190c69e5410914d9e00120099307d6f7a663c5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[9] ) begin
                    I54296c97ecd9a699f171f4d7271c761aeea50255010a0a90d2dabc16a0cbef79  <=  ~I74677cda9719646b1c842acbed5d3b13462ef153d0a8907019b2553c808f84c6 + 1;
                end else begin
                    I54296c97ecd9a699f171f4d7271c761aeea50255010a0a90d2dabc16a0cbef79  <= I74677cda9719646b1c842acbed5d3b13462ef153d0a8907019b2553c808f84c6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681 != I553a83634252c50164bdde3576d7e1552a147490d02eac6dfd1140a46b813d08[0] ) begin
                    Ib823a58e9d4db87e4d73a81a772a02435af32a11d3c2265fb8a16021cfe4503d  <=  ~I4e0c405b4f7107ae7d9a35eff8fc48672c1ff35ede5dcbaa4340926c9d9e65d4 + 1;
                end else begin
                    Ib823a58e9d4db87e4d73a81a772a02435af32a11d3c2265fb8a16021cfe4503d  <= I4e0c405b4f7107ae7d9a35eff8fc48672c1ff35ede5dcbaa4340926c9d9e65d4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[10] ) begin
                    I345c0aef41ee2863a96a076a78d92c7498f50ef90e82e75565df1d1f38a08161  <=  ~I1db1a5d4e476af4fb7bbf80331760238438096833616b30904a4b6fbe0057e63 + 1;
                end else begin
                    I345c0aef41ee2863a96a076a78d92c7498f50ef90e82e75565df1d1f38a08161  <= I1db1a5d4e476af4fb7bbf80331760238438096833616b30904a4b6fbe0057e63 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1 != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[4] ) begin
                    Ibca01267ba9d7e2fe9f8df34a548836390ba12b9b782f16ba40965c00735213a  <=  ~I083b6e833d8b3bda9d56f159a5e297305e44fad9f2024a3204c6e5b7afca9405 + 1;
                end else begin
                    Ibca01267ba9d7e2fe9f8df34a548836390ba12b9b782f16ba40965c00735213a  <= I083b6e833d8b3bda9d56f159a5e297305e44fad9f2024a3204c6e5b7afca9405 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[9] ) begin
                    Ic36cf3da50983e4168cc0a31ec0a86c171714355c0fab18398b8daf57bee1a45  <=  ~I410bc8d9b13d79713c47cab785cae1ee4db55ba3e7a207519bdbc646dfa815dc + 1;
                end else begin
                    Ic36cf3da50983e4168cc0a31ec0a86c171714355c0fab18398b8daf57bee1a45  <= I410bc8d9b13d79713c47cab785cae1ee4db55ba3e7a207519bdbc646dfa815dc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1 != Ib450c1ee41d04516060a410bbdfb605f0ce13cd8781596ce5218928ed207de8a[0] ) begin
                    I3427390162b0952481e5f0728a20075c9cfb814431ecbb1a4014d407ab3b3afd  <=  ~Iab1ad3fda6ef48c15a116045600ab96f057c4e2769b1736742ece54e049a9884 + 1;
                end else begin
                    I3427390162b0952481e5f0728a20075c9cfb814431ecbb1a4014d407ab3b3afd  <= Iab1ad3fda6ef48c15a116045600ab96f057c4e2769b1736742ece54e049a9884 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[10] ) begin
                    Ia7900b5a01cfc1c4db79ca653f072956c13e2040cbd94cf07de2f1d969222fa8  <=  ~If01282d291c85bcab01b47104be9ed13915609c85c61d979b60b02847a685e4f + 1;
                end else begin
                    Ia7900b5a01cfc1c4db79ca653f072956c13e2040cbd94cf07de2f1d969222fa8  <= If01282d291c85bcab01b47104be9ed13915609c85c61d979b60b02847a685e4f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851 != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[4] ) begin
                    I783b89f0c1e5463646e0fceb976f2b27aac523a677eff6e597e434672b0daac1  <=  ~I2c3551c0a960cbdcab2b802148c759ca7c8dc401d98b251d9ea21d6de16d3bf8 + 1;
                end else begin
                    I783b89f0c1e5463646e0fceb976f2b27aac523a677eff6e597e434672b0daac1  <= I2c3551c0a960cbdcab2b802148c759ca7c8dc401d98b251d9ea21d6de16d3bf8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[9] ) begin
                    I238a5c9cd1dcce0d745817081a4b240f74de3de6f18a3abcc42cafbb19a0ad69  <=  ~Ic7977549066f72a2e4c0d91c592a5d93a2a64fd1ac48cafd6f0f4600912f3fc1 + 1;
                end else begin
                    I238a5c9cd1dcce0d745817081a4b240f74de3de6f18a3abcc42cafbb19a0ad69  <= Ic7977549066f72a2e4c0d91c592a5d93a2a64fd1ac48cafd6f0f4600912f3fc1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851 != Ica745abd4de790f1cd3e2a5a32a9d0b5edf1b64e85759c49f3b4e51779443709[0] ) begin
                    I35a9ae1cf23d8697091de65a1d0678632bd6889ae32408d7658e542a756e95ca  <=  ~I08c54adda4326fbc5985605f17f5b1c47ce821476ba25053aaa7449a571bf33c + 1;
                end else begin
                    I35a9ae1cf23d8697091de65a1d0678632bd6889ae32408d7658e542a756e95ca  <= I08c54adda4326fbc5985605f17f5b1c47ce821476ba25053aaa7449a571bf33c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[10] ) begin
                    I9eb30c75f8d71ade925633d7c8bc6b948ae519cdff33ddb885761bf72a8b0869  <=  ~I74a65dbb33c6088646be4339ced1e6167ed3c67fe3f520e10d4fb2c96358ce62 + 1;
                end else begin
                    I9eb30c75f8d71ade925633d7c8bc6b948ae519cdff33ddb885761bf72a8b0869  <= I74a65dbb33c6088646be4339ced1e6167ed3c67fe3f520e10d4fb2c96358ce62 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104 != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[4] ) begin
                    I64aaf806ebf0ead2a4836251dccd62a394b984823592340be94f4ea02e12d766  <=  ~I378dc69acacc690da268354f08a9f1fd08b11a899cd2253c2cca3c979245a06b + 1;
                end else begin
                    I64aaf806ebf0ead2a4836251dccd62a394b984823592340be94f4ea02e12d766  <= I378dc69acacc690da268354f08a9f1fd08b11a899cd2253c2cca3c979245a06b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[9] ) begin
                    I8b3bb7a4701d3ef22c71a9631482e13afc2ff80f40e2f0ae75cb2211af5ce6d9  <=  ~I8519733c2d4de3643ecf515bc788e665d7661c947a6532dcefce59b255fc05c5 + 1;
                end else begin
                    I8b3bb7a4701d3ef22c71a9631482e13afc2ff80f40e2f0ae75cb2211af5ce6d9  <= I8519733c2d4de3643ecf515bc788e665d7661c947a6532dcefce59b255fc05c5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104 != I6399b29558311ea40cda1388848ce13bb7593bfed01ca2a10fa5d8ed6700df56[0] ) begin
                    I37e54e8ae28cf1a36cb9101d5afd4d523ca9a6ae244efe641c547a4114726bea  <=  ~I2b3f1cb9e25ac68c67abdee581e7dbb74b039b9f1f04459e3a4049769f27c474 + 1;
                end else begin
                    I37e54e8ae28cf1a36cb9101d5afd4d523ca9a6ae244efe641c547a4114726bea  <= I2b3f1cb9e25ac68c67abdee581e7dbb74b039b9f1f04459e3a4049769f27c474 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[12] ) begin
                    I7e7be31550be1cacb2acdb27d5120769dd7a0a49efb833051ceb83c8cf691e21  <=  ~Id79e7da27c2a195d433419bcc0481ffe12155390f0a10ac6be75723cf2ad53f2 + 1;
                end else begin
                    I7e7be31550be1cacb2acdb27d5120769dd7a0a49efb833051ceb83c8cf691e21  <= Id79e7da27c2a195d433419bcc0481ffe12155390f0a10ac6be75723cf2ad53f2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[5] ) begin
                    I86e764dc3320206d9b52013c2d735ff4d27bf6e4a82227486e64b4ceb68dfe8a  <=  ~I9aa3880979a20743da2aa753686d0ecaf0702008920d80af34d834ef1e2249be + 1;
                end else begin
                    I86e764dc3320206d9b52013c2d735ff4d27bf6e4a82227486e64b4ceb68dfe8a  <= I9aa3880979a20743da2aa753686d0ecaf0702008920d80af34d834ef1e2249be ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[10] ) begin
                    I6a24b9c3ea194d09d619dff007c4c6f53a3cbbbae5c9d3ba718bc3546eaad989  <=  ~Ie591b9c2c777632b671f8aa86f6befb3d02e16c23329cbc7c07438588aea4c9b + 1;
                end else begin
                    I6a24b9c3ea194d09d619dff007c4c6f53a3cbbbae5c9d3ba718bc3546eaad989  <= Ie591b9c2c777632b671f8aa86f6befb3d02e16c23329cbc7c07438588aea4c9b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[3] ) begin
                    Ia244be7d571a1e41348c37534a23f7cc942b689cbcd5dff8c10043325b80e322  <=  ~Ibaccfedeb751c2506a2342df2f75fe492accc5c68614fcb90b4f5c332c088808 + 1;
                end else begin
                    Ia244be7d571a1e41348c37534a23f7cc942b689cbcd5dff8c10043325b80e322  <= Ibaccfedeb751c2506a2342df2f75fe492accc5c68614fcb90b4f5c332c088808 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f != I6f529a4dd77f75d9af4350baf53ba61c1e9c5ea6227c26690987d244dfe71528[0] ) begin
                    I9544a194d3d75c6c414169ea2536e111c09711ee602eb3462c4022350906a21e  <=  ~Ifa134df77ff670a0cb559c384c786af4de916cea66ca13147d43f4030d474d0f + 1;
                end else begin
                    I9544a194d3d75c6c414169ea2536e111c09711ee602eb3462c4022350906a21e  <= Ifa134df77ff670a0cb559c384c786af4de916cea66ca13147d43f4030d474d0f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[12] ) begin
                    I7b8225b7ff4972426858a8550dc67a231d85fe94426bf0812906f1aee0e2d097  <=  ~Ib378be3532348ccba868d918209ee3f013c1844044c8a93467a93c3463f7a36c + 1;
                end else begin
                    I7b8225b7ff4972426858a8550dc67a231d85fe94426bf0812906f1aee0e2d097  <= Ib378be3532348ccba868d918209ee3f013c1844044c8a93467a93c3463f7a36c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[5] ) begin
                    I9bcd5f3f4630ce7a24ea4479c9ddfce59ed809dfaad9d767e80295c41b332f4a  <=  ~Ib85e84ee2add613edb76e2321f7a5d6b4de3be9b1ab97905b5980277ed273dd1 + 1;
                end else begin
                    I9bcd5f3f4630ce7a24ea4479c9ddfce59ed809dfaad9d767e80295c41b332f4a  <= Ib85e84ee2add613edb76e2321f7a5d6b4de3be9b1ab97905b5980277ed273dd1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[10] ) begin
                    I50a310ea41e0637bf28b5f56cf11560bc936e15c73acee063c60668bfa905fed  <=  ~I10ee9fd16ea681268e4bcdcc30b515d990dc30d3fd41e059e9f1dcc80042ae1f + 1;
                end else begin
                    I50a310ea41e0637bf28b5f56cf11560bc936e15c73acee063c60668bfa905fed  <= I10ee9fd16ea681268e4bcdcc30b515d990dc30d3fd41e059e9f1dcc80042ae1f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[3] ) begin
                    I6b264ac5221269381b155a30c051523f4488ecdc6eb2cf60da80a8b84c49bd96  <=  ~Ic33e33bdd936748553ff29221e983dc115121fc84bd1a2799a3da8120be82c04 + 1;
                end else begin
                    I6b264ac5221269381b155a30c051523f4488ecdc6eb2cf60da80a8b84c49bd96  <= Ic33e33bdd936748553ff29221e983dc115121fc84bd1a2799a3da8120be82c04 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd != I7a94e46f1351801c2edf76bf3b70e3b5100b8e6108d60d9341591aa59f4e95d1[0] ) begin
                    I1e4bc72a55efb8462410905dcb2c9a8412e2533ded854d23ca648e0e36802960  <=  ~I0705a3be469f22a69c0c4d2366fd0eaee02065685349db5abd81049530fbf842 + 1;
                end else begin
                    I1e4bc72a55efb8462410905dcb2c9a8412e2533ded854d23ca648e0e36802960  <= I0705a3be469f22a69c0c4d2366fd0eaee02065685349db5abd81049530fbf842 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[12] ) begin
                    I41b365f8c613bf86dc5e2ed41719ec6823046127babf87a083503ebcfd38ae75  <=  ~Ic0edcffe7bf2caf311b42675297cde79af81c022f660757cdbed53dbf5c04eaf + 1;
                end else begin
                    I41b365f8c613bf86dc5e2ed41719ec6823046127babf87a083503ebcfd38ae75  <= Ic0edcffe7bf2caf311b42675297cde79af81c022f660757cdbed53dbf5c04eaf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[5] ) begin
                    I15123100f4377e14c62cf47fb1fb652badc3bd0e8f0ab4b970a0bece065a6380  <=  ~I600367d873f901e6b7f92a4f9c0ac92c9f8efa6da1d6e6945f83b863e8bb8519 + 1;
                end else begin
                    I15123100f4377e14c62cf47fb1fb652badc3bd0e8f0ab4b970a0bece065a6380  <= I600367d873f901e6b7f92a4f9c0ac92c9f8efa6da1d6e6945f83b863e8bb8519 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[10] ) begin
                    I7469c1791d81d0924eb0faa6303565dc78fe9eb371fa13039ff89b92b7f51a6b  <=  ~I8e30a7f3eb36b84c9df9d59f6164c757c8612fb12567ddfd03c32388af750bb6 + 1;
                end else begin
                    I7469c1791d81d0924eb0faa6303565dc78fe9eb371fa13039ff89b92b7f51a6b  <= I8e30a7f3eb36b84c9df9d59f6164c757c8612fb12567ddfd03c32388af750bb6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[3] ) begin
                    I8d8dbd62189397b5e9189ead2126a615d5b6cea393901e21cd89c255d6672615  <=  ~I8d123ed314ee10c10f04151727cd5ce1e836c01f0f8143285b54425633591008 + 1;
                end else begin
                    I8d8dbd62189397b5e9189ead2126a615d5b6cea393901e21cd89c255d6672615  <= I8d123ed314ee10c10f04151727cd5ce1e836c01f0f8143285b54425633591008 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 != I0b761d71a88d70e6228dcf7325206f840d9da85892ba151c317e06079291fc2e[0] ) begin
                    If2cec64e868d25d7fbad45ce4889c6a4cac0084aae00d2aa8963678edbb88875  <=  ~I0ae31ee6a1c597ec90ca13dd69a651079d801c279292523953428af55188ddea + 1;
                end else begin
                    If2cec64e868d25d7fbad45ce4889c6a4cac0084aae00d2aa8963678edbb88875  <= I0ae31ee6a1c597ec90ca13dd69a651079d801c279292523953428af55188ddea ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[12] ) begin
                    Ie3290070e785df28e64ff4df124d14c370c9edb924d5f35b059a6c82e8373f91  <=  ~I7bbfdff59068ad7e527ada31d96fd47cb737e6b7ba56b1b2b9e522fe3a63a954 + 1;
                end else begin
                    Ie3290070e785df28e64ff4df124d14c370c9edb924d5f35b059a6c82e8373f91  <= I7bbfdff59068ad7e527ada31d96fd47cb737e6b7ba56b1b2b9e522fe3a63a954 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[5] ) begin
                    Ia9bf10fecfe62530ea6be4687ecf78a2ac08c6fc6e38328c2d64a80cb5a3d72b  <=  ~I09001eb04237069c413098f07bb41538c6d39b0ac000f175d61ee3c0b47cfae2 + 1;
                end else begin
                    Ia9bf10fecfe62530ea6be4687ecf78a2ac08c6fc6e38328c2d64a80cb5a3d72b  <= I09001eb04237069c413098f07bb41538c6d39b0ac000f175d61ee3c0b47cfae2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[10] ) begin
                    I53c29303c76ac3c1c02fc9a74eaff9595153ba06d67c08e07790c58e53b674f1  <=  ~Iddcd6e6693d5f625ba82ec2cdb0a93ca1826dca4989d19221c8127513648eab2 + 1;
                end else begin
                    I53c29303c76ac3c1c02fc9a74eaff9595153ba06d67c08e07790c58e53b674f1  <= Iddcd6e6693d5f625ba82ec2cdb0a93ca1826dca4989d19221c8127513648eab2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[3] ) begin
                    I468b28bee4fe1c0d20fe7abd9338bf844ce0a2e322ed6b6de11e2ac621572c48  <=  ~I89df294963327dee66a931b858b05dddd97e3fe4d048ecbfaa9c15e28c57602e + 1;
                end else begin
                    I468b28bee4fe1c0d20fe7abd9338bf844ce0a2e322ed6b6de11e2ac621572c48  <= I89df294963327dee66a931b858b05dddd97e3fe4d048ecbfaa9c15e28c57602e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 != Ic2ae521a3a6fef956f28a89da365b0838d535c9f7801a405cf60cc776ba0af2a[0] ) begin
                    I73ad61911b0822e313aab2c484d1699cf2655a42a2bb0a1c9ab36228e41d0f7f  <=  ~I1f0110f45df674628a1a02cf01dc58577628dd88049b93ebf02b5c4143781ade + 1;
                end else begin
                    I73ad61911b0822e313aab2c484d1699cf2655a42a2bb0a1c9ab36228e41d0f7f  <= I1f0110f45df674628a1a02cf01dc58577628dd88049b93ebf02b5c4143781ade ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[13] ) begin
                    I02ed3128371185efeae1e27046aa378006ec78d7c458dcba137f69c29c4363bc  <=  ~Ib0995588ac28564326a4dec88344ddd733075750fab9f4f8fec64cc91b3b48e2 + 1;
                end else begin
                    I02ed3128371185efeae1e27046aa378006ec78d7c458dcba137f69c29c4363bc  <= Ib0995588ac28564326a4dec88344ddd733075750fab9f4f8fec64cc91b3b48e2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[5] ) begin
                    I4a6a17ada186c2bb60e521443c0a5a0248d03242c4ae01b751fcce4abe853065  <=  ~I3a2ddd5962242d66fa4b8bca39a81765dfbc6c0b6b012ee42329dcdfc12ae9b3 + 1;
                end else begin
                    I4a6a17ada186c2bb60e521443c0a5a0248d03242c4ae01b751fcce4abe853065  <= I3a2ddd5962242d66fa4b8bca39a81765dfbc6c0b6b012ee42329dcdfc12ae9b3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[11] ) begin
                    I9b8a4dcee9668bb71803c25e0ece0eebbf704eb29cfa7b91c47cf48d61076803  <=  ~I83cd839beef638f212312a0093595ec3d71dc80e240aba892f6404de6d614bec + 1;
                end else begin
                    I9b8a4dcee9668bb71803c25e0ece0eebbf704eb29cfa7b91c47cf48d61076803  <= I83cd839beef638f212312a0093595ec3d71dc80e240aba892f6404de6d614bec ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[4] ) begin
                    Ie79db7f22cab9cd57482ce0141d83d5c1ff720a7c3dca2c3664feb4a1e2f4850  <=  ~I3420837ce14103293c9ee75848088cd144ed5b975add2adfd479ad10eff552ca + 1;
                end else begin
                    Ie79db7f22cab9cd57482ce0141d83d5c1ff720a7c3dca2c3664feb4a1e2f4850  <= I3420837ce14103293c9ee75848088cd144ed5b975add2adfd479ad10eff552ca ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa != I01d9f8a8900be1981c601c0ccb45c1f39a0fdc16179245d80fbb2ad6d7060899[0] ) begin
                    I218255d96e659dc8f60cddd40cac94a56d93556ed609b60157d88b298ec95f0c  <=  ~I641204b71e0368d174adf904e08c12465fc7a18e1adf1372e1649efad206ba0a + 1;
                end else begin
                    I218255d96e659dc8f60cddd40cac94a56d93556ed609b60157d88b298ec95f0c  <= I641204b71e0368d174adf904e08c12465fc7a18e1adf1372e1649efad206ba0a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[13] ) begin
                    I26d08096b43367ba37b8f6dcd919bf4ecb9c660a39f2c0ae29f655e42b88887a  <=  ~I10bd3ad7827da7bbb0e1170d7e495b88ab6ac55e0421b4f208f5c1ccd722198d + 1;
                end else begin
                    I26d08096b43367ba37b8f6dcd919bf4ecb9c660a39f2c0ae29f655e42b88887a  <= I10bd3ad7827da7bbb0e1170d7e495b88ab6ac55e0421b4f208f5c1ccd722198d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[5] ) begin
                    Ibe932d914d189b275138de8d6f3ffb914940d4b2bbecb574fba3c6aed885c44e  <=  ~Iee26e4077668d0e7329068693c4279480b26e4f16adb0161c8e7f87de802a14a + 1;
                end else begin
                    Ibe932d914d189b275138de8d6f3ffb914940d4b2bbecb574fba3c6aed885c44e  <= Iee26e4077668d0e7329068693c4279480b26e4f16adb0161c8e7f87de802a14a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[11] ) begin
                    Ia92993e9a66294adf7a4dbe1ea88a9e8be6367da1c05b8df343b3c7a38bfd8b6  <=  ~Ia8e573753ddee4fe18b1f9fbafcd135efc7fb7e7eec52e45b5148b0dcf346050 + 1;
                end else begin
                    Ia92993e9a66294adf7a4dbe1ea88a9e8be6367da1c05b8df343b3c7a38bfd8b6  <= Ia8e573753ddee4fe18b1f9fbafcd135efc7fb7e7eec52e45b5148b0dcf346050 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[4] ) begin
                    I08c55e08731cbdc9703e607b481a65177e7e1e242fdab9bfb014964bb0d1d22c  <=  ~Ie8e89070910f06608a4df5951936faf465b4f235d92b3cf8a3820d03bcaa83ed + 1;
                end else begin
                    I08c55e08731cbdc9703e607b481a65177e7e1e242fdab9bfb014964bb0d1d22c  <= Ie8e89070910f06608a4df5951936faf465b4f235d92b3cf8a3820d03bcaa83ed ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe != Icdfc2f0ce24f01af7df8a99b58de3a74e1dda0eea5b41ff2c342106cb226abdc[0] ) begin
                    I11284a18d6115421b4c76054c1a580c41987dec66caa7d5bd9107bbd4ac8bc2c  <=  ~I1a0b36a215887b4419ebcfbddb0ab8b4b9b21c4643051db135c9d9ee53c6bb3e + 1;
                end else begin
                    I11284a18d6115421b4c76054c1a580c41987dec66caa7d5bd9107bbd4ac8bc2c  <= I1a0b36a215887b4419ebcfbddb0ab8b4b9b21c4643051db135c9d9ee53c6bb3e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[13] ) begin
                    I3358739f5e55263208e661a339d6b29f188f07ef07e2ee7a63a24011a4f8568f  <=  ~I84694b26e240bcc3e7c9b224ce3c2f5891fb546a4fc11e4597819fd9827c3105 + 1;
                end else begin
                    I3358739f5e55263208e661a339d6b29f188f07ef07e2ee7a63a24011a4f8568f  <= I84694b26e240bcc3e7c9b224ce3c2f5891fb546a4fc11e4597819fd9827c3105 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[5] ) begin
                    I377aa224e1817d2ab5cb02a5a290a723621782607fcd59b319d8cec1b092bc1b  <=  ~Ie69f3ad2e3dcb172e525302a533963ab9a2a08af8d1ec71e07d0946d393c056f + 1;
                end else begin
                    I377aa224e1817d2ab5cb02a5a290a723621782607fcd59b319d8cec1b092bc1b  <= Ie69f3ad2e3dcb172e525302a533963ab9a2a08af8d1ec71e07d0946d393c056f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[11] ) begin
                    Ic7af968d25c444d210ebbc7ae563688f4f8a48f38035ce5bccee100e10555047  <=  ~I6e0e1c5361317aa91a6e54e23fe2585744a1ec47fcb2412ed152b660781c7832 + 1;
                end else begin
                    Ic7af968d25c444d210ebbc7ae563688f4f8a48f38035ce5bccee100e10555047  <= I6e0e1c5361317aa91a6e54e23fe2585744a1ec47fcb2412ed152b660781c7832 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[4] ) begin
                    I14730b2825dc07428388347472491ef3abe06da3bcea9b7dc9c919079c22325c  <=  ~Ia338a53ab734049efb28655e209908f1fd2c5d19f8056463d711cc1e50dde602 + 1;
                end else begin
                    I14730b2825dc07428388347472491ef3abe06da3bcea9b7dc9c919079c22325c  <= Ia338a53ab734049efb28655e209908f1fd2c5d19f8056463d711cc1e50dde602 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 != I929ef5474f10c76c4686fb044b2833b6ba1571f2e1c82b6d92cfaadfa44946e6[0] ) begin
                    I8516ef195e4ba8f6e29a02ab5ea349a26bb68f6ebb4da847d56c03c942e9c20c  <=  ~If63dbf3e3c6000184af28e72b5f2960f6a376f509d5693a96d2ab9f92ae7b237 + 1;
                end else begin
                    I8516ef195e4ba8f6e29a02ab5ea349a26bb68f6ebb4da847d56c03c942e9c20c  <= If63dbf3e3c6000184af28e72b5f2960f6a376f509d5693a96d2ab9f92ae7b237 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[13] ) begin
                    If9bd4d7f3740f15bdf597de00eecf1cbf2e3b4efdbacbbad889c0946a6b34a24  <=  ~Ib89d5800576f979f189d88e7976f8d49b8470bcbf6b365f7cc6031735e3adb4a + 1;
                end else begin
                    If9bd4d7f3740f15bdf597de00eecf1cbf2e3b4efdbacbbad889c0946a6b34a24  <= Ib89d5800576f979f189d88e7976f8d49b8470bcbf6b365f7cc6031735e3adb4a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[5] ) begin
                    Icd30277c9d839d833f27f571231dd138497796d3e7818460d836a48b87e34d03  <=  ~I622321198c6f868e554b595d1e1616dd63ad46a80c33bbe896df9b6558418ccc + 1;
                end else begin
                    Icd30277c9d839d833f27f571231dd138497796d3e7818460d836a48b87e34d03  <= I622321198c6f868e554b595d1e1616dd63ad46a80c33bbe896df9b6558418ccc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[11] ) begin
                    I25d2b0d3ff7f684e508a62271f3d29c729dc46478248627013dd91075f8d2146  <=  ~Iafcf26b8f2df7719a0b660b41de28c5a325e50d75382579e53aa9d065bd81cbf + 1;
                end else begin
                    I25d2b0d3ff7f684e508a62271f3d29c729dc46478248627013dd91075f8d2146  <= Iafcf26b8f2df7719a0b660b41de28c5a325e50d75382579e53aa9d065bd81cbf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[4] ) begin
                    I5c3a945e8bd4c55e9cb38d19100b13668bd652bc1162d16b30f1562a6595a032  <=  ~I859639da611c77242efe899343358a650652277ea45277d9792b619196c66a1a + 1;
                end else begin
                    I5c3a945e8bd4c55e9cb38d19100b13668bd652bc1162d16b30f1562a6595a032  <= I859639da611c77242efe899343358a650652277ea45277d9792b619196c66a1a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 != I55312932ff9d69c8ffa1e42efdb5e775ccb21a8f9e8791b080b67654462e537a[0] ) begin
                    I2411dfbbf605c7590bc678373dd20b7241356a433756332f9a3445ba8dad57fb  <=  ~I2899ec4e420edc766050ec0042965f87c79455271a54ba7c947e94d37450a033 + 1;
                end else begin
                    I2411dfbbf605c7590bc678373dd20b7241356a433756332f9a3445ba8dad57fb  <= I2899ec4e420edc766050ec0042965f87c79455271a54ba7c947e94d37450a033 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[11] ) begin
                    Ifb94a220081758ce91634fef64be084898a662f7c0e8cc9f86859bf3852b3efe  <=  ~Ibb256fb3d4bbe6ddc65378ced36e01255d8164d29755891e06fbd4caf2a290cf + 1;
                end else begin
                    Ifb94a220081758ce91634fef64be084898a662f7c0e8cc9f86859bf3852b3efe  <= Ibb256fb3d4bbe6ddc65378ced36e01255d8164d29755891e06fbd4caf2a290cf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995 != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[5] ) begin
                    I91716015389a9d3b1d0cc77327f439e02e54be0d3524b2cdbeed886eea673b10  <=  ~I60f4bae66121b814e2faa564c162bccbd2ef0a73bcaf10c3c78e30ff2edcde4a + 1;
                end else begin
                    I91716015389a9d3b1d0cc77327f439e02e54be0d3524b2cdbeed886eea673b10  <= I60f4bae66121b814e2faa564c162bccbd2ef0a73bcaf10c3c78e30ff2edcde4a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[7] ) begin
                    I35e7fd3f09acca79a1003b0a4b7ac62c4a2be93bcf333abbfb13a5eefd7d5eaf  <=  ~Iac70da997560fcd3949fde686e6f8a3dc834a2ab7ff2beaeedf7614710bbfaff + 1;
                end else begin
                    I35e7fd3f09acca79a1003b0a4b7ac62c4a2be93bcf333abbfb13a5eefd7d5eaf  <= Iac70da997560fcd3949fde686e6f8a3dc834a2ab7ff2beaeedf7614710bbfaff ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995 != Icbdbaf4eb2f30bb78db34a582e06dc91689b9eab2f8fdfe4fbfb41a8cce93ca5[0] ) begin
                    I69d896cdb2303b99b73c4d6886f2686381230feca86c62fc064a85e4d11266f4  <=  ~Ie32e4f67efcbea2f033a66104b3315b46a1c857781ac63283f4d955384bcdd4f + 1;
                end else begin
                    I69d896cdb2303b99b73c4d6886f2686381230feca86c62fc064a85e4d11266f4  <= Ie32e4f67efcbea2f033a66104b3315b46a1c857781ac63283f4d955384bcdd4f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[11] ) begin
                    I1aa136009f34c39a8dbc39b4444642cd09c9cd2f01bd6310287d4ddc9bedad85  <=  ~I4720d84525310ad5428da40677f1cd99365d1467c29d214ab4ae300277322cbe + 1;
                end else begin
                    I1aa136009f34c39a8dbc39b4444642cd09c9cd2f01bd6310287d4ddc9bedad85  <= I4720d84525310ad5428da40677f1cd99365d1467c29d214ab4ae300277322cbe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2 != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[5] ) begin
                    Ied710d5ba03554d4103468029a9d895c25c10765b6e3d73bbdebc54d7cc7d8db  <=  ~Ia1f10017528e76925426be916c558186f2196a0c4d7520e57e0895e14e7c1d53 + 1;
                end else begin
                    Ied710d5ba03554d4103468029a9d895c25c10765b6e3d73bbdebc54d7cc7d8db  <= Ia1f10017528e76925426be916c558186f2196a0c4d7520e57e0895e14e7c1d53 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[7] ) begin
                    Ice24cd0bd76a7d12a0199df195b34f41f7f72f037177656693b3154d102ba729  <=  ~I46a3710c0e472a92b83354b668ac21c775b2c4e3dceadc49dc0cb712c08c319e + 1;
                end else begin
                    Ice24cd0bd76a7d12a0199df195b34f41f7f72f037177656693b3154d102ba729  <= I46a3710c0e472a92b83354b668ac21c775b2c4e3dceadc49dc0cb712c08c319e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2 != Ifa4cbbd5c3ab5e47a7d5135e4dbaf365e79c4c6a806bfae88c9c0e1c9ffe2fa5[0] ) begin
                    If6ca882e537cdf5f458a2e11b7a11f057a3d2a00923825fe236afa0b0e1442c0  <=  ~I594b73c43f22c1cc15daf1eb602be4366502100a0ad3a3bad7b7992c9839dbbb + 1;
                end else begin
                    If6ca882e537cdf5f458a2e11b7a11f057a3d2a00923825fe236afa0b0e1442c0  <= I594b73c43f22c1cc15daf1eb602be4366502100a0ad3a3bad7b7992c9839dbbb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[11] ) begin
                    I5456c559bdce4d65af540e4c71c19e44227c62e5c129b7de968ac7f311dd76f4  <=  ~Id6264ccfced253e14f1f9be10f967d475695838c367808b97abbd7578447179a + 1;
                end else begin
                    I5456c559bdce4d65af540e4c71c19e44227c62e5c129b7de968ac7f311dd76f4  <= Id6264ccfced253e14f1f9be10f967d475695838c367808b97abbd7578447179a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218 != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[5] ) begin
                    I8ca8dfb7a3a8ecb9eac34d1d1ef4768d31b86a757cb7b9ce61ef159816ceea7f  <=  ~Ied0e2037bbb2f2b7d0cef3d7d3f5b7123c006255cb7f2297df7e1a1eb03dee16 + 1;
                end else begin
                    I8ca8dfb7a3a8ecb9eac34d1d1ef4768d31b86a757cb7b9ce61ef159816ceea7f  <= Ied0e2037bbb2f2b7d0cef3d7d3f5b7123c006255cb7f2297df7e1a1eb03dee16 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[7] ) begin
                    Iab97067540ba8c9551711cdbff0c6aa3993534d3e8b352bda090a0997c681afa  <=  ~Ica6a39f57caae5761078aaf00587554f1acef5d9b2e1fb73931f5715ebc762dc + 1;
                end else begin
                    Iab97067540ba8c9551711cdbff0c6aa3993534d3e8b352bda090a0997c681afa  <= Ica6a39f57caae5761078aaf00587554f1acef5d9b2e1fb73931f5715ebc762dc ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218 != I2341907334935e19ef0e392216e39bb35c215730c464a85c0e1b804b364b492c[0] ) begin
                    Ie35443efbbf821e07284652a4b37347c4cfb959495dafa4fd2f81ffa2edc56db  <=  ~I0fe26cc77a5b117d82b8f0da27f4cc5e9465360eba32d35aeefc16ff600ad5f2 + 1;
                end else begin
                    Ie35443efbbf821e07284652a4b37347c4cfb959495dafa4fd2f81ffa2edc56db  <= I0fe26cc77a5b117d82b8f0da27f4cc5e9465360eba32d35aeefc16ff600ad5f2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[11] ) begin
                    Ia0c4bcb29e2939b889fb7a5a7b62b49a3eeb3ee6f4555518c9059cb34dfebc7a  <=  ~I8bfbee6346d016ff8cd0ef681e0efdf28d0f27b3e887397fa1aff647739e25a1 + 1;
                end else begin
                    Ia0c4bcb29e2939b889fb7a5a7b62b49a3eeb3ee6f4555518c9059cb34dfebc7a  <= I8bfbee6346d016ff8cd0ef681e0efdf28d0f27b3e887397fa1aff647739e25a1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[5] ) begin
                    I7ff25e517e328eda581e7637a2114a7cffe873df520114410c0487e503c01aa6  <=  ~I57f07e2955da5218122f614720d5890af9d7b5ac4f033e9d1c10db08e7ad1882 + 1;
                end else begin
                    I7ff25e517e328eda581e7637a2114a7cffe873df520114410c0487e503c01aa6  <= I57f07e2955da5218122f614720d5890af9d7b5ac4f033e9d1c10db08e7ad1882 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[7] ) begin
                    Ia1d4bd5d90332afbfaaac3cd0d8f5fcbc626ec4adbb0b0f16fc80923925f703f  <=  ~I9c71f3f968f3265215ce730a5f922db81aa408218fc76de3b64ee4f9396d3f78 + 1;
                end else begin
                    Ia1d4bd5d90332afbfaaac3cd0d8f5fcbc626ec4adbb0b0f16fc80923925f703f  <= I9c71f3f968f3265215ce730a5f922db81aa408218fc76de3b64ee4f9396d3f78 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a != Ic0bbaf8314688690b5a15a5613ab149f604a8bfb92a2b9ed014e7ce2757d0743[0] ) begin
                    Id6d0b1fe00e5324e0ed7c37d41ee3e848f9c7dcfb4a85f5da2b82ed4d8942b21  <=  ~I3afdbbfca5c952e1800c1e15ca629173eac62810b6bf8097421addeae979ca81 + 1;
                end else begin
                    Id6d0b1fe00e5324e0ed7c37d41ee3e848f9c7dcfb4a85f5da2b82ed4d8942b21  <= I3afdbbfca5c952e1800c1e15ca629173eac62810b6bf8097421addeae979ca81 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[12] ) begin
                    I3de9fbe37d08009f5fa66bf7c59debe7da836dc078e212968afdc608b100e3bd  <=  ~Ie9d906bda89623d793bc65968cd86bd0c63458c7a6b12fd38f7054069dfcd132 + 1;
                end else begin
                    I3de9fbe37d08009f5fa66bf7c59debe7da836dc078e212968afdc608b100e3bd  <= Ie9d906bda89623d793bc65968cd86bd0c63458c7a6b12fd38f7054069dfcd132 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[14] ) begin
                    I5eff39d324b6a8910fad41786d651086c622d331987e649ba4b3baae11ca40ce  <=  ~I969b9fa05c651f6e2f2dc426e35c43864f9b5c6d4f6278b0f7ec4e7c5e872eec + 1;
                end else begin
                    I5eff39d324b6a8910fad41786d651086c622d331987e649ba4b3baae11ca40ce  <= I969b9fa05c651f6e2f2dc426e35c43864f9b5c6d4f6278b0f7ec4e7c5e872eec ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[5] ) begin
                    Ib0ee967a174d7c841ebe71e144d6303bfc80a6083ff6ad745c76d488dea66d9e  <=  ~I436c98ccee6d1a138f1c47ef4e5b7ac39db15122b2b134828b257dd629e310a5 + 1;
                end else begin
                    Ib0ee967a174d7c841ebe71e144d6303bfc80a6083ff6ad745c76d488dea66d9e  <= I436c98ccee6d1a138f1c47ef4e5b7ac39db15122b2b134828b257dd629e310a5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e != I19ff0bebf62a994a2b5814ea41289f72cd62a38d2f37dc0027beb0f488926d4f[0] ) begin
                    I0a309e8aa7f7e07abd837c99be6d8bb8c29dc1679b449111a02f49442d5cb432  <=  ~Ide4ad5678bce6a696f0c6cb163eaf670c47c2506acf7977c1031c6ec03e03a58 + 1;
                end else begin
                    I0a309e8aa7f7e07abd837c99be6d8bb8c29dc1679b449111a02f49442d5cb432  <= Ide4ad5678bce6a696f0c6cb163eaf670c47c2506acf7977c1031c6ec03e03a58 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[12] ) begin
                    I5f1b294a0702ab37f94304ae67fe91abc04c397dd682d371126a7ceacf7c43ec  <=  ~I043258a364cd91821e9bb3e9c46441ac7d330c706e4b0b7e29c4b92f7c5ce562 + 1;
                end else begin
                    I5f1b294a0702ab37f94304ae67fe91abc04c397dd682d371126a7ceacf7c43ec  <= I043258a364cd91821e9bb3e9c46441ac7d330c706e4b0b7e29c4b92f7c5ce562 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[14] ) begin
                    I31c470f2adda0a23b85c3245646a168f2478bfdff11a434c1455be20db703c64  <=  ~I2f639b76b1afd86d9ba4d07d54f5b45df8cb99d7bc58cafd0c1a9a9001842260 + 1;
                end else begin
                    I31c470f2adda0a23b85c3245646a168f2478bfdff11a434c1455be20db703c64  <= I2f639b76b1afd86d9ba4d07d54f5b45df8cb99d7bc58cafd0c1a9a9001842260 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[5] ) begin
                    I152b3a1e710e5a39bac6338591c6597ee2a38fc25555f563beb7a1a967bf4e94  <=  ~I1dd0421d7e31a316541c339f8b4f1e3afbe37ce09254ed825c1b6086a0c0f3f2 + 1;
                end else begin
                    I152b3a1e710e5a39bac6338591c6597ee2a38fc25555f563beb7a1a967bf4e94  <= I1dd0421d7e31a316541c339f8b4f1e3afbe37ce09254ed825c1b6086a0c0f3f2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c != I4f9435bbcce379d6d591547481382ab188003b97877c0f32462ef9e33aa8bc1a[0] ) begin
                    I416c7ff28cd1d182ba2e08c3882c04d5073a014f7b9b41e56a3850cdc289ffb4  <=  ~I50ccddac87e61ba10dd9410a224c74ca88b521dfed962bf601c38ae78299384f + 1;
                end else begin
                    I416c7ff28cd1d182ba2e08c3882c04d5073a014f7b9b41e56a3850cdc289ffb4  <= I50ccddac87e61ba10dd9410a224c74ca88b521dfed962bf601c38ae78299384f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[12] ) begin
                    Ic195e053a186bcb0e653c0ddec75c57d1b3210c583162dd90978858c98fa53f2  <=  ~I5fd9960aaa562ff70e5d0e913dd4d88aac1b73a95c41ba903c0b7fc4dd4d93b2 + 1;
                end else begin
                    Ic195e053a186bcb0e653c0ddec75c57d1b3210c583162dd90978858c98fa53f2  <= I5fd9960aaa562ff70e5d0e913dd4d88aac1b73a95c41ba903c0b7fc4dd4d93b2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[14] ) begin
                    I8dcb7a5498da4a9d3e4a76923e84c88a30ec174503cd435864a066ff0ff464ba  <=  ~Icdff2336860758127c20c1d45d5723511fa42577417bf4f77d0c770abcbb175b + 1;
                end else begin
                    I8dcb7a5498da4a9d3e4a76923e84c88a30ec174503cd435864a066ff0ff464ba  <= Icdff2336860758127c20c1d45d5723511fa42577417bf4f77d0c770abcbb175b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[5] ) begin
                    I4f96b4022f127e7d965786f2cac8ee6afdbee96980608c876c6b699495f80b0f  <=  ~I9351e784be3825e94dcf67151cf38c9fddcf244bf5512db57dcc612882b449ce + 1;
                end else begin
                    I4f96b4022f127e7d965786f2cac8ee6afdbee96980608c876c6b699495f80b0f  <= I9351e784be3825e94dcf67151cf38c9fddcf244bf5512db57dcc612882b449ce ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636 != I9e497e3ee797c274b82ecca58218c47f9b663bcac21b1431b45c17d5e54e5a4a[0] ) begin
                    Ie44d1a587dcdbb709546c6c567988fb0a19c276a1df7aced4c09a029196dfd4b  <=  ~I23f7465a60acd0fb198e753834d30932ddab8939bb2df2172f54c7bdbe02e154 + 1;
                end else begin
                    Ie44d1a587dcdbb709546c6c567988fb0a19c276a1df7aced4c09a029196dfd4b  <= I23f7465a60acd0fb198e753834d30932ddab8939bb2df2172f54c7bdbe02e154 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[12] ) begin
                    I98e4b84e98742d38b206ac059ad123966ee63903c616b9c31b4ba9615edb9f40  <=  ~I40687a0e9fee803f38df7cf7dbc3d3107b859b4e80822bc59a157fdc606416b6 + 1;
                end else begin
                    I98e4b84e98742d38b206ac059ad123966ee63903c616b9c31b4ba9615edb9f40  <= I40687a0e9fee803f38df7cf7dbc3d3107b859b4e80822bc59a157fdc606416b6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[14] ) begin
                    I2c200a5ade27683d4afd55e06371f9880a7bb99259e2ccda5c368fe46bb385bd  <=  ~I807d8cd303e5c8c8379a9a2954804c606d897fc06412c924a89f3dc9e29909bd + 1;
                end else begin
                    I2c200a5ade27683d4afd55e06371f9880a7bb99259e2ccda5c368fe46bb385bd  <= I807d8cd303e5c8c8379a9a2954804c606d897fc06412c924a89f3dc9e29909bd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05 != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[5] ) begin
                    I105a7d84244a0d9143b9b2a3c64ea6964f7e1f43b7f8f5cb15d579885bbf746f  <=  ~I1244d935c6db7b5441533aab87f518ea215aa6f5903b071f2ee8cb3359b3bcb2 + 1;
                end else begin
                    I105a7d84244a0d9143b9b2a3c64ea6964f7e1f43b7f8f5cb15d579885bbf746f  <= I1244d935c6db7b5441533aab87f518ea215aa6f5903b071f2ee8cb3359b3bcb2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05 != Ib929181cef39d751d2726a054cd0478d309e58350ecd11d3363ecba8bd4cb7fa[0] ) begin
                    Ic2b8d811fd01f5cd88dd60bb1b89b33163b3cbeae48d04e2316f15500c6a1a40  <=  ~Ia7cdab2a88c99d9780bb267234b2cb87946009484d21f4419c50e7570438e645 + 1;
                end else begin
                    Ic2b8d811fd01f5cd88dd60bb1b89b33163b3cbeae48d04e2316f15500c6a1a40  <= Ia7cdab2a88c99d9780bb267234b2cb87946009484d21f4419c50e7570438e645 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[15] ) begin
                    I94024b61447a332a2c36a75bbf305f3fd80606bfbfcc4ee8c5783e3910e9840b  <=  ~Iacdbe6e2ae2cd5fa475cde0217452a14f05bc8d499b9ddeca568f6cd96ad6a2e + 1;
                end else begin
                    I94024b61447a332a2c36a75bbf305f3fd80606bfbfcc4ee8c5783e3910e9840b  <= Iacdbe6e2ae2cd5fa475cde0217452a14f05bc8d499b9ddeca568f6cd96ad6a2e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0 != Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[3] ) begin
                    If83264f9ff9f7b77429559aff8b14fce54040210c6ba3476b77824c28b95bea9  <=  ~I5aaf6ccf4cefc2732732ddd816c3eb7aea7146c6e7abf913a5193f6906fe9497 + 1;
                end else begin
                    If83264f9ff9f7b77429559aff8b14fce54040210c6ba3476b77824c28b95bea9  <= I5aaf6ccf4cefc2732732ddd816c3eb7aea7146c6e7abf913a5193f6906fe9497 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[12] ) begin
                    I7f9f83601cb61fece60f94c3120b43ca0c737ee36b8c67ccc917d3a428d8750a  <=  ~I96d8c1b67b028322f3d3e46d6306eac0333a8f3fe45073c08c5267157f73b71e + 1;
                end else begin
                    I7f9f83601cb61fece60f94c3120b43ca0c737ee36b8c67ccc917d3a428d8750a  <= I96d8c1b67b028322f3d3e46d6306eac0333a8f3fe45073c08c5267157f73b71e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0 != I64fa7f4fa09b7909840d8edb83f29f6a2379419e65b80f592b37d8ea00e59475[0] ) begin
                    I85ff9ab4f9a4a3301bb8fcdc7107202263af0c37f091445efb5fa163a6b47a51  <=  ~I600b1d1ff12460bfbaf32de67aff0e32087306628f0ba7db6736a81354309a41 + 1;
                end else begin
                    I85ff9ab4f9a4a3301bb8fcdc7107202263af0c37f091445efb5fa163a6b47a51  <= I600b1d1ff12460bfbaf32de67aff0e32087306628f0ba7db6736a81354309a41 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[15] ) begin
                    I92d28f6c97dab90de260df37f619e0a9000db48e278327a5c5d1528a34bb6dd2  <=  ~I225db641808b767d3f529e5ef2ac066e3abe953b8b434fd7bf4e02b57edc0f27 + 1;
                end else begin
                    I92d28f6c97dab90de260df37f619e0a9000db48e278327a5c5d1528a34bb6dd2  <= I225db641808b767d3f529e5ef2ac066e3abe953b8b434fd7bf4e02b57edc0f27 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f != I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[3] ) begin
                    I0f54db0f4bdec3ff62a8f1b5f4974982e3600a906dcfc79789fb9fac058c353c  <=  ~I1b7380bca98b56ba1a2c2ad5d78fdadc1112b208e8d98b84c8d950f3f12f1658 + 1;
                end else begin
                    I0f54db0f4bdec3ff62a8f1b5f4974982e3600a906dcfc79789fb9fac058c353c  <= I1b7380bca98b56ba1a2c2ad5d78fdadc1112b208e8d98b84c8d950f3f12f1658 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[12] ) begin
                    Icf4d3544466d430d71abf2513cfbc16b575af540d369d405ed831753f304673c  <=  ~I651492ce35fed9d77d5167dd211125ace0af8d55b8aff148e760d8919d53b6b8 + 1;
                end else begin
                    Icf4d3544466d430d71abf2513cfbc16b575af540d369d405ed831753f304673c  <= I651492ce35fed9d77d5167dd211125ace0af8d55b8aff148e760d8919d53b6b8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f != I35beac843abd6268c39acb691d3105a5c386f05461bca8c63b951ce1c2ed07bc[0] ) begin
                    I39ab1bf4bdde9805c5bc7695c4700975d5a6094c40e107b82477192005d9ce21  <=  ~Id732b4b9de3f715537d32d6eb6eca4f6f9fa6d634bc283ceaef531bdef605537 + 1;
                end else begin
                    I39ab1bf4bdde9805c5bc7695c4700975d5a6094c40e107b82477192005d9ce21  <= Id732b4b9de3f715537d32d6eb6eca4f6f9fa6d634bc283ceaef531bdef605537 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[15] ) begin
                    I4a5c4f290852b8c1baa90ae00400045825f13c24b546dc4a7848f91824185f7c  <=  ~I78c5859a565a68329d5f75effa2fbe77e16d86bbfcaf79d5480374f8bb87039c + 1;
                end else begin
                    I4a5c4f290852b8c1baa90ae00400045825f13c24b546dc4a7848f91824185f7c  <= I78c5859a565a68329d5f75effa2fbe77e16d86bbfcaf79d5480374f8bb87039c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474 != I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[3] ) begin
                    If45b8fca9a85788040c10a47569139b44384357512af96ee7bd8cd98d88f8f0f  <=  ~I411faecc88c5a9fcbc433d784eccf7024675c9b009564295eeb765079b8069c8 + 1;
                end else begin
                    If45b8fca9a85788040c10a47569139b44384357512af96ee7bd8cd98d88f8f0f  <= I411faecc88c5a9fcbc433d784eccf7024675c9b009564295eeb765079b8069c8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[12] ) begin
                    I329448311438699d3d590bba6ab4bfc9cead805f96015b77617f42d957bde7d5  <=  ~Ic429f74c6e97fa699700391c81e8a8ac449270476ebded49a8bcf8161a19260e + 1;
                end else begin
                    I329448311438699d3d590bba6ab4bfc9cead805f96015b77617f42d957bde7d5  <= Ic429f74c6e97fa699700391c81e8a8ac449270476ebded49a8bcf8161a19260e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474 != I9d8fbde44d35c50f5f24ceae6f2e16ca2f280573caeb8a3021b6f69dec3d04b4[0] ) begin
                    I602591ae56f1a42c64e50378841e065e79aee138622a0a571effe20cb48645a3  <=  ~I6efa3ca79fc64053e7e2744a4248a5c0df63ef15c66542967b53b2fcefe0d286 + 1;
                end else begin
                    I602591ae56f1a42c64e50378841e065e79aee138622a0a571effe20cb48645a3  <= I6efa3ca79fc64053e7e2744a4248a5c0df63ef15c66542967b53b2fcefe0d286 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[15] ) begin
                    I9fa9c98579041b6735eb78f7b3727824dd61991c6a6d91a158c6ac65cb20b05d  <=  ~I00827962c46c637f5d74d450ff4eae848b4cb15add5bf1f607708b76c8551c21 + 1;
                end else begin
                    I9fa9c98579041b6735eb78f7b3727824dd61991c6a6d91a158c6ac65cb20b05d  <= I00827962c46c637f5d74d450ff4eae848b4cb15add5bf1f607708b76c8551c21 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987 != Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[3] ) begin
                    Id6b81456b5d3050b4e1fe80ccc8f992cf56eb0f08a1d29ec1e7cabe1baeb0872  <=  ~I6cb1364420f9bdd072770a684de242f89990e3f144f160c2f5311bb00fe4daa0 + 1;
                end else begin
                    Id6b81456b5d3050b4e1fe80ccc8f992cf56eb0f08a1d29ec1e7cabe1baeb0872  <= I6cb1364420f9bdd072770a684de242f89990e3f144f160c2f5311bb00fe4daa0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[12] ) begin
                    Icb61d0767612534695d9de0380a1febbda612604f373afa55f0339c7a679e99e  <=  ~I41bc9fc093e9f311e6376edb8aa0640709fb3bd420ff8a7cb2092844fbe0e121 + 1;
                end else begin
                    Icb61d0767612534695d9de0380a1febbda612604f373afa55f0339c7a679e99e  <= I41bc9fc093e9f311e6376edb8aa0640709fb3bd420ff8a7cb2092844fbe0e121 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987 != I507d851a78a765c18af6d529292384fb4cbb06cfec0e22d516adc79b8ea13c7f[0] ) begin
                    If37e9ed3af8a31c989dc6ad554207cd464c591b630ca1e5cf56b2eca57a18d8c  <=  ~I84519b5d45c05d737fb27ebd20ddbddfdaf7a22125df9eea17400856eed27992 + 1;
                end else begin
                    If37e9ed3af8a31c989dc6ad554207cd464c591b630ca1e5cf56b2eca57a18d8c  <= I84519b5d45c05d737fb27ebd20ddbddfdaf7a22125df9eea17400856eed27992 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[13] ) begin
                    I81aa911c9f6f4bd88314aa3c5310efef6c40219ca93521bbea3c1afcea7bb48f  <=  ~I3af2de27ab7a899c5e55f150a53b7ef65e88309f4280269afb3eda2b1b408d05 + 1;
                end else begin
                    I81aa911c9f6f4bd88314aa3c5310efef6c40219ca93521bbea3c1afcea7bb48f  <= I3af2de27ab7a899c5e55f150a53b7ef65e88309f4280269afb3eda2b1b408d05 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e != I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[5] ) begin
                    I2e557a901de23b8442e8002b3560bbf9cb8592b7bfb7a6e2f8aad12843a5a041  <=  ~I988d8e969e2a2ecac68a36a5f4eb0d6cb2c325e4be24c4716625070057ab9538 + 1;
                end else begin
                    I2e557a901de23b8442e8002b3560bbf9cb8592b7bfb7a6e2f8aad12843a5a041  <= I988d8e969e2a2ecac68a36a5f4eb0d6cb2c325e4be24c4716625070057ab9538 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[6] ) begin
                    I0d25b3618b50ff21e3f301fe44087368e38fd6b37b6f6fab004824aa9df51f0b  <=  ~I63ec7fce46bb02bd1662b19d58025abb479c4b57a0e4fd0642404ddf7f607077 + 1;
                end else begin
                    I0d25b3618b50ff21e3f301fe44087368e38fd6b37b6f6fab004824aa9df51f0b  <= I63ec7fce46bb02bd1662b19d58025abb479c4b57a0e4fd0642404ddf7f607077 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e != I80fb8d450dd144ffade989cc2cec363cf6bbcdc267f5372163fde38313387499[0] ) begin
                    I80099c7b01770cc5f7edb3a3551d8edfe9dccbcd2a12daf8ebbafdfccd141bd4  <=  ~I086c1b2b7346139212d810647d98824eff245a9e24fa84006583fd56f1e76926 + 1;
                end else begin
                    I80099c7b01770cc5f7edb3a3551d8edfe9dccbcd2a12daf8ebbafdfccd141bd4  <= I086c1b2b7346139212d810647d98824eff245a9e24fa84006583fd56f1e76926 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[13] ) begin
                    Ic859d34db6baa83e73a8627c251c877e93f15653973d0634c42a8ffc9f628bae  <=  ~I401154446147692cdd273c1d6dbe5a225e466799d41dd00f9477c586add460a4 + 1;
                end else begin
                    Ic859d34db6baa83e73a8627c251c877e93f15653973d0634c42a8ffc9f628bae  <= I401154446147692cdd273c1d6dbe5a225e466799d41dd00f9477c586add460a4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229 != I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[5] ) begin
                    I823e337e6437e5ba36ecaf0b1ac6b7a4e74cd2ed7019dd5447355626a8877d89  <=  ~If832820141ab4f3c34efb429966b47ce584cf58fd34d38a7ecd976235613c541 + 1;
                end else begin
                    I823e337e6437e5ba36ecaf0b1ac6b7a4e74cd2ed7019dd5447355626a8877d89  <= If832820141ab4f3c34efb429966b47ce584cf58fd34d38a7ecd976235613c541 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[6] ) begin
                    I068f00aade8307d2a2e2ddb37d7429a04c2f6786232134a041e62733cadb03ac  <=  ~If13409b9d8c65fe2127031b0e4f953f55c8a66c06811c6a5d261372aa2986511 + 1;
                end else begin
                    I068f00aade8307d2a2e2ddb37d7429a04c2f6786232134a041e62733cadb03ac  <= If13409b9d8c65fe2127031b0e4f953f55c8a66c06811c6a5d261372aa2986511 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229 != I7844074cddcce1b95a010729a9e4ce2bfc4f7e1962b84af0e0a3cbb2c2c08206[0] ) begin
                    Ie479ccbabaa8a00009152557e4de08bd240fd28f1b131c674dafbcc2505711f7  <=  ~Id2bc1d218fffb230a1505feb20cfb5229db9f3e2b0c7bb005bc8c59403fa35ad + 1;
                end else begin
                    Ie479ccbabaa8a00009152557e4de08bd240fd28f1b131c674dafbcc2505711f7  <= Id2bc1d218fffb230a1505feb20cfb5229db9f3e2b0c7bb005bc8c59403fa35ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[13] ) begin
                    I40d7eae63827c6efe2ac480c8eb9f8a8f77bbfa845caae02d137397c9da822a9  <=  ~Ia1846f3088723131b0fc158b2d942749466887bf940e29340846070ac9d5090b + 1;
                end else begin
                    I40d7eae63827c6efe2ac480c8eb9f8a8f77bbfa845caae02d137397c9da822a9  <= Ia1846f3088723131b0fc158b2d942749466887bf940e29340846070ac9d5090b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96 != I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[5] ) begin
                    I259a9b6041f341013e6ea0706c4e9ef9a77148bc003b3f0cf9593ebd915b30c1  <=  ~I5d5edfd68cef65681c36f4bcd770ec84a721eb515bc1d0fb7603ee0f5a63fabb + 1;
                end else begin
                    I259a9b6041f341013e6ea0706c4e9ef9a77148bc003b3f0cf9593ebd915b30c1  <= I5d5edfd68cef65681c36f4bcd770ec84a721eb515bc1d0fb7603ee0f5a63fabb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[6] ) begin
                    I5b4c4554a78c551dd34a93ceb225237a2d2540a0e05311c4595bdaa5a4cb14ea  <=  ~I9efcedaa1cc036ad8613f9ba801ca4ff4afcd709f5e4aaadbcdcd130d1263fc8 + 1;
                end else begin
                    I5b4c4554a78c551dd34a93ceb225237a2d2540a0e05311c4595bdaa5a4cb14ea  <= I9efcedaa1cc036ad8613f9ba801ca4ff4afcd709f5e4aaadbcdcd130d1263fc8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96 != I88be0c0499713ce396832a79853e9918ecdfed2519fba6fd7c0bae51450478e7[0] ) begin
                    I6364406b04427fe3a4cecbed48e12a67cb08dc632b2914b0fe52fab0ca541c0d  <=  ~I26dc2d992b646fe215751740a4406ce2a30e06fa2251f0382248aed7a08071be + 1;
                end else begin
                    I6364406b04427fe3a4cecbed48e12a67cb08dc632b2914b0fe52fab0ca541c0d  <= I26dc2d992b646fe215751740a4406ce2a30e06fa2251f0382248aed7a08071be ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[13] ) begin
                    I7c6d90cd79e1b85ce9a5452570cfeec8faf9ce3e6bc886f66495ec2a66fc8c7e  <=  ~If25d531f7d1101b94167fde8f48549338e9b003202bc68bcb851f94fccb01007 + 1;
                end else begin
                    I7c6d90cd79e1b85ce9a5452570cfeec8faf9ce3e6bc886f66495ec2a66fc8c7e  <= If25d531f7d1101b94167fde8f48549338e9b003202bc68bcb851f94fccb01007 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5 != I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[5] ) begin
                    I3225ba7b6d0e0c7a94dfbc8e074ade02b79a66f6aaf97580a451c2d1781a625c  <=  ~I3e49103842dcd70cc7795bfb356ef7d178c1e87d94c08cbef0794b0956dff7b9 + 1;
                end else begin
                    I3225ba7b6d0e0c7a94dfbc8e074ade02b79a66f6aaf97580a451c2d1781a625c  <= I3e49103842dcd70cc7795bfb356ef7d178c1e87d94c08cbef0794b0956dff7b9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[6] ) begin
                    Ice3b06f04279add8283c8173340c2bfd4b4801d85610179943f070aef508a893  <=  ~I84b78cf1294735491099a4ece1a26f5a1bed53ffd09724d3383bc63756866721 + 1;
                end else begin
                    Ice3b06f04279add8283c8173340c2bfd4b4801d85610179943f070aef508a893  <= I84b78cf1294735491099a4ece1a26f5a1bed53ffd09724d3383bc63756866721 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5 != Ib585733bf4c3eb59a772866965420fc7397b01272410cdb701f289daf9549fc9[0] ) begin
                    I610dd39f1d44d84764b0acd6b3fb1219fb6b6d6ca92e1b226ca76a389bf6c937  <=  ~I964fe2ac03da8dd1965fd87a79f3fb2adf8e1607b64404233c3a09867227531e + 1;
                end else begin
                    I610dd39f1d44d84764b0acd6b3fb1219fb6b6d6ca92e1b226ca76a389bf6c937  <= I964fe2ac03da8dd1965fd87a79f3fb2adf8e1607b64404233c3a09867227531e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icf75206b75ca695f888c3d924d2f1822806f452b5d29a0d6084dbd1c00a15790 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[16] ) begin
                    Ibcddbd4e851466c5ff49f13244c2478ab6c089e6d8ad294cdfbdc8451ac6a895  <=  ~I58df6e4342bc054f0177b7c91a68a1afdac21b2d1d52434ef5d8272b92fef6d9 + 1;
                end else begin
                    Ibcddbd4e851466c5ff49f13244c2478ab6c089e6d8ad294cdfbdc8451ac6a895  <= I58df6e4342bc054f0177b7c91a68a1afdac21b2d1d52434ef5d8272b92fef6d9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icf75206b75ca695f888c3d924d2f1822806f452b5d29a0d6084dbd1c00a15790 != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[2] ) begin
                    I492e47d35231729b266a9f31aba61a3ac2c93a9786a20f6a152d342cd1d0b911  <=  ~Iac61de7786d6ba1a40fc62f7d70b3cb366469c6674ebc4ecdaa21346903a58ff + 1;
                end else begin
                    I492e47d35231729b266a9f31aba61a3ac2c93a9786a20f6a152d342cd1d0b911  <= Iac61de7786d6ba1a40fc62f7d70b3cb366469c6674ebc4ecdaa21346903a58ff ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icf75206b75ca695f888c3d924d2f1822806f452b5d29a0d6084dbd1c00a15790 != Ida673298c761bab46fb26d4e73caa99f5b3ade7f924d99fcedae4e47c70b5b67[0] ) begin
                    Ib9f9384ac4ec4bad29fbb4ce683ffda7dcab311135f02b6336e6209f5742fddd  <=  ~I3c94620659b19b26861b2f4dc674bd9b9ddd8a378f11b67d27bc0f7639e0842c + 1;
                end else begin
                    Ib9f9384ac4ec4bad29fbb4ce683ffda7dcab311135f02b6336e6209f5742fddd  <= I3c94620659b19b26861b2f4dc674bd9b9ddd8a378f11b67d27bc0f7639e0842c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4a1896458491f2613d2c7274b81fbb7a9d405272b871b504455b388a3695acae != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[16] ) begin
                    Ib053c04dd4e330e6784846706317bb6c8b12f9b36a57ee12807bff7de8ba7f0c  <=  ~I4aeb03994ab1826b4bc249e1cdcbda394b864bcec0ca3bd6a0897fafa6d280f6 + 1;
                end else begin
                    Ib053c04dd4e330e6784846706317bb6c8b12f9b36a57ee12807bff7de8ba7f0c  <= I4aeb03994ab1826b4bc249e1cdcbda394b864bcec0ca3bd6a0897fafa6d280f6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4a1896458491f2613d2c7274b81fbb7a9d405272b871b504455b388a3695acae != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[2] ) begin
                    I18777be7a1745485d18289e0b4a6e43e8a2e6758be0967b8cea04a3b0faf973f  <=  ~I4d24219bb14476929c0d4b4bbef3ecee057061ad24af5601a8de67871680ee10 + 1;
                end else begin
                    I18777be7a1745485d18289e0b4a6e43e8a2e6758be0967b8cea04a3b0faf973f  <= I4d24219bb14476929c0d4b4bbef3ecee057061ad24af5601a8de67871680ee10 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4a1896458491f2613d2c7274b81fbb7a9d405272b871b504455b388a3695acae != I60bb81cc7cd9a6212f7b4261a21655accd6cd09e7aaf5f78f7f1f4dec0e8489b[0] ) begin
                    I60980f76d468775bcc8a7052681fbb6ef4b2243e5e30e5365cda6cf598bd0bde  <=  ~I6729f7458757e512a921fff6abb9aa05fb498db59115c3b041bad959c15fad3f + 1;
                end else begin
                    I60980f76d468775bcc8a7052681fbb6ef4b2243e5e30e5365cda6cf598bd0bde  <= I6729f7458757e512a921fff6abb9aa05fb498db59115c3b041bad959c15fad3f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If122210c8dc39e7ab2fecb27dac5c167b39ccd9e8e4cd076b2b3b92632357248 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[16] ) begin
                    I9af65d3592633577409561b2069e30c73196d1a4798cb92f4d2f14db8771895c  <=  ~I543c9825f790b1e9264e3f6b5e66e64c773dd0866bda372b2eda0201910105e9 + 1;
                end else begin
                    I9af65d3592633577409561b2069e30c73196d1a4798cb92f4d2f14db8771895c  <= I543c9825f790b1e9264e3f6b5e66e64c773dd0866bda372b2eda0201910105e9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If122210c8dc39e7ab2fecb27dac5c167b39ccd9e8e4cd076b2b3b92632357248 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[2] ) begin
                    I9b13cfb3566db96edc7c018b88f158faa57e4db029e3982290989c6fc08163b2  <=  ~I8097cf47b760092e87e117165f17e1f66afbaa3ee78160fd0e2a597f613883ee + 1;
                end else begin
                    I9b13cfb3566db96edc7c018b88f158faa57e4db029e3982290989c6fc08163b2  <= I8097cf47b760092e87e117165f17e1f66afbaa3ee78160fd0e2a597f613883ee ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If122210c8dc39e7ab2fecb27dac5c167b39ccd9e8e4cd076b2b3b92632357248 != I85d3c885ce504524ab43daed7bbcb599cd7e5d6d3635cf46e278345134e97e22[0] ) begin
                    I892a754f0322d92126d4731e8066760a24897f93e2afb858ee1393604d2cbb26  <=  ~I4eb210e31e4ad434958f477b79dcf5b2694caf5c18f801a8d3b3b612eb0812af + 1;
                end else begin
                    I892a754f0322d92126d4731e8066760a24897f93e2afb858ee1393604d2cbb26  <= I4eb210e31e4ad434958f477b79dcf5b2694caf5c18f801a8d3b3b612eb0812af ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iea6e52ee89805cbf2f2a65f695323d8dd7669c23df341897eff049fbcbd1db98 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[16] ) begin
                    I9fc6fbd6f2f888b9750fa59a966971aa6ba6fe4eee8c8f3ed4c3ea60141a7d23  <=  ~I40b6ad89db699e7f672e55f672bfc979d85a462330e526aefd63b9724ff7de89 + 1;
                end else begin
                    I9fc6fbd6f2f888b9750fa59a966971aa6ba6fe4eee8c8f3ed4c3ea60141a7d23  <= I40b6ad89db699e7f672e55f672bfc979d85a462330e526aefd63b9724ff7de89 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iea6e52ee89805cbf2f2a65f695323d8dd7669c23df341897eff049fbcbd1db98 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[2] ) begin
                    I3baaba73f51f47e6a3f2310f692de9f7b9a871c65605e14d204d6965153ff4f0  <=  ~I014e96c75acbbe2bf38e1c89b52e1a331eb3d31b984a67946eef2a5223b87855 + 1;
                end else begin
                    I3baaba73f51f47e6a3f2310f692de9f7b9a871c65605e14d204d6965153ff4f0  <= I014e96c75acbbe2bf38e1c89b52e1a331eb3d31b984a67946eef2a5223b87855 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Iea6e52ee89805cbf2f2a65f695323d8dd7669c23df341897eff049fbcbd1db98 != Iaa08a49e0ca4f92f38c7f4d115ae1b275e45c42dfa6fd4b6a2ff40536b7f5f15[0] ) begin
                    Ib0f8816eafd3b950f67cfbdb6a44c59ab7c0918979817a4a998d8305da847e72  <=  ~Ia3588e449670d7edbf99e52ccf0d7c8462b51e3d24ec5f0f7293290d47154f72 + 1;
                end else begin
                    Ib0f8816eafd3b950f67cfbdb6a44c59ab7c0918979817a4a998d8305da847e72  <= Ia3588e449670d7edbf99e52ccf0d7c8462b51e3d24ec5f0f7293290d47154f72 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[14] ) begin
                    I57d80f41498f8d7b91410dc02e646a45a3f05d45e9b5871ae95d6432ecd2af56  <=  ~I6b3108db71d5eaffc5606fb88fe909a0462a77232258fd85cb6792954ad28c0b + 1;
                end else begin
                    I57d80f41498f8d7b91410dc02e646a45a3f05d45e9b5871ae95d6432ecd2af56  <= I6b3108db71d5eaffc5606fb88fe909a0462a77232258fd85cb6792954ad28c0b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa != I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[4] ) begin
                    Ib924c4eaf872874debc3b6ee65921f0381331e1421cbfc3bd17e8caf273049cb  <=  ~I55a1e3e076ea304ccd72b18524bfa076977a0f791806719d752ed020cb6c3e37 + 1;
                end else begin
                    Ib924c4eaf872874debc3b6ee65921f0381331e1421cbfc3bd17e8caf273049cb  <= I55a1e3e076ea304ccd72b18524bfa076977a0f791806719d752ed020cb6c3e37 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[6] ) begin
                    Ib1310cd21337a1faa061ffd12a2670171f582e03471ab315b90de9f8fc30959a  <=  ~I318f0ddae7fd42b63d856ad6923268574eb4f8f71cbdddcaa420e917a1d7ea51 + 1;
                end else begin
                    Ib1310cd21337a1faa061ffd12a2670171f582e03471ab315b90de9f8fc30959a  <= I318f0ddae7fd42b63d856ad6923268574eb4f8f71cbdddcaa420e917a1d7ea51 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa != I197b3231cb1da107c5001075809e9fa75e4089871d473490981a8b44d3ff5e4c[0] ) begin
                    I04b55f2c45002f1f1f7a6176773a22730dcfea14662f0badb102ddb60b84cf9d  <=  ~Iee19c6e30e6fb9258878db36251e2e15a071b41364b59473c9de2c0f0b8c9ce8 + 1;
                end else begin
                    I04b55f2c45002f1f1f7a6176773a22730dcfea14662f0badb102ddb60b84cf9d  <= Iee19c6e30e6fb9258878db36251e2e15a071b41364b59473c9de2c0f0b8c9ce8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[14] ) begin
                    I97f674eaee005fc7a54ccb648f5a0a67cec041e895d62eacbcc9a37068b912a7  <=  ~I4a9362c36b4a88ee5422688ee5550c97e8fe10b4cc23b6538ee81bfeef1472a9 + 1;
                end else begin
                    I97f674eaee005fc7a54ccb648f5a0a67cec041e895d62eacbcc9a37068b912a7  <= I4a9362c36b4a88ee5422688ee5550c97e8fe10b4cc23b6538ee81bfeef1472a9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2 != I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[4] ) begin
                    I730fa6d01ade8f1439b29b955c5cff62700a90e523a4f4208ca2f9978e59afcd  <=  ~I9dda3335af58c2daa92010ef90e217e0842b7740a65ce2a029ebde5b65e9fc86 + 1;
                end else begin
                    I730fa6d01ade8f1439b29b955c5cff62700a90e523a4f4208ca2f9978e59afcd  <= I9dda3335af58c2daa92010ef90e217e0842b7740a65ce2a029ebde5b65e9fc86 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[6] ) begin
                    I2862bdd9be64c24d98e80e8b662a7c97c70943bab3d49cc8d39443abcd5c2c3c  <=  ~I996cd6ee71fdd8f4b109acfd52bf495951439b9e49b87a6db4565bebbc7d1e1d + 1;
                end else begin
                    I2862bdd9be64c24d98e80e8b662a7c97c70943bab3d49cc8d39443abcd5c2c3c  <= I996cd6ee71fdd8f4b109acfd52bf495951439b9e49b87a6db4565bebbc7d1e1d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2 != I384c04b75344f97c691f70965d7e08266ab9cd8862e04ba73b502a0f36ac5ea7[0] ) begin
                    I5edc072d158ac583bd1cdb2449086d4f0b17e36d724f4cfde79820788ce57f31  <=  ~I705cf789e535bcc9523034b7f4743daa8f66f1dfa3d15c77b87e9f1845563690 + 1;
                end else begin
                    I5edc072d158ac583bd1cdb2449086d4f0b17e36d724f4cfde79820788ce57f31  <= I705cf789e535bcc9523034b7f4743daa8f66f1dfa3d15c77b87e9f1845563690 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[14] ) begin
                    Ibeb23788ce301c724494a2852312b38344c27416a5604c0145fa330ccd1f290d  <=  ~I4345f323dbf4da279580851ea1d0b7a2e5109f518ca914c88b6ac91e9ce8625c + 1;
                end else begin
                    Ibeb23788ce301c724494a2852312b38344c27416a5604c0145fa330ccd1f290d  <= I4345f323dbf4da279580851ea1d0b7a2e5109f518ca914c88b6ac91e9ce8625c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236 != Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[4] ) begin
                    I425913b12fc3c865d95f1caead00d8c49de08765b634aa444243f4a03a53d0df  <=  ~I8a484469fd2c86173f27a68b9ae6c15c3813761e5dc1035c2f9fe04b24a6d73d + 1;
                end else begin
                    I425913b12fc3c865d95f1caead00d8c49de08765b634aa444243f4a03a53d0df  <= I8a484469fd2c86173f27a68b9ae6c15c3813761e5dc1035c2f9fe04b24a6d73d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[6] ) begin
                    I33d759e40b55a0d83119f5c19cf87e6e3181c7e3eed94eec60fb52f9c376addd  <=  ~Ic6518d2e4de9b3feb98b24f5ff4fd43edb699fad33847f2e67ff731825f15177 + 1;
                end else begin
                    I33d759e40b55a0d83119f5c19cf87e6e3181c7e3eed94eec60fb52f9c376addd  <= Ic6518d2e4de9b3feb98b24f5ff4fd43edb699fad33847f2e67ff731825f15177 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236 != Ibf95afb3941a2272d76cd7256d0789f11fb35a3020c3ccca5b099d335d4a2330[0] ) begin
                    Ieb128919ed64e331affb6adba798c267e8c3ec924a7ef58f50b1bc0b29702c23  <=  ~Ie147f013af77ffb57ecdf0bac185fd60648505960bec48f3f18094b1b7e319ca + 1;
                end else begin
                    Ieb128919ed64e331affb6adba798c267e8c3ec924a7ef58f50b1bc0b29702c23  <= Ie147f013af77ffb57ecdf0bac185fd60648505960bec48f3f18094b1b7e319ca ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[14] ) begin
                    I30a9d5330fac5c3ec7b63cfab0edcef0eda61dddb23d2aabf733b9982c12b4ad  <=  ~I0a51859ca31f0b470011ae2b3bcbd11fd2c79f03c854103f016b54af79028ba1 + 1;
                end else begin
                    I30a9d5330fac5c3ec7b63cfab0edcef0eda61dddb23d2aabf733b9982c12b4ad  <= I0a51859ca31f0b470011ae2b3bcbd11fd2c79f03c854103f016b54af79028ba1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915 != Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[4] ) begin
                    I2abc1178fa35959d8eb41342a7d7289e29054439c7bc06adc61f3a1d2e55bd6f  <=  ~I1f5d36144836b1c2e41164adaa02934f77b47f317c3f6e7452ea483c756b4ba3 + 1;
                end else begin
                    I2abc1178fa35959d8eb41342a7d7289e29054439c7bc06adc61f3a1d2e55bd6f  <= I1f5d36144836b1c2e41164adaa02934f77b47f317c3f6e7452ea483c756b4ba3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[6] ) begin
                    Ie2abebb2c2604e435cea102275e0726254ad91df1973aece477e1e5315f82d0b  <=  ~Ie1c46630d4cd6028c341687f4df0c2220054b63f8263fab4a11d3ad89f6518cd + 1;
                end else begin
                    Ie2abebb2c2604e435cea102275e0726254ad91df1973aece477e1e5315f82d0b  <= Ie1c46630d4cd6028c341687f4df0c2220054b63f8263fab4a11d3ad89f6518cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915 != I885622bb1c7371f4afa3e9966f870d2bf7750c2d2280a2a993a5bd9854187994[0] ) begin
                    I90cc372cc2f3b23eaaf2cb32da95ee715af64ca2eaee77195d9813647d2a0d08  <=  ~Iedab2e8aa599a943abe7d0d1dabb0f7a5a7d4b97f36e982d5f548a4acccfe2c2 + 1;
                end else begin
                    I90cc372cc2f3b23eaaf2cb32da95ee715af64ca2eaee77195d9813647d2a0d08  <= Iedab2e8aa599a943abe7d0d1dabb0f7a5a7d4b97f36e982d5f548a4acccfe2c2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[17] ) begin
                    I50ff347e89fb452beb071f112e4a51e074cb3d66bd903552db23c17670286e7b  <=  ~Ic7ecf5c9528425bf54c120398b0e5f75dcd4acd18b3088fd8a16fe8207a592bf + 1;
                end else begin
                    I50ff347e89fb452beb071f112e4a51e074cb3d66bd903552db23c17670286e7b  <= Ic7ecf5c9528425bf54c120398b0e5f75dcd4acd18b3088fd8a16fe8207a592bf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204 != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[3] ) begin
                    I2624a2d841eeb09774127e5d709364f803826266b46f0fc3122fcdcf0aa129e6  <=  ~I355cc82d012dbfaa00529a9197d4fe0b654fc609360a0775d398ae0b3e95f2cd + 1;
                end else begin
                    I2624a2d841eeb09774127e5d709364f803826266b46f0fc3122fcdcf0aa129e6  <= I355cc82d012dbfaa00529a9197d4fe0b654fc609360a0775d398ae0b3e95f2cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204 != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[6] ) begin
                    Ic0a892c18037ef674c8d94cdfc94cfca47d977ca2da9e678303255b96575f022  <=  ~Ic0c2a03a257040df478653886a3a2400777322b4d4333c0da94211227433697f + 1;
                end else begin
                    Ic0a892c18037ef674c8d94cdfc94cfca47d977ca2da9e678303255b96575f022  <= Ic0c2a03a257040df478653886a3a2400777322b4d4333c0da94211227433697f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204 != I719a3e78d6a298f7db920bf7e355f6fca2c46135abb8ccd1cc3ea470912d05c1[0] ) begin
                    Idaf65411d995039ea730b6ee4b5ae727325da17dc79c8664270d60f063828453  <=  ~Ic09079bc0fb0e140e7285e2e5af8caa802db98a774db8ce0bc5158e08becb4c1 + 1;
                end else begin
                    Idaf65411d995039ea730b6ee4b5ae727325da17dc79c8664270d60f063828453  <= Ic09079bc0fb0e140e7285e2e5af8caa802db98a774db8ce0bc5158e08becb4c1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[17] ) begin
                    I0f71479f871309f1717e7a1a2372ebfff4623c315cc31914588df3896740a074  <=  ~Ia7d33f990e505c818a46c2a54c13bd6680e3a34847708d89ee6f38999242e0b4 + 1;
                end else begin
                    I0f71479f871309f1717e7a1a2372ebfff4623c315cc31914588df3896740a074  <= Ia7d33f990e505c818a46c2a54c13bd6680e3a34847708d89ee6f38999242e0b4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[3] ) begin
                    I1c30d2957a73fc51bb7044b869e28e0a8f6e0378a6098ee5e244efb43ab6a690  <=  ~I0c87558b4bcfed105da91186dbea82b0f8d38c2473b578fb874ebd3e844edf51 + 1;
                end else begin
                    I1c30d2957a73fc51bb7044b869e28e0a8f6e0378a6098ee5e244efb43ab6a690  <= I0c87558b4bcfed105da91186dbea82b0f8d38c2473b578fb874ebd3e844edf51 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460 != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[6] ) begin
                    Ie1447c9e1eb4ed110e6b0353bc5dd2cd14ec645355c3cf897df6f6c5808475ad  <=  ~I5a7f5ab868cc2f4e823808a238df41f5e29c98d896557abab5eb1b5ac4231eeb + 1;
                end else begin
                    Ie1447c9e1eb4ed110e6b0353bc5dd2cd14ec645355c3cf897df6f6c5808475ad  <= I5a7f5ab868cc2f4e823808a238df41f5e29c98d896557abab5eb1b5ac4231eeb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460 != I1729b841d155c32b617727459f01aa9a9a6af56de5f464e20e900e3a4da30dba[0] ) begin
                    I977557441002c273f9b9b8748ffa9edceadb342e028ceb581c3bbce9af103a74  <=  ~If3574e7d834ff9a2b7247d3262dcd4265a5aa04a73495afc4e8098f7da4cd0ce + 1;
                end else begin
                    I977557441002c273f9b9b8748ffa9edceadb342e028ceb581c3bbce9af103a74  <= If3574e7d834ff9a2b7247d3262dcd4265a5aa04a73495afc4e8098f7da4cd0ce ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[17] ) begin
                    Ie2261f6d4e2c2ce04997cd365593486e02a7d85106b9c3b568ccdfcda7a9c352  <=  ~I5187aa2268c0345b27861b3f411a57adfe94104cd1a48c7573407a0f79e345d6 + 1;
                end else begin
                    Ie2261f6d4e2c2ce04997cd365593486e02a7d85106b9c3b568ccdfcda7a9c352  <= I5187aa2268c0345b27861b3f411a57adfe94104cd1a48c7573407a0f79e345d6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[3] ) begin
                    I8a1ba53134dcd1141a6f03dbed0f18ff7be9728dd9a6d6b138ff266c5307ba24  <=  ~If54927516082a9fec583e3cdeaf09539203d2f351771381d6c29c7961dc6f98a + 1;
                end else begin
                    I8a1ba53134dcd1141a6f03dbed0f18ff7be9728dd9a6d6b138ff266c5307ba24  <= If54927516082a9fec583e3cdeaf09539203d2f351771381d6c29c7961dc6f98a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3 != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[6] ) begin
                    I4a98524c02346f4b9468666ffaa9d996b9b868a5a8730264d798d7a66b7454bc  <=  ~I8e63aa98e26c7163ac7e004f9b363177513859fd81ce1d6be355e187166ee55a + 1;
                end else begin
                    I4a98524c02346f4b9468666ffaa9d996b9b868a5a8730264d798d7a66b7454bc  <= I8e63aa98e26c7163ac7e004f9b363177513859fd81ce1d6be355e187166ee55a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3 != I96affe6d042e09b07278ae45744977fd3719a31fa5d578adaa2b3a66b2c3ebd0[0] ) begin
                    Icc10ac19a64065f5923ecef4f1353f13c7796c23f2555f8ae6566eb538d77677  <=  ~I6e3f1705d8ba2b2cbd6b7749bf249716ede50edeca032e277396a885c69399ef + 1;
                end else begin
                    Icc10ac19a64065f5923ecef4f1353f13c7796c23f2555f8ae6566eb538d77677  <= I6e3f1705d8ba2b2cbd6b7749bf249716ede50edeca032e277396a885c69399ef ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[17] ) begin
                    I8c133563a8b5e359a6a45a7f3b4e939fc84766f9fa09634d18e5d2101d0c0645  <=  ~Idc29a95902384ae5ae3858cc3583cfc2fb39d4634b67c3c9858b9b6b9468fc87 + 1;
                end else begin
                    I8c133563a8b5e359a6a45a7f3b4e939fc84766f9fa09634d18e5d2101d0c0645  <= Idc29a95902384ae5ae3858cc3583cfc2fb39d4634b67c3c9858b9b6b9468fc87 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[3] ) begin
                    I82d316ed1475017844ea73f32085b755d17c9fdafd8191df2e363496e1950869  <=  ~I3ee26418f368f28b1dbc386529fe4d0034170fceeaa1cf5f4edd2132db250ab6 + 1;
                end else begin
                    I82d316ed1475017844ea73f32085b755d17c9fdafd8191df2e363496e1950869  <= I3ee26418f368f28b1dbc386529fe4d0034170fceeaa1cf5f4edd2132db250ab6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253 != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[6] ) begin
                    Iac7a05e270cb898af4ba32c16445d0dbdffdafdcc5fae209f09367abcff9d6b7  <=  ~I82393d9631be548b7d2f25eff102ffad6a2a1b7a683c82d8046dfd07b66e26a3 + 1;
                end else begin
                    Iac7a05e270cb898af4ba32c16445d0dbdffdafdcc5fae209f09367abcff9d6b7  <= I82393d9631be548b7d2f25eff102ffad6a2a1b7a683c82d8046dfd07b66e26a3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253 != I12e1e01b28d2d443785fac1d0314b477b221b17b715f1153c5379a85b4b5e3aa[0] ) begin
                    I725c369a5013eeb6b581209bc8a921fccfcf1754137191e26757abdb72ced94b  <=  ~I61291a36d4d546d1cb7c79a8a8c9ccbb4da2bf3fe853e05a56296804d5fde212 + 1;
                end else begin
                    I725c369a5013eeb6b581209bc8a921fccfcf1754137191e26757abdb72ced94b  <= I61291a36d4d546d1cb7c79a8a8c9ccbb4da2bf3fe853e05a56296804d5fde212 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idc77bba153be5873f87a4cf88c6ddc6a89bf8aa3ffcd29702126b01053f012f2 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[15] ) begin
                    I7628fd0a5ee3ec547c1b4798a4d76de651807424cd18f0b3b8a3bea849e6fe0d  <=  ~I454cdecfffd5c06b833e81e8990b07a9b326eec23f31a7b6589b969f610d8ed6 + 1;
                end else begin
                    I7628fd0a5ee3ec547c1b4798a4d76de651807424cd18f0b3b8a3bea849e6fe0d  <= I454cdecfffd5c06b833e81e8990b07a9b326eec23f31a7b6589b969f610d8ed6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idc77bba153be5873f87a4cf88c6ddc6a89bf8aa3ffcd29702126b01053f012f2 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[7] ) begin
                    I84920b6036437109dbc48865b69f249d82da5c7288a7eb7744ea7ea567e03657  <=  ~I0d0472e7c0ef483f8cb46ed393b7bcd5ea93f12dc2885368d5bf587c24198980 + 1;
                end else begin
                    I84920b6036437109dbc48865b69f249d82da5c7288a7eb7744ea7ea567e03657  <= I0d0472e7c0ef483f8cb46ed393b7bcd5ea93f12dc2885368d5bf587c24198980 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idc77bba153be5873f87a4cf88c6ddc6a89bf8aa3ffcd29702126b01053f012f2 != Ie244ea5cb57e0b4c14c0c8c22592347d1389a6b0f53b821335b821ca5130ad6e[0] ) begin
                    Iaa02b7ddfffcecb763aa916a2bc4c3aea58027c89b515c40b72214d9dd44ba21  <=  ~I33dc9b3b4f5aac0a30c5ab73b222441f5fbeedb26b7b8749a0ab253f239598d4 + 1;
                end else begin
                    Iaa02b7ddfffcecb763aa916a2bc4c3aea58027c89b515c40b72214d9dd44ba21  <= I33dc9b3b4f5aac0a30c5ab73b222441f5fbeedb26b7b8749a0ab253f239598d4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8674756fbdb78fab124727c8154adc4dcfd4674e3a4d9977d2fff619cbc42e5a != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[15] ) begin
                    I5ccf8e87b0b8e8ce9bdf4b3329e4458a628f2568184f82b998ac62ea28bc0307  <=  ~I70ea317892671f95b146604245efea2c83830d5e6b03a1dd19f2ecb28b47a9a1 + 1;
                end else begin
                    I5ccf8e87b0b8e8ce9bdf4b3329e4458a628f2568184f82b998ac62ea28bc0307  <= I70ea317892671f95b146604245efea2c83830d5e6b03a1dd19f2ecb28b47a9a1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8674756fbdb78fab124727c8154adc4dcfd4674e3a4d9977d2fff619cbc42e5a != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[7] ) begin
                    I8befad7180232073f2f7db5a3f546a5a1af79b21cc9cb00a13e266db4eebba48  <=  ~Idf920a1de857f846c8ab2646a68ee3a6053d935968cdc3d6b46308a473be4099 + 1;
                end else begin
                    I8befad7180232073f2f7db5a3f546a5a1af79b21cc9cb00a13e266db4eebba48  <= Idf920a1de857f846c8ab2646a68ee3a6053d935968cdc3d6b46308a473be4099 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I8674756fbdb78fab124727c8154adc4dcfd4674e3a4d9977d2fff619cbc42e5a != I5a07f349b1fd7d668d35583c50dfa3ceda070e5dc241bff1ecdddace6624bd57[0] ) begin
                    If8737fa82b71d9b0e7223baabca7405e148621600bdaef02e65cd7bd175b2d88  <=  ~Ifade018f22d237bddeb6fd8736ba424241846d20f2f32d2bb7fe779462ed7261 + 1;
                end else begin
                    If8737fa82b71d9b0e7223baabca7405e148621600bdaef02e65cd7bd175b2d88  <= Ifade018f22d237bddeb6fd8736ba424241846d20f2f32d2bb7fe779462ed7261 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4a3c7a36a82811aff327ec55776f5077aec859d5557df45568abcbcbb0fc5d5a != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[15] ) begin
                    Icbdf29918b91006ffdc8b68c707840ee6bb9c27779dabd372e2033888743409f  <=  ~I9318e8402c23072dcc49ace45bb9814c535167574af63bc61463059dbcb0067e + 1;
                end else begin
                    Icbdf29918b91006ffdc8b68c707840ee6bb9c27779dabd372e2033888743409f  <= I9318e8402c23072dcc49ace45bb9814c535167574af63bc61463059dbcb0067e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4a3c7a36a82811aff327ec55776f5077aec859d5557df45568abcbcbb0fc5d5a != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[7] ) begin
                    Iabc9fc6e9581216af19559d8e709ea0842cba4f29f3fdfb05bd71d6d9f7594ae  <=  ~Ic0071db5dbcb92ea14e4b31a24b9f9febc208bf86bb0634f07d9cd3763461055 + 1;
                end else begin
                    Iabc9fc6e9581216af19559d8e709ea0842cba4f29f3fdfb05bd71d6d9f7594ae  <= Ic0071db5dbcb92ea14e4b31a24b9f9febc208bf86bb0634f07d9cd3763461055 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4a3c7a36a82811aff327ec55776f5077aec859d5557df45568abcbcbb0fc5d5a != I6e5f194e3acb27a7fdd060e05aff00bb9fcd0904b3f920d7db0fee84c1534558[0] ) begin
                    Id85c2b905d61bcdc87d500d6ede3ca02d52bc3eaf278f087f27fe6f277c91262  <=  ~I64cc4cfd27023e75e5cb557e7bac31506d466107aa2cfe7809e148d8977f8393 + 1;
                end else begin
                    Id85c2b905d61bcdc87d500d6ede3ca02d52bc3eaf278f087f27fe6f277c91262  <= I64cc4cfd27023e75e5cb557e7bac31506d466107aa2cfe7809e148d8977f8393 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I931f943f5db8edf3580ebe67b3da2a0cc9a1b68ac6485930d6d9dc792bd36eb3 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[15] ) begin
                    Ief90cf0b0997823c3071eb46b636e384077579beae3d85d29e639a7719763396  <=  ~I560502a76e2a6f15d91f55a12133213d8896b50299e0a7ed30c5c5958d5f5ec5 + 1;
                end else begin
                    Ief90cf0b0997823c3071eb46b636e384077579beae3d85d29e639a7719763396  <= I560502a76e2a6f15d91f55a12133213d8896b50299e0a7ed30c5c5958d5f5ec5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I931f943f5db8edf3580ebe67b3da2a0cc9a1b68ac6485930d6d9dc792bd36eb3 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[7] ) begin
                    I4f73c51d25db7485bf4a0d63f95f14fc0661431870ce704f70cbb787eb336f09  <=  ~I7813b9f4f76a24bbf99a0f2d9cfe1d3a53eb0ec0fa5c72e06f1f86fdd1801c56 + 1;
                end else begin
                    I4f73c51d25db7485bf4a0d63f95f14fc0661431870ce704f70cbb787eb336f09  <= I7813b9f4f76a24bbf99a0f2d9cfe1d3a53eb0ec0fa5c72e06f1f86fdd1801c56 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I931f943f5db8edf3580ebe67b3da2a0cc9a1b68ac6485930d6d9dc792bd36eb3 != I09780397509ca78f4b4aed5b08cf22d8eae797d1d1864cdba4a951ac8d583c91[0] ) begin
                    I5923f41aa444bebfc18d13202747ff84e20a4753bc9cedf697b9ae8ec3418afa  <=  ~Ia81295e4b9400e1737a8a8d335ed9765fbb59b817f0251f1f032ba3e48c6bdf3 + 1;
                end else begin
                    I5923f41aa444bebfc18d13202747ff84e20a4753bc9cedf697b9ae8ec3418afa  <= Ia81295e4b9400e1737a8a8d335ed9765fbb59b817f0251f1f032ba3e48c6bdf3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[4] ) begin
                    Ifd2ca31ff3eec501f34892055a36979681d27574ed8007e4df5cc0109b71bd89  <=  ~I0b7c06b48a33586be508f2334fc3eac5befd9ff87751db1859c5f01cc6d44b15 + 1;
                end else begin
                    Ifd2ca31ff3eec501f34892055a36979681d27574ed8007e4df5cc0109b71bd89  <= I0b7c06b48a33586be508f2334fc3eac5befd9ff87751db1859c5f01cc6d44b15 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[8] ) begin
                    I6148a04ce3733485aeb6c4d20b6117eea37a510aba76ac29e82d44980bec0934  <=  ~I63860f7f2cc2e0814f98ead1e90694f745ef7a70e90f0af487d002ca46bf2c57 + 1;
                end else begin
                    I6148a04ce3733485aeb6c4d20b6117eea37a510aba76ac29e82d44980bec0934  <= I63860f7f2cc2e0814f98ead1e90694f745ef7a70e90f0af487d002ca46bf2c57 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[5] ) begin
                    Idcdcb2dd5e2f2aff0d7b362ddb4ae1ee4db08edc2c3df3589a7143bafeec0bcf  <=  ~I48e0ff7c513e9892c552947f3bb0a96d7b00d0ccfa3d7fbcf067d996b3d58dc6 + 1;
                end else begin
                    Idcdcb2dd5e2f2aff0d7b362ddb4ae1ee4db08edc2c3df3589a7143bafeec0bcf  <= I48e0ff7c513e9892c552947f3bb0a96d7b00d0ccfa3d7fbcf067d996b3d58dc6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[7] ) begin
                    Iba62c53d136b455b7d575b868f2ebd2dadc6003981aa2aae72863a0eb812bd1a  <=  ~I904078f4d964b6f66502423cb801a285f9cf21964df0a9fc1b8fdb9e35090265 + 1;
                end else begin
                    Iba62c53d136b455b7d575b868f2ebd2dadc6003981aa2aae72863a0eb812bd1a  <= I904078f4d964b6f66502423cb801a285f9cf21964df0a9fc1b8fdb9e35090265 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 != Iefcb9b5b2f238005d0f37bc519349bbbc130e3e072814ec48b4edf9c853a6913[0] ) begin
                    I4ac498dc826a9dbeaddf2f013ae7116e92dc772ea55987a4661f18e56a4123a8  <=  ~Iaed17e55ab4220ad1c1485ce0b5e5518cfc682531407f36561bfff3ed5026ff6 + 1;
                end else begin
                    I4ac498dc826a9dbeaddf2f013ae7116e92dc772ea55987a4661f18e56a4123a8  <= Iaed17e55ab4220ad1c1485ce0b5e5518cfc682531407f36561bfff3ed5026ff6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[4] ) begin
                    Id9e3ea08b52843b4a9426b735967bd4ac3d49bd67ab8fc85688b0f55e6df186a  <=  ~I101c35283ea20516f74f90cdf4ea7f1ac3a008d80dcb4b80235a17483b1f5211 + 1;
                end else begin
                    Id9e3ea08b52843b4a9426b735967bd4ac3d49bd67ab8fc85688b0f55e6df186a  <= I101c35283ea20516f74f90cdf4ea7f1ac3a008d80dcb4b80235a17483b1f5211 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[8] ) begin
                    I25c667a6616c9a94f6618166c99298b28d897f9ac8276bb85816e4b42582cdfe  <=  ~I1184b619aa3fb52506bcb002a57a421ae2f9d3a85502d2ae8132f38092c38fb5 + 1;
                end else begin
                    I25c667a6616c9a94f6618166c99298b28d897f9ac8276bb85816e4b42582cdfe  <= I1184b619aa3fb52506bcb002a57a421ae2f9d3a85502d2ae8132f38092c38fb5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[5] ) begin
                    I6c252caff8f1ab047efc25a950ce3e3ffb47a5b779e37a667c48bc1487528218  <=  ~I08fc2b9a844e2c482e2bf89714e92b5baa0ff2b9bc456c523d6360e5b5bbe2d0 + 1;
                end else begin
                    I6c252caff8f1ab047efc25a950ce3e3ffb47a5b779e37a667c48bc1487528218  <= I08fc2b9a844e2c482e2bf89714e92b5baa0ff2b9bc456c523d6360e5b5bbe2d0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[7] ) begin
                    I07087056bd31363bfb1f76f8fbeb18d1deafd5e4816ca1200d362c0797a77bb4  <=  ~I5617f2c448f426aa20d4dc124625b298648c40b73307feddaa9806bf571a71f4 + 1;
                end else begin
                    I07087056bd31363bfb1f76f8fbeb18d1deafd5e4816ca1200d362c0797a77bb4  <= I5617f2c448f426aa20d4dc124625b298648c40b73307feddaa9806bf571a71f4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 != I9835f6f38580d8765566723f5a9adbfb4935af8bf719b3e4918e1b746cf12241[0] ) begin
                    Iaadbb1b235a85c555a6f37d003e87a987b7d9b07148207555eb717b7332f67ec  <=  ~Ic9219b1b4792455d5f1c104798cfb3ace66806e030172b83b652747280a3ea8f + 1;
                end else begin
                    Iaadbb1b235a85c555a6f37d003e87a987b7d9b07148207555eb717b7332f67ec  <= Ic9219b1b4792455d5f1c104798cfb3ace66806e030172b83b652747280a3ea8f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[4] ) begin
                    Ia6414b3aff6031e10856953f6b15ffdb0971aeb680d784a7199386be15624ff6  <=  ~Ia1e3983b6aaba9149d835f0e79d761b34c608f894259979b9e02f9891b0e04be + 1;
                end else begin
                    Ia6414b3aff6031e10856953f6b15ffdb0971aeb680d784a7199386be15624ff6  <= Ia1e3983b6aaba9149d835f0e79d761b34c608f894259979b9e02f9891b0e04be ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[8] ) begin
                    I87af49f5f04df14686aef62aa27c16723af3ad05398f00e29788666b27784de5  <=  ~Ibd87e183657088945b5a8789b001bbe566368ecbc0a773fb784a3d26cb6886e1 + 1;
                end else begin
                    I87af49f5f04df14686aef62aa27c16723af3ad05398f00e29788666b27784de5  <= Ibd87e183657088945b5a8789b001bbe566368ecbc0a773fb784a3d26cb6886e1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[5] ) begin
                    I22670670d7018cb361ca0ffd92516837302d5528c26915b62d22505471ab7384  <=  ~Ic67c3bded52308b7875b1fe59eac4e253898565ad36a0f3cb39051d5a1a0289d + 1;
                end else begin
                    I22670670d7018cb361ca0ffd92516837302d5528c26915b62d22505471ab7384  <= Ic67c3bded52308b7875b1fe59eac4e253898565ad36a0f3cb39051d5a1a0289d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[7] ) begin
                    If27288056468d3ef3052303952f2e4be67796c40d6224383047d71d996f98cf3  <=  ~I496a0976329e8a4f6d29dbe1b1e9319f3f99afc9f4d3c645f264f4675b7ebf7b + 1;
                end else begin
                    If27288056468d3ef3052303952f2e4be67796c40d6224383047d71d996f98cf3  <= I496a0976329e8a4f6d29dbe1b1e9319f3f99afc9f4d3c645f264f4675b7ebf7b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 != I2266ca44e019a30bb553f955a158a5b075035c4b20a0b3fca6a3675ec79b9997[0] ) begin
                    I6afb533ec993de4f9b04007b355a9cadf08488ee6ca02aec2d7916a4c98a7fad  <=  ~I93889e1f0f60b124844920662add026c1da1fa6650f347a6a616da18e8b96c02 + 1;
                end else begin
                    I6afb533ec993de4f9b04007b355a9cadf08488ee6ca02aec2d7916a4c98a7fad  <= I93889e1f0f60b124844920662add026c1da1fa6650f347a6a616da18e8b96c02 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[4] ) begin
                    I69f7964c2f630ef03f49c2a6cac12420e0998397470245e6afaed2546b33775c  <=  ~I9bea46de6ec248c77242ae2154d5c6e1dc17ff892dc903bd685badcbaf62291e + 1;
                end else begin
                    I69f7964c2f630ef03f49c2a6cac12420e0998397470245e6afaed2546b33775c  <= I9bea46de6ec248c77242ae2154d5c6e1dc17ff892dc903bd685badcbaf62291e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[8] ) begin
                    I7e269b2e2d9ec70c47570bad75bce0ddf53e85e3cb4ba87f784ca520c5ff1084  <=  ~I88a966d14bd155320f8f49d164cf93516a3822b9098c6417bcdb8a64f9eb1a38 + 1;
                end else begin
                    I7e269b2e2d9ec70c47570bad75bce0ddf53e85e3cb4ba87f784ca520c5ff1084  <= I88a966d14bd155320f8f49d164cf93516a3822b9098c6417bcdb8a64f9eb1a38 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[5] ) begin
                    Ief691d56b56a000651b0a4c6cc9f26bc44da82f4a6382550d96ea4101b81ecb9  <=  ~I23c475c49d2504d72c81fcf2a1ca3122e6dfbc9f1e9faa0253d0d36c27881126 + 1;
                end else begin
                    Ief691d56b56a000651b0a4c6cc9f26bc44da82f4a6382550d96ea4101b81ecb9  <= I23c475c49d2504d72c81fcf2a1ca3122e6dfbc9f1e9faa0253d0d36c27881126 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[7] ) begin
                    I4fa5ada2d589c7a90e700745aba8e09edcfb0252f532e4c74eb0809c712a36f0  <=  ~Ib19a40aaae7bc965afa2506ee77fab296894319861766d0f6ede0e69e01ad17a + 1;
                end else begin
                    I4fa5ada2d589c7a90e700745aba8e09edcfb0252f532e4c74eb0809c712a36f0  <= Ib19a40aaae7bc965afa2506ee77fab296894319861766d0f6ede0e69e01ad17a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 != I684ec077e37638f022f10b5eb31403e6f9117a83a606f2a5013c2c33b8d1a8ab[0] ) begin
                    I01313177417c899543a67763ede925dea3ee58ef4a31714ad15a7a3746bb5be5  <=  ~Ie10eac9c8e0f2526d443d3c8d9c007e29481ae4fd9bed2afac5a0861f80705c0 + 1;
                end else begin
                    I01313177417c899543a67763ede925dea3ee58ef4a31714ad15a7a3746bb5be5  <= Ie10eac9c8e0f2526d443d3c8d9c007e29481ae4fd9bed2afac5a0861f80705c0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b3ff601c78f414f5f48cde79235444d13872a0527c054356b3af150315b0949 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[16] ) begin
                    I1d8a992801d3f6a457848578ce286b496d4e2a69937344bdcbab4e8b1af1fe4e  <=  ~I873fa9e73fcb148c0eab3dfc8d6163714e0a0dd5889d5d5dd73244c4f700f3bf + 1;
                end else begin
                    I1d8a992801d3f6a457848578ce286b496d4e2a69937344bdcbab4e8b1af1fe4e  <= I873fa9e73fcb148c0eab3dfc8d6163714e0a0dd5889d5d5dd73244c4f700f3bf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b3ff601c78f414f5f48cde79235444d13872a0527c054356b3af150315b0949 != I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[6] ) begin
                    Id7dcf87d2a40e82e7f01327d834d5207ae5873a7e5133c3dddead9d0cb9703f9  <=  ~I2d891a9027bcd15bb7deaddca0e282e872204770ad4e90ffcd4826beb3c492cf + 1;
                end else begin
                    Id7dcf87d2a40e82e7f01327d834d5207ae5873a7e5133c3dddead9d0cb9703f9  <= I2d891a9027bcd15bb7deaddca0e282e872204770ad4e90ffcd4826beb3c492cf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7b3ff601c78f414f5f48cde79235444d13872a0527c054356b3af150315b0949 != I9331428911b817ea45d1b5ae75eb3ee6e05c189785c995e5d2625f12ce4e0846[0] ) begin
                    Ibd0ba147d1a08acea707b8c60da14ebcc4ad62e67ef26634777b5dae38af6d61  <=  ~Ieae87e6a29536e19a2589665b2af980e34700c9a614fe1b7c4704a7a538a8f8c + 1;
                end else begin
                    Ibd0ba147d1a08acea707b8c60da14ebcc4ad62e67ef26634777b5dae38af6d61  <= Ieae87e6a29536e19a2589665b2af980e34700c9a614fe1b7c4704a7a538a8f8c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I434491ac49be9939ffdcf469991bc3d23ef217b8414c677d78ec9a062e74ba07 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[16] ) begin
                    Iaea7277e745e05f803325e0f19dbc5a54234878a9a3cb2cedcc013e3942e9cc0  <=  ~Ia30f6d6396acef716d7383513ac1f4caface96330dcacfdc5302bbb0408697cb + 1;
                end else begin
                    Iaea7277e745e05f803325e0f19dbc5a54234878a9a3cb2cedcc013e3942e9cc0  <= Ia30f6d6396acef716d7383513ac1f4caface96330dcacfdc5302bbb0408697cb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I434491ac49be9939ffdcf469991bc3d23ef217b8414c677d78ec9a062e74ba07 != I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[6] ) begin
                    I2cb1ae23e53b89ca0fd3d1df98b32d5b9e478e9eb579b0875981a6b056e8ef4e  <=  ~I794ed9d1df776d692b623e89b6d6ade5d265c9869957ddd8e256061bb513d7ea + 1;
                end else begin
                    I2cb1ae23e53b89ca0fd3d1df98b32d5b9e478e9eb579b0875981a6b056e8ef4e  <= I794ed9d1df776d692b623e89b6d6ade5d265c9869957ddd8e256061bb513d7ea ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I434491ac49be9939ffdcf469991bc3d23ef217b8414c677d78ec9a062e74ba07 != I7769e8ceb72790c37b351c32983860280aef172974d19a2e99348607863a97d4[0] ) begin
                    I1e92e18a915678cc96aa493a00627dffecbd341dc8e022615610061e52c1ac3f  <=  ~Iaaffc28ce6e25495dfad668af2f560c988f5a5abb76db94b71563231400c28b1 + 1;
                end else begin
                    I1e92e18a915678cc96aa493a00627dffecbd341dc8e022615610061e52c1ac3f  <= Iaaffc28ce6e25495dfad668af2f560c988f5a5abb76db94b71563231400c28b1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icd717b9b3dc725b8579e62b042051399a3b21cc10076de8e0bae480fcd24d607 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[16] ) begin
                    I7f6b89a61d6313029102fc48e92a54ffdece30e9eac1191d840c488be69d8223  <=  ~I45324df36dd601c219634e39418995a9ab1bd58be03cb5dee89ac2d01bec1dde + 1;
                end else begin
                    I7f6b89a61d6313029102fc48e92a54ffdece30e9eac1191d840c488be69d8223  <= I45324df36dd601c219634e39418995a9ab1bd58be03cb5dee89ac2d01bec1dde ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icd717b9b3dc725b8579e62b042051399a3b21cc10076de8e0bae480fcd24d607 != I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[6] ) begin
                    I463662fa980f8a5e4be086aa5f37db53b1d6ea8dfe11725b8c407f779a168998  <=  ~Idc26ae0a7d9ab347f3c75ed2ac7c48f6937f9cc035d46be065fb4b15699cc989 + 1;
                end else begin
                    I463662fa980f8a5e4be086aa5f37db53b1d6ea8dfe11725b8c407f779a168998  <= Idc26ae0a7d9ab347f3c75ed2ac7c48f6937f9cc035d46be065fb4b15699cc989 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icd717b9b3dc725b8579e62b042051399a3b21cc10076de8e0bae480fcd24d607 != If09c36408407b246848b29df63e789fd1041815243beb4f27db0e774e853f1cd[0] ) begin
                    Ia7b91fa4a1ef16f859ee162b91daedc97927244dc19aaedede898049daf85a19  <=  ~I8e22237e0bc0b24825cc53a9b88f0ad973a825d25aee1abcfddcbb6ddc14ea48 + 1;
                end else begin
                    Ia7b91fa4a1ef16f859ee162b91daedc97927244dc19aaedede898049daf85a19  <= I8e22237e0bc0b24825cc53a9b88f0ad973a825d25aee1abcfddcbb6ddc14ea48 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0c556fb5fa4a1297825cab8dc64089faa86f1cbe67bf106748d927849e16e007 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[16] ) begin
                    I295d7aef060ca978805bdf65138e5bf134551eda9c396a22165a77a3091dfd28  <=  ~Ieff55ba27500b6d175abdc30224d7d4c703ff1ce6a3b5d86475b739903839b52 + 1;
                end else begin
                    I295d7aef060ca978805bdf65138e5bf134551eda9c396a22165a77a3091dfd28  <= Ieff55ba27500b6d175abdc30224d7d4c703ff1ce6a3b5d86475b739903839b52 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0c556fb5fa4a1297825cab8dc64089faa86f1cbe67bf106748d927849e16e007 != I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[6] ) begin
                    Ibc3e77c4d6cb28599b7a21c7992802beffb168f54d8dfa650750ffdc6730df29  <=  ~I79948c8c3800c594e6e33eff537e1b38872775f3674ce78ad963f09de0091486 + 1;
                end else begin
                    Ibc3e77c4d6cb28599b7a21c7992802beffb168f54d8dfa650750ffdc6730df29  <= I79948c8c3800c594e6e33eff537e1b38872775f3674ce78ad963f09de0091486 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0c556fb5fa4a1297825cab8dc64089faa86f1cbe67bf106748d927849e16e007 != I533b63eedc528cb36abc0a469b66b144a6ae5122c038eef85d8d0557c3dff3ea[0] ) begin
                    I9918d91748722a47f8526008bc3fd4c498bc80205211d5c92acbc511fdb667bf  <=  ~Icf4362e74e763b339d2ba9634282b8441d0c293aacbc2879f95a53ef1a2122e6 + 1;
                end else begin
                    I9918d91748722a47f8526008bc3fd4c498bc80205211d5c92acbc511fdb667bf  <= Icf4362e74e763b339d2ba9634282b8441d0c293aacbc2879f95a53ef1a2122e6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[18] ) begin
                    I8b5ee5d271abdbdc518ce02f900da21e858d3e2530585fd859690a1a71502434  <=  ~Id6a3fad936fae13ba6503265a6a9a2bd1c54dc3fcb3d196623bf8aad32225687 + 1;
                end else begin
                    I8b5ee5d271abdbdc518ce02f900da21e858d3e2530585fd859690a1a71502434  <= Id6a3fad936fae13ba6503265a6a9a2bd1c54dc3fcb3d196623bf8aad32225687 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[5] ) begin
                    I6b2620e847ea73b8618ac7bdcd8236c4278de3bef0bf1511ee9779306438fa38  <=  ~Ic26999f764390a0c1461876b7687ee02acb7586ae1e24d171988084ca9d4aa82 + 1;
                end else begin
                    I6b2620e847ea73b8618ac7bdcd8236c4278de3bef0bf1511ee9779306438fa38  <= Ic26999f764390a0c1461876b7687ee02acb7586ae1e24d171988084ca9d4aa82 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[8] ) begin
                    I2647390c3800518f2251794a7ee4aa2d71ca9589534cf73eda0accbd2b3342da  <=  ~Ic77bba83655ba517bc6313df02ee80ace5ba5e383e3794f971225d42bdf82690 + 1;
                end else begin
                    I2647390c3800518f2251794a7ee4aa2d71ca9589534cf73eda0accbd2b3342da  <= Ic77bba83655ba517bc6313df02ee80ace5ba5e383e3794f971225d42bdf82690 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e != I051e3b709db2e7861d31165ec1e5ee679f1e6dffa5a951072831ce479c16f27f[0] ) begin
                    I95d109e37a87827de1455b5ec479dda78a0218cb9db245b80710cdb1e8ead67a  <=  ~I01ac098466c350975d0ecff2227564446e39a21fd133aab22628a9cf3a866b90 + 1;
                end else begin
                    I95d109e37a87827de1455b5ec479dda78a0218cb9db245b80710cdb1e8ead67a  <= I01ac098466c350975d0ecff2227564446e39a21fd133aab22628a9cf3a866b90 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[18] ) begin
                    If49d6a59c1d539e369406ee4e8a2ebb30199f46c335584e62921f98fd811001d  <=  ~I97389ae6e03b0e2bee0e882909d2adf1aa34eecf73084ceab73088e850c24e87 + 1;
                end else begin
                    If49d6a59c1d539e369406ee4e8a2ebb30199f46c335584e62921f98fd811001d  <= I97389ae6e03b0e2bee0e882909d2adf1aa34eecf73084ceab73088e850c24e87 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[5] ) begin
                    I77e34c24ea46e99b6bfc0f960d428d6ba3ea4f9261d5a183d83c386f259ab431  <=  ~I059c355ce17871c1a494b1a39b4ad3408ab5d28b886b143e04c71a29731f4651 + 1;
                end else begin
                    I77e34c24ea46e99b6bfc0f960d428d6ba3ea4f9261d5a183d83c386f259ab431  <= I059c355ce17871c1a494b1a39b4ad3408ab5d28b886b143e04c71a29731f4651 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[8] ) begin
                    I78f0dcc6533ef218ce6959768639c983d2119dd518e988eb3dcd6f0b4de98c82  <=  ~Ie5a7256fb2ee0e45b0cc306c46856bd7cc606efccd221b75d515f608ad567603 + 1;
                end else begin
                    I78f0dcc6533ef218ce6959768639c983d2119dd518e988eb3dcd6f0b4de98c82  <= Ie5a7256fb2ee0e45b0cc306c46856bd7cc606efccd221b75d515f608ad567603 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec != I2fa018ce903921d0a174a63dbbb29eea8d5700b376335b2ba9bd448e8782018a[0] ) begin
                    Ia0c7162290e415f24699688e45850c243397b5cccf07daf0398dda04810b0690  <=  ~Ib419bb101d14a1958ca5b3a7c6a72d8fc15ca6e217fcac0f7eb84c776f3b0826 + 1;
                end else begin
                    Ia0c7162290e415f24699688e45850c243397b5cccf07daf0398dda04810b0690  <= Ib419bb101d14a1958ca5b3a7c6a72d8fc15ca6e217fcac0f7eb84c776f3b0826 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[18] ) begin
                    Icf0b2747a9e17f2d2672f7a17111c6bf54bed7d8fedcb5260f25fdc4280ae727  <=  ~Ie5a479b36bb003e0b2d92a68e955c1906c3969ee52a96b4aef5a84bc275f3f9f + 1;
                end else begin
                    Icf0b2747a9e17f2d2672f7a17111c6bf54bed7d8fedcb5260f25fdc4280ae727  <= Ie5a479b36bb003e0b2d92a68e955c1906c3969ee52a96b4aef5a84bc275f3f9f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[5] ) begin
                    Iaf94ae58c1d9c9206d02651cd03cf2e02bba505f76b849158530a38382396ffa  <=  ~I380a702cee9dcf67af75101568b0a417c567c5ebc9e777dd1fd2d297c2455e90 + 1;
                end else begin
                    Iaf94ae58c1d9c9206d02651cd03cf2e02bba505f76b849158530a38382396ffa  <= I380a702cee9dcf67af75101568b0a417c567c5ebc9e777dd1fd2d297c2455e90 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[8] ) begin
                    I3a9293b8f323c7e097a099fa6beb33ca299723796aec9396365d43334eb55e35  <=  ~I44aed07314ea5c6ed70e468558116a9b956c9a2d67e52229ac85b62c1b511d36 + 1;
                end else begin
                    I3a9293b8f323c7e097a099fa6beb33ca299723796aec9396365d43334eb55e35  <= I44aed07314ea5c6ed70e468558116a9b956c9a2d67e52229ac85b62c1b511d36 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b != I36e06c1d77080ff75778f3dfa4ed60e66f9a3bedc39b214e3fdb5b6c21f1cd3e[0] ) begin
                    Ib9dc17b2b9fc7c228eba40cf625a49a27ec16f8c8a91957de14fb6849ea49212  <=  ~I7f63700c8702ba858d076a1901ee015cd80dd29b33e109b7ce64aa14493461af + 1;
                end else begin
                    Ib9dc17b2b9fc7c228eba40cf625a49a27ec16f8c8a91957de14fb6849ea49212  <= I7f63700c8702ba858d076a1901ee015cd80dd29b33e109b7ce64aa14493461af ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[18] ) begin
                    I84238bd7e53e0dd7ba07efd813661c8cd1648b76c44665dfe51fd07dfaa9b249  <=  ~If8bbc0d7554b094c7dbd8b4a06c4ef791cd6e66621e4c3b97464052276957603 + 1;
                end else begin
                    I84238bd7e53e0dd7ba07efd813661c8cd1648b76c44665dfe51fd07dfaa9b249  <= If8bbc0d7554b094c7dbd8b4a06c4ef791cd6e66621e4c3b97464052276957603 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[5] ) begin
                    I6f63c71eab6c2d7e3eb41fd78c9e18d6362d2dd4100c72b43d3e4b9d06663165  <=  ~Ib65f0444b24cc43c4ebe5dc5fb7a2e0aad7c8d125bf92c527ba5dabd52d8f98a + 1;
                end else begin
                    I6f63c71eab6c2d7e3eb41fd78c9e18d6362d2dd4100c72b43d3e4b9d06663165  <= Ib65f0444b24cc43c4ebe5dc5fb7a2e0aad7c8d125bf92c527ba5dabd52d8f98a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[8] ) begin
                    Id165331f616d7e8f347cbe46daff955009fef6f8c0310c64c01dd35990231279  <=  ~I088890dd5f7391be17333396dc9b8cba40ddef39e657378c312707e1ea43bb56 + 1;
                end else begin
                    Id165331f616d7e8f347cbe46daff955009fef6f8c0310c64c01dd35990231279  <= I088890dd5f7391be17333396dc9b8cba40ddef39e657378c312707e1ea43bb56 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e != Id647e3bd88fdc7a3642092d071f66f74657c8364937caf63c723f1e027c157bc[0] ) begin
                    Ied32ced79448b3f92faf0dca1673559e07372ec338e8c51a750be1c6975a298e  <=  ~I64fcddc23b1b1d72f4a5cd8707f8ec3dfb77bd105d279d01a99750b9ec4894d6 + 1;
                end else begin
                    Ied32ced79448b3f92faf0dca1673559e07372ec338e8c51a750be1c6975a298e  <= I64fcddc23b1b1d72f4a5cd8707f8ec3dfb77bd105d279d01a99750b9ec4894d6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id3bfe7fc5e0a1ea258f912127a3c77f7cc5ad791dc6166266f64c574b8ed0e81 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[17] ) begin
                    I9471414594b824d60836981bf4b9931c135520ad1ae7dea177e0bc591c2572c2  <=  ~I323a7ad384b7514bf52fc27d18b29da7effc88c35471be18c85d0b61ece11db3 + 1;
                end else begin
                    I9471414594b824d60836981bf4b9931c135520ad1ae7dea177e0bc591c2572c2  <= I323a7ad384b7514bf52fc27d18b29da7effc88c35471be18c85d0b61ece11db3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id3bfe7fc5e0a1ea258f912127a3c77f7cc5ad791dc6166266f64c574b8ed0e81 != Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[4] ) begin
                    Iaa0b6d0f2fe24db548975f410ac5b79f687b7646169247f3891ce9e4644ee0fa  <=  ~Iede33454e4e4f5856e3700d92d14d4b4ee573de70aa6715525cb1164348e6561 + 1;
                end else begin
                    Iaa0b6d0f2fe24db548975f410ac5b79f687b7646169247f3891ce9e4644ee0fa  <= Iede33454e4e4f5856e3700d92d14d4b4ee573de70aa6715525cb1164348e6561 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id3bfe7fc5e0a1ea258f912127a3c77f7cc5ad791dc6166266f64c574b8ed0e81 != I015b73e7e4bc4c2a3073a304e58d24f5c8c32e90299f004bc0f75eb9e18e6d41[0] ) begin
                    Iaddb000276bde734c13ec1395f06c1b3bf5606ad5cb138579d711cecf26ac88a  <=  ~I6254bd01448c9d8e8b348c9cf6f62da72b3e66c76cfc692be2250a30039c48db + 1;
                end else begin
                    Iaddb000276bde734c13ec1395f06c1b3bf5606ad5cb138579d711cecf26ac88a  <= I6254bd01448c9d8e8b348c9cf6f62da72b3e66c76cfc692be2250a30039c48db ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I370bb7df3320249e804ee9d3d371b1e82809433e4f7e00f74ea0ab59252f4176 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[17] ) begin
                    I73a855a590363c762c34008e77f73f961950c0dd71b795acab3adf40c4540453  <=  ~Ib50a67b0b1f097d85a05aefb1686e6d51cbbda0406226d20772af68de6e6d139 + 1;
                end else begin
                    I73a855a590363c762c34008e77f73f961950c0dd71b795acab3adf40c4540453  <= Ib50a67b0b1f097d85a05aefb1686e6d51cbbda0406226d20772af68de6e6d139 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I370bb7df3320249e804ee9d3d371b1e82809433e4f7e00f74ea0ab59252f4176 != Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[4] ) begin
                    I1cf0e3016bbd2d8e5debffedb198273a2d019ce75f2f8352a285d17264d262f0  <=  ~Ib0809c22530a4fef601b75ff7573a7e9606b2da1938ed0918b43a958b9c2ddb9 + 1;
                end else begin
                    I1cf0e3016bbd2d8e5debffedb198273a2d019ce75f2f8352a285d17264d262f0  <= Ib0809c22530a4fef601b75ff7573a7e9606b2da1938ed0918b43a958b9c2ddb9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I370bb7df3320249e804ee9d3d371b1e82809433e4f7e00f74ea0ab59252f4176 != I7c211cef6a581c5a6871d4c9a2b7ba29a9d05d36b0a758106e006caebfc592e5[0] ) begin
                    I211ada7f9095ced6b3d20f8f7f67b56cd2e73595481ed5d4c08175ca874d16ae  <=  ~Ia0febef423616e7d4ab3957eea2ba1de8a8bba8b027652658ac2ab5aab11b9bf + 1;
                end else begin
                    I211ada7f9095ced6b3d20f8f7f67b56cd2e73595481ed5d4c08175ca874d16ae  <= Ia0febef423616e7d4ab3957eea2ba1de8a8bba8b027652658ac2ab5aab11b9bf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d17552542ca2452e4f458fbd0aacb1a5b62ebee4be942ac561b87376658c9d8 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[17] ) begin
                    Ia28f68b737aaaaa6b98aa5e9696b937e564754edef217740c414c16fe2e485b6  <=  ~I8cdc972ad763857aa9a0cf1145ac106bedcf7897da19e06cdac06cbbc52e0141 + 1;
                end else begin
                    Ia28f68b737aaaaa6b98aa5e9696b937e564754edef217740c414c16fe2e485b6  <= I8cdc972ad763857aa9a0cf1145ac106bedcf7897da19e06cdac06cbbc52e0141 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d17552542ca2452e4f458fbd0aacb1a5b62ebee4be942ac561b87376658c9d8 != I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[4] ) begin
                    I9a4f77c8ba9a40c1b543070a42451ed37c0f22850a4734cdda393e69c7b54733  <=  ~I10d197005aafecec4bf8c18547bda5a551dac520da311ee42db394ac67f413f1 + 1;
                end else begin
                    I9a4f77c8ba9a40c1b543070a42451ed37c0f22850a4734cdda393e69c7b54733  <= I10d197005aafecec4bf8c18547bda5a551dac520da311ee42db394ac67f413f1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d17552542ca2452e4f458fbd0aacb1a5b62ebee4be942ac561b87376658c9d8 != I3f2014435aac47a3c807e9ad3f0829179f9285582b7ff2e3bae250a25e800aee[0] ) begin
                    I0d49182fe7486bcf54c8f68904b4b90436de6f3bc42fab67a4e47f61154e22c4  <=  ~Idb166c946a1916a593a1931a1651288e452553572b5b4e272aaa917a4afbc42e + 1;
                end else begin
                    I0d49182fe7486bcf54c8f68904b4b90436de6f3bc42fab67a4e47f61154e22c4  <= Idb166c946a1916a593a1931a1651288e452553572b5b4e272aaa917a4afbc42e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5ae887c145ca6af35eef2229e55c297f4b6ffe0a2cc47e55e6dbf09e1f11a9e7 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[17] ) begin
                    Ic94e7c887d7f24b573b470820c36fe8a0fef750e2c46675f8867d78f2100f1f9  <=  ~I3ca7faf1b6e8e04fdab54e1a4b313720f91992013d31b492f9aa49e54676aea4 + 1;
                end else begin
                    Ic94e7c887d7f24b573b470820c36fe8a0fef750e2c46675f8867d78f2100f1f9  <= I3ca7faf1b6e8e04fdab54e1a4b313720f91992013d31b492f9aa49e54676aea4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5ae887c145ca6af35eef2229e55c297f4b6ffe0a2cc47e55e6dbf09e1f11a9e7 != I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[4] ) begin
                    I926233df0c5e8461173cedabbf49fead4b0ab577d82f2585af3a1fb6e3130e21  <=  ~I77a2d0c0f26725cfe51712e4d1fd8663cdcd4668405e3fabd33e72bf7d008343 + 1;
                end else begin
                    I926233df0c5e8461173cedabbf49fead4b0ab577d82f2585af3a1fb6e3130e21  <= I77a2d0c0f26725cfe51712e4d1fd8663cdcd4668405e3fabd33e72bf7d008343 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5ae887c145ca6af35eef2229e55c297f4b6ffe0a2cc47e55e6dbf09e1f11a9e7 != Ib27fb4891a6edd486a99f23a750057de12a5a3e3fc6a5fad7976aa7e961e0c54[0] ) begin
                    If79b91295d25c503f6bf5ca7c6eebd2ebf6807dd9990ce31e844cee0d8f89dac  <=  ~I3c9445224e3dc806a499c5a5faae2cd5691cfb5497852d3aced39ec164d9a5ce + 1;
                end else begin
                    If79b91295d25c503f6bf5ca7c6eebd2ebf6807dd9990ce31e844cee0d8f89dac  <= I3c9445224e3dc806a499c5a5faae2cd5691cfb5497852d3aced39ec164d9a5ce ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[6] ) begin
                    Ia0a40c2a77389cda4a8333aeaecf37a2595fbda87854a43162ad1299544bd9e6  <=  ~If86de9d134174799b06582013809be1a492e36de3aeae4cab7bdd6a827223976 + 1;
                end else begin
                    Ia0a40c2a77389cda4a8333aeaecf37a2595fbda87854a43162ad1299544bd9e6  <= If86de9d134174799b06582013809be1a492e36de3aeae4cab7bdd6a827223976 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[9] ) begin
                    If64a23ad02d1da21fe63cb33f95d37c576739eb181b0fe50d7a5101817b4ede9  <=  ~I6c7e61c506c8d841d4747e5963d49e0237b106ba6cb15a0fc9e4680ccab02c5e + 1;
                end else begin
                    If64a23ad02d1da21fe63cb33f95d37c576739eb181b0fe50d7a5101817b4ede9  <= I6c7e61c506c8d841d4747e5963d49e0237b106ba6cb15a0fc9e4680ccab02c5e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[9] ) begin
                    Ic1211f3a0703e281ce073a20afbabe9b2a698d1cf74f07f099d21fd89ffc8908  <=  ~I9c17caab5e5aed3ddf7a867cf514cdb5f65c3591789f1058a756265f97aabea9 + 1;
                end else begin
                    Ic1211f3a0703e281ce073a20afbabe9b2a698d1cf74f07f099d21fd89ffc8908  <= I9c17caab5e5aed3ddf7a867cf514cdb5f65c3591789f1058a756265f97aabea9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 != I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[7] ) begin
                    I2c316e8b8cb6b499a7a8fbb513b3067829197cfacee877c35874a2ec686ada4a  <=  ~Ic818ff3260f1543c8d940d36c72d644a7a3a243220548792289117ca6a793c02 + 1;
                end else begin
                    I2c316e8b8cb6b499a7a8fbb513b3067829197cfacee877c35874a2ec686ada4a  <= Ic818ff3260f1543c8d940d36c72d644a7a3a243220548792289117ca6a793c02 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 != Ib58cd067e009a5f4b72af8cfb1e5c49c18f51a2ad8880f65aee683bf8ecd40ad[0] ) begin
                    Iec1d04d20ec09595743b7a35860b5cb2ec862c20da87c6f899284069c60bdd71  <=  ~Ief965ff00c0da0a12a68cadf50622567e99dd688e9bb810dd46f69e3eacb7285 + 1;
                end else begin
                    Iec1d04d20ec09595743b7a35860b5cb2ec862c20da87c6f899284069c60bdd71  <= Ief965ff00c0da0a12a68cadf50622567e99dd688e9bb810dd46f69e3eacb7285 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[6] ) begin
                    I23c91b29deaa2df1f4d96e343f6fb852a2b594937a4f62dc4be1fcbe0347c439  <=  ~Ib4d1942b7949b0a4e79441e13e3b6b7b36bbb136c2bed6ad1adba30a840f4b55 + 1;
                end else begin
                    I23c91b29deaa2df1f4d96e343f6fb852a2b594937a4f62dc4be1fcbe0347c439  <= Ib4d1942b7949b0a4e79441e13e3b6b7b36bbb136c2bed6ad1adba30a840f4b55 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[9] ) begin
                    I52698fa0d5291f0dc20fb5f24c33e968ea63f47765bb7d231720330b624b2fae  <=  ~Idc7991125ae81f1c0d5f221c7fccd90e5aaf92e72e0421aa687e6c1e0f8afa9d + 1;
                end else begin
                    I52698fa0d5291f0dc20fb5f24c33e968ea63f47765bb7d231720330b624b2fae  <= Idc7991125ae81f1c0d5f221c7fccd90e5aaf92e72e0421aa687e6c1e0f8afa9d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[9] ) begin
                    I0c23517b9814053cd1f89a8b80a64fcff6ae65937dc97199c0b79ba8f7a34ff3  <=  ~Ic1e2fa322b42a15a886ec6ba9f67656a39c8bd6a13af883081336da43d9d0406 + 1;
                end else begin
                    I0c23517b9814053cd1f89a8b80a64fcff6ae65937dc97199c0b79ba8f7a34ff3  <= Ic1e2fa322b42a15a886ec6ba9f67656a39c8bd6a13af883081336da43d9d0406 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 != I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[7] ) begin
                    Ic8f640e7a0c71ddb20a985259b5e48746d28d2898383765c3b78c577f281d27f  <=  ~Ibdbd014d7bbe12aa223eaa43939e3459f35b9970ed075d4733932cb66042d281 + 1;
                end else begin
                    Ic8f640e7a0c71ddb20a985259b5e48746d28d2898383765c3b78c577f281d27f  <= Ibdbd014d7bbe12aa223eaa43939e3459f35b9970ed075d4733932cb66042d281 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 != I7e40bd6625b1d7deff82f67d46817c7af70f1da57561ab528b553b3d244b3f1d[0] ) begin
                    I2126b1597a95d7aeb7d20d4e0f4270e1fc5cb0fe6eb5003b05abbb7e5e9a2819  <=  ~I4dcdb2c22db70cdfa468f9249fea4262e91120e0d995981b34919e26c9b5bc5b + 1;
                end else begin
                    I2126b1597a95d7aeb7d20d4e0f4270e1fc5cb0fe6eb5003b05abbb7e5e9a2819  <= I4dcdb2c22db70cdfa468f9249fea4262e91120e0d995981b34919e26c9b5bc5b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[6] ) begin
                    Id2cf59876d070e0f34ee834d2691f7fbdb039bc9273329e2ce8eddfe736f0a45  <=  ~I2f6966ba5ca0aea5cb187d9d90bb6b743b80bbc7fc4547396dac13a22603e7d4 + 1;
                end else begin
                    Id2cf59876d070e0f34ee834d2691f7fbdb039bc9273329e2ce8eddfe736f0a45  <= I2f6966ba5ca0aea5cb187d9d90bb6b743b80bbc7fc4547396dac13a22603e7d4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[9] ) begin
                    If17c7df712b5dd40132ac60628bd514bc70092122a0cb89ba7d4559439779fc9  <=  ~Ibec37c7599a7f7cad52a48cb44ea0ffe117ac5ea206590a3eb8a2c661913c9ad + 1;
                end else begin
                    If17c7df712b5dd40132ac60628bd514bc70092122a0cb89ba7d4559439779fc9  <= Ibec37c7599a7f7cad52a48cb44ea0ffe117ac5ea206590a3eb8a2c661913c9ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[9] ) begin
                    Ia6391e6b0ad4d9fe4136b90a57d121f2b5f16ed4662429f1b85677591fee37a6  <=  ~Ieea63392582d451f7570a458bd235afaec2d11a7427d4e706bc1d73128993792 + 1;
                end else begin
                    Ia6391e6b0ad4d9fe4136b90a57d121f2b5f16ed4662429f1b85677591fee37a6  <= Ieea63392582d451f7570a458bd235afaec2d11a7427d4e706bc1d73128993792 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 != I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[7] ) begin
                    I1187dbcc72f33b4cc3442982af526be4cfca1b5ac65be943d4ec380421632117  <=  ~I2fc14612ec75b59c28fa90d7a5bfd1bce6d5d1fe0c46ba45f77ee2f9aa9e481a + 1;
                end else begin
                    I1187dbcc72f33b4cc3442982af526be4cfca1b5ac65be943d4ec380421632117  <= I2fc14612ec75b59c28fa90d7a5bfd1bce6d5d1fe0c46ba45f77ee2f9aa9e481a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 != I01949f24f74578cb63dd095e8ce639ce0d273c14da81e75d00097535e391aa4c[0] ) begin
                    I72a115d9b3659f31366e1d73d6d9a0793e20be233c3ccab2b513fd79786224bb  <=  ~I876dccf88204e4113c5f80bdf348624dfbd5a1439638577670da4c6afe1d5f70 + 1;
                end else begin
                    I72a115d9b3659f31366e1d73d6d9a0793e20be233c3ccab2b513fd79786224bb  <= I876dccf88204e4113c5f80bdf348624dfbd5a1439638577670da4c6afe1d5f70 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[6] ) begin
                    I930ad334ce972f0b5dbddf698f6101a196d8072e90d8144b31ce3f4b48a73e59  <=  ~If0c1eced668b91b966c13a44ef09ca1209f96723c7e3d030a757d45d0b61141f + 1;
                end else begin
                    I930ad334ce972f0b5dbddf698f6101a196d8072e90d8144b31ce3f4b48a73e59  <= If0c1eced668b91b966c13a44ef09ca1209f96723c7e3d030a757d45d0b61141f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[9] ) begin
                    Ie05c1da46b594d3c94aac179f6c98334d0d667cea08108719b44541b7b0a2049  <=  ~I5f3fc42a6dc35a49dba82814b80238d6a9f6e9c8cfddd4d72749a3197115b969 + 1;
                end else begin
                    Ie05c1da46b594d3c94aac179f6c98334d0d667cea08108719b44541b7b0a2049  <= I5f3fc42a6dc35a49dba82814b80238d6a9f6e9c8cfddd4d72749a3197115b969 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[9] ) begin
                    I2d2137ac29a7c23160dedc43e9caf010f72f7d08b057e49fcac89984e616fa5a  <=  ~I677e11f6dcc443a45cc24e28c955adce7dc006e6b26e0ade792740c59d91ed6d + 1;
                end else begin
                    I2d2137ac29a7c23160dedc43e9caf010f72f7d08b057e49fcac89984e616fa5a  <= I677e11f6dcc443a45cc24e28c955adce7dc006e6b26e0ade792740c59d91ed6d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 != I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[7] ) begin
                    Iad7f008b5f08f3ba94a0832261fb4add17f0897e3c7d54a250377b813e284331  <=  ~I703d9bd8f5b9435c814d93ae7e2327a45e0febce37b67b770c2b93f30ba39972 + 1;
                end else begin
                    Iad7f008b5f08f3ba94a0832261fb4add17f0897e3c7d54a250377b813e284331  <= I703d9bd8f5b9435c814d93ae7e2327a45e0febce37b67b770c2b93f30ba39972 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 != Id8f2a0d3524b27621ca5a576bf16e15789e6257060225da04da2a5fcc8cf751e[0] ) begin
                    I469b0bcfe9cfc27a8596782bab479f30aedaa132a5cd404feb1fec4b52a17d3a  <=  ~I4d518a62a0a46b493ab538e6ccaec00b9b2cd08aba9695482997b884ae7b006e + 1;
                end else begin
                    I469b0bcfe9cfc27a8596782bab479f30aedaa132a5cd404feb1fec4b52a17d3a  <= I4d518a62a0a46b493ab538e6ccaec00b9b2cd08aba9695482997b884ae7b006e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00fca56df853315156adf3a6a5cdecaf6256b108f16f65b1e93272f0c7796e9c != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[19] ) begin
                    I54e64fd01d9aff7ddfc4babeff6703891da38578bb141d250c4ef5949d818cfb  <=  ~I67fa42eadbdacb43b464b7246fbecac6c261d3cc37d501efdc1e83b9b1ff6055 + 1;
                end else begin
                    I54e64fd01d9aff7ddfc4babeff6703891da38578bb141d250c4ef5949d818cfb  <= I67fa42eadbdacb43b464b7246fbecac6c261d3cc37d501efdc1e83b9b1ff6055 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00fca56df853315156adf3a6a5cdecaf6256b108f16f65b1e93272f0c7796e9c != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[8] ) begin
                    I71c6f88cbabd48d41f42f2b16170c8955b79d20b8a8b211e174d1c1473567ad4  <=  ~Idb5ffff327b8edefda5ee44436f5f31deac21a01781b65e2429b1e1a025c997c + 1;
                end else begin
                    I71c6f88cbabd48d41f42f2b16170c8955b79d20b8a8b211e174d1c1473567ad4  <= Idb5ffff327b8edefda5ee44436f5f31deac21a01781b65e2429b1e1a025c997c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00fca56df853315156adf3a6a5cdecaf6256b108f16f65b1e93272f0c7796e9c != I6020dcffd9e047c03740cffcdfe790eaf614ea1036a50fefcec9e13e5b5ac4bc[0] ) begin
                    Ib4c52550766a2cbe0de236d6783edfb1a6a7cb4c2bb9333a9379e1b75680dad1  <=  ~I0384038afb05788ee28f773a244ec49cd78da115f5d864f8497df2b36f37ae54 + 1;
                end else begin
                    Ib4c52550766a2cbe0de236d6783edfb1a6a7cb4c2bb9333a9379e1b75680dad1  <= I0384038afb05788ee28f773a244ec49cd78da115f5d864f8497df2b36f37ae54 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia6934e7e07061fec0575e9ceb1910150463d7c530d30091ee48fcc50bc2d0cf8 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[19] ) begin
                    I051f072f564eefd657cb4d59c1c851b56df2e70861d875f3b4c9b95e8945db08  <=  ~Ibee29fffd6b844b0fc4666fbb35c295ccc5a7b99dbedce125b370508cf6b0b90 + 1;
                end else begin
                    I051f072f564eefd657cb4d59c1c851b56df2e70861d875f3b4c9b95e8945db08  <= Ibee29fffd6b844b0fc4666fbb35c295ccc5a7b99dbedce125b370508cf6b0b90 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia6934e7e07061fec0575e9ceb1910150463d7c530d30091ee48fcc50bc2d0cf8 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[8] ) begin
                    Ia6f2e4979fa9229a647a81a4fa3f8b2af809199049d2554ea15fa9a6ba2f90a9  <=  ~Ia8f9f47f8cf0ac244089271b1cb952cac9d90aa94b91eef48733afbbcd992952 + 1;
                end else begin
                    Ia6f2e4979fa9229a647a81a4fa3f8b2af809199049d2554ea15fa9a6ba2f90a9  <= Ia8f9f47f8cf0ac244089271b1cb952cac9d90aa94b91eef48733afbbcd992952 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia6934e7e07061fec0575e9ceb1910150463d7c530d30091ee48fcc50bc2d0cf8 != I815f772d86db329f78fa75c3326c129ccf0f6c5f383b42ef18033e48d11525d2[0] ) begin
                    Iaa72101e8c3e7fa248ac4d4336b3847c4f602b6db009e9cd74cdd25251d5178e  <=  ~Ie80058ecf96cf544095e34ccc9662fb679b8da3cf6f10797805cbcaddfd63804 + 1;
                end else begin
                    Iaa72101e8c3e7fa248ac4d4336b3847c4f602b6db009e9cd74cdd25251d5178e  <= Ie80058ecf96cf544095e34ccc9662fb679b8da3cf6f10797805cbcaddfd63804 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8358c4f85a5a177702d111cdd3e705172bedf92a6d01f2c5d25b5e33c75538d != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[19] ) begin
                    Ifb6bf654293ed3bacd2a4ffc883b8ca5e4dedea39e338bd1a30b21e8f8df2f62  <=  ~I680b7384eb5b44faf98980956603d7db164a819fe394beff4e94872edcbece0b + 1;
                end else begin
                    Ifb6bf654293ed3bacd2a4ffc883b8ca5e4dedea39e338bd1a30b21e8f8df2f62  <= I680b7384eb5b44faf98980956603d7db164a819fe394beff4e94872edcbece0b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8358c4f85a5a177702d111cdd3e705172bedf92a6d01f2c5d25b5e33c75538d != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[8] ) begin
                    I01c264f9a89aec9dc11fa16206ffee1c8fb03bcb279e9e9f53fea1e94e9d8b23  <=  ~I7bdb6b57635075a7bb8408a878d4ef7f2ff136804287cfbacddb40bb20dd053a + 1;
                end else begin
                    I01c264f9a89aec9dc11fa16206ffee1c8fb03bcb279e9e9f53fea1e94e9d8b23  <= I7bdb6b57635075a7bb8408a878d4ef7f2ff136804287cfbacddb40bb20dd053a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8358c4f85a5a177702d111cdd3e705172bedf92a6d01f2c5d25b5e33c75538d != I2c8a33831a21c4c21dd58a300467abcc82d52e7636a73a12a003a4144d43e0dc[0] ) begin
                    Ic1381219782d18c1cb880970c062eb260d9d3be0b597e1465fc604c0c0c32c68  <=  ~I27f0b66e246c474ca71e1ae20503843b31921b5552092c5ae6eb872e76808395 + 1;
                end else begin
                    Ic1381219782d18c1cb880970c062eb260d9d3be0b597e1465fc604c0c0c32c68  <= I27f0b66e246c474ca71e1ae20503843b31921b5552092c5ae6eb872e76808395 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2e37b13b583174f0ca14a3fff3bbdd50d584c2a917a020de586b559bb7df4c45 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[19] ) begin
                    I6c3a9695a1c1d22809b1378e82cbdbebc1ca78428194df50cce0a69d6a159398  <=  ~Id81f3fed6908e777951bdff6448776a9a80348c44058ba0f9450999a26f6155f + 1;
                end else begin
                    I6c3a9695a1c1d22809b1378e82cbdbebc1ca78428194df50cce0a69d6a159398  <= Id81f3fed6908e777951bdff6448776a9a80348c44058ba0f9450999a26f6155f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2e37b13b583174f0ca14a3fff3bbdd50d584c2a917a020de586b559bb7df4c45 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[8] ) begin
                    I12dfae8d4c1a0612c6d65c6f5493247af5e06ca1d8c72dc28f9ca41b0bbc6ea3  <=  ~Ie4655a76ed253aad70f2340070cd7b6f2041e6782a87be16ea66ee0fa2e2ad74 + 1;
                end else begin
                    I12dfae8d4c1a0612c6d65c6f5493247af5e06ca1d8c72dc28f9ca41b0bbc6ea3  <= Ie4655a76ed253aad70f2340070cd7b6f2041e6782a87be16ea66ee0fa2e2ad74 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I2e37b13b583174f0ca14a3fff3bbdd50d584c2a917a020de586b559bb7df4c45 != I8c7b9ead4ab28ae2c2aa5185a0746c9cfe9fd90bdd68f2ba05291045a296d566[0] ) begin
                    Icf0c3c82c9e458a347212415d3029f192c40152e8525a20b5c9bfed88ccdb32e  <=  ~I8acc445f4b9f01af1a8f4f34ab10028472b79a2c1d1d3b8aed7d040f5ff4cff9 + 1;
                end else begin
                    Icf0c3c82c9e458a347212415d3029f192c40152e8525a20b5c9bfed88ccdb32e  <= I8acc445f4b9f01af1a8f4f34ab10028472b79a2c1d1d3b8aed7d040f5ff4cff9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[18] ) begin
                    I0e9135a0817e96971dc8c4fe6eec717a563c44738f7e38d5bfb2f4dda8c77876  <=  ~I11f1c07733856926d4d980234959cd48f8b0247270d6485cc57dc3456ba7adbf + 1;
                end else begin
                    I0e9135a0817e96971dc8c4fe6eec717a563c44738f7e38d5bfb2f4dda8c77876  <= I11f1c07733856926d4d980234959cd48f8b0247270d6485cc57dc3456ba7adbf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[10] ) begin
                    Id4cd4fdc9fdb1198c2894543e212f665c925298f1c92b4da9c432eca9442963d  <=  ~I26f2f2938065d9336a83a2edcb5595f6976c5c434c76d4c44e771cb8a0c685c4 + 1;
                end else begin
                    Id4cd4fdc9fdb1198c2894543e212f665c925298f1c92b4da9c432eca9442963d  <= I26f2f2938065d9336a83a2edcb5595f6976c5c434c76d4c44e771cb8a0c685c4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[6] ) begin
                    Ibc34c6979b8f5adc5421ca8603b6dca91161055286758ac10d0c612263077758  <=  ~I059b4a33ad6774feb79158ff05ecb4287420d94dc0c57650fb90f11fb7fb83ec + 1;
                end else begin
                    Ibc34c6979b8f5adc5421ca8603b6dca91161055286758ac10d0c612263077758  <= I059b4a33ad6774feb79158ff05ecb4287420d94dc0c57650fb90f11fb7fb83ec ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8 != I32ed4ecd4363760151c1accda085c9afa3efe63daf7a312feefc00b804401c27[0] ) begin
                    Ic5a87abf4c6018e9555de321c141d9754a7de91f1743d980e339ff9cebd63b7a  <=  ~I9a9e162c226e402630bd217ff502dc5aa823ee7c089801803c5ee091b5ea4026 + 1;
                end else begin
                    Ic5a87abf4c6018e9555de321c141d9754a7de91f1743d980e339ff9cebd63b7a  <= I9a9e162c226e402630bd217ff502dc5aa823ee7c089801803c5ee091b5ea4026 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[18] ) begin
                    Ie38c638da580ca7d25fc0754497163d0369f31a6cdb4bd26663a759b74efd588  <=  ~If30f29822c81c32a3f153165fbdd82ff6cd9527a6a065627852ca8d5d1a0b122 + 1;
                end else begin
                    Ie38c638da580ca7d25fc0754497163d0369f31a6cdb4bd26663a759b74efd588  <= If30f29822c81c32a3f153165fbdd82ff6cd9527a6a065627852ca8d5d1a0b122 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[10] ) begin
                    Id8d0e36ce1faa76feb8cbe0331f2179ddfc066b70e93e990b5d5bce17f505440  <=  ~Iec9d3d3ad44a5c22fbedf1fc73a01cf348f8c4b16c5f3f0cf55c85f8d92ca22b + 1;
                end else begin
                    Id8d0e36ce1faa76feb8cbe0331f2179ddfc066b70e93e990b5d5bce17f505440  <= Iec9d3d3ad44a5c22fbedf1fc73a01cf348f8c4b16c5f3f0cf55c85f8d92ca22b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601 != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[6] ) begin
                    Icf55933dce8b9f95a57d7d019c9b29f72e08454428013009cf0e4d2c5b6edf0b  <=  ~I94452304db6f03a077cc46cd087cc756c098f85885a9c8a60e1860ebb0b23a60 + 1;
                end else begin
                    Icf55933dce8b9f95a57d7d019c9b29f72e08454428013009cf0e4d2c5b6edf0b  <= I94452304db6f03a077cc46cd087cc756c098f85885a9c8a60e1860ebb0b23a60 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601 != I6aa6d6c6213348ea0cc3e8b207bca2c1db81499441e4ed721ca0ee01ae831291[0] ) begin
                    I3a27e4e3322c28e7fe85d7e76b7d5477f4d4f6acb8cdb876b9a54cba98b189b9  <=  ~I59d79bf88b865cc38882adc0e8d69f2a1556f9cef906cd558730ea7a902de6ce + 1;
                end else begin
                    I3a27e4e3322c28e7fe85d7e76b7d5477f4d4f6acb8cdb876b9a54cba98b189b9  <= I59d79bf88b865cc38882adc0e8d69f2a1556f9cef906cd558730ea7a902de6ce ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[18] ) begin
                    I099e314496f03784e5504a35292defa79dc063aa81e6aa8764802f7fe3a47114  <=  ~I022500b8d9cd3b589fb75b90c1b633a96fdc76c0e3e2ec514cf7b4ff3ccce1b6 + 1;
                end else begin
                    I099e314496f03784e5504a35292defa79dc063aa81e6aa8764802f7fe3a47114  <= I022500b8d9cd3b589fb75b90c1b633a96fdc76c0e3e2ec514cf7b4ff3ccce1b6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[10] ) begin
                    I9d7506b5ed3de0e32e821ce6ddd1c28aed177910ccacc4d4aa2a8ee57212d162  <=  ~Id9936f1014242296259237c4aa19452ea56509e2d970ce60c72e7c4d18a66752 + 1;
                end else begin
                    I9d7506b5ed3de0e32e821ce6ddd1c28aed177910ccacc4d4aa2a8ee57212d162  <= Id9936f1014242296259237c4aa19452ea56509e2d970ce60c72e7c4d18a66752 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[6] ) begin
                    I525b9b85b14df7a6533a7e54bdc9bf40a303c890a4a410251c8d556d38b33125  <=  ~Idad105c150f27de4777164385ed4e2123966f63d2b2ff32add6d18a95be2624d + 1;
                end else begin
                    I525b9b85b14df7a6533a7e54bdc9bf40a303c890a4a410251c8d556d38b33125  <= Idad105c150f27de4777164385ed4e2123966f63d2b2ff32add6d18a95be2624d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f != Ib4f23d2e5f8c73110ae24212c4ec0e7ef29c09c8178ec3850f061a5b0386feca[0] ) begin
                    I11edfeb948852dab396975b53b12d09da7a5fbedc2dae9fe7c687768cfef05b4  <=  ~Ice1023bfed1f964ccc66c7d914378cc899ac310a76f3d694302cc688bb560e45 + 1;
                end else begin
                    I11edfeb948852dab396975b53b12d09da7a5fbedc2dae9fe7c687768cfef05b4  <= Ice1023bfed1f964ccc66c7d914378cc899ac310a76f3d694302cc688bb560e45 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[18] ) begin
                    Ifa0b8243f5ab6adb88a70fc1245e3480ea3fb3f3af846fdefd0613ca91d7b122  <=  ~I372b0e45c0d1e8d30830bd3cac2c3082ec36f9af195380d0e1b7d62712123fa7 + 1;
                end else begin
                    Ifa0b8243f5ab6adb88a70fc1245e3480ea3fb3f3af846fdefd0613ca91d7b122  <= I372b0e45c0d1e8d30830bd3cac2c3082ec36f9af195380d0e1b7d62712123fa7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[10] ) begin
                    I1bfa3da571b0e3d943ec7b9a8c641283e080bcc6502fa8317ced3c0a6eb2c4cf  <=  ~Ie98369c31ad7be164b6fc0f16fd6d1a5193f2b00a3eb10ee1cb478b4653b60fe + 1;
                end else begin
                    I1bfa3da571b0e3d943ec7b9a8c641283e080bcc6502fa8317ced3c0a6eb2c4cf  <= Ie98369c31ad7be164b6fc0f16fd6d1a5193f2b00a3eb10ee1cb478b4653b60fe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6 != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[6] ) begin
                    I2ade6ee1b52da04fce9491cad314947a07eb9aaa8b0a430db2f96e2d290384dc  <=  ~I80f30106eccbcdd1f0aabed1521d2b09a4bb56a421079ec90f81527a903c6643 + 1;
                end else begin
                    I2ade6ee1b52da04fce9491cad314947a07eb9aaa8b0a430db2f96e2d290384dc  <= I80f30106eccbcdd1f0aabed1521d2b09a4bb56a421079ec90f81527a903c6643 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6 != If2be986b27ce8aa2117f87e9a144015a10acf0a07847f83acec2804b9e987e8b[0] ) begin
                    I578437932d2d1156445b41a1238e0fd96ab5702bc3158ea337a9e37d14d6731e  <=  ~I81349ebf72720f77a8902dc12d9cf986ddec6f8fe30f7f76f9f4dc54881708b5 + 1;
                end else begin
                    I578437932d2d1156445b41a1238e0fd96ab5702bc3158ea337a9e37d14d6731e  <= I81349ebf72720f77a8902dc12d9cf986ddec6f8fe30f7f76f9f4dc54881708b5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[7] ) begin
                    I8411087f9f6fa41d454a74dc89e5152e5e8edfa501c8753bd0735cec3789f14b  <=  ~Ic941f62ac4a004ce3dfdcdfc5312a3be16a5307024d1ad292754532cec3fc90b + 1;
                end else begin
                    I8411087f9f6fa41d454a74dc89e5152e5e8edfa501c8753bd0735cec3789f14b  <= Ic941f62ac4a004ce3dfdcdfc5312a3be16a5307024d1ad292754532cec3fc90b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[10] ) begin
                    I11775c069ab4acd951a3ca47bfa65c7632a6a8a369bb103d0bb719806dfe0c57  <=  ~I65c4ade7c4c23e62f5cd1846b0a739c70cd498087298f54c41f89bbd9677e705 + 1;
                end else begin
                    I11775c069ab4acd951a3ca47bfa65c7632a6a8a369bb103d0bb719806dfe0c57  <= I65c4ade7c4c23e62f5cd1846b0a739c70cd498087298f54c41f89bbd9677e705 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[6] ) begin
                    I6a2505f0de03f3e2d303fd207ee819f5a1777b650930b87a235ab3cca5de6e87  <=  ~I4d548bf4a643564a906a42a32acc4fe6919c91f43890f1b921b9e42100b92e68 + 1;
                end else begin
                    I6a2505f0de03f3e2d303fd207ee819f5a1777b650930b87a235ab3cca5de6e87  <= I4d548bf4a643564a906a42a32acc4fe6919c91f43890f1b921b9e42100b92e68 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9 != I9f17331c6a9858b60705d889b5b77078042cffe9e956de20eb067ad7e70626b7[0] ) begin
                    I3c2c5b5cd798851c7fcb0d0e66ddf81a516ef9bdf4aa4ebd4901532bfb2a651b  <=  ~Id89fd01703e5a1c53c89a64885698fdf565b791620408fb963b53208a33e7f47 + 1;
                end else begin
                    I3c2c5b5cd798851c7fcb0d0e66ddf81a516ef9bdf4aa4ebd4901532bfb2a651b  <= Id89fd01703e5a1c53c89a64885698fdf565b791620408fb963b53208a33e7f47 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26 != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[7] ) begin
                    Iae213c2ac7729f8efe23deca256bf56f030403ef6ac00a3bc181414b6a3aa75e  <=  ~I8467f29aa6da06588468e21697c56464c67e4809c135d2d41e38d9881715aee7 + 1;
                end else begin
                    Iae213c2ac7729f8efe23deca256bf56f030403ef6ac00a3bc181414b6a3aa75e  <= I8467f29aa6da06588468e21697c56464c67e4809c135d2d41e38d9881715aee7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[10] ) begin
                    I2985f4f17b726f40ab6609b57a796727fe46605944c5e25c594caa8dfbea9f58  <=  ~I55ee374c21e5aee6b0ada78409b18bdefed20abbf3dc5716c62daa87b418dcfa + 1;
                end else begin
                    I2985f4f17b726f40ab6609b57a796727fe46605944c5e25c594caa8dfbea9f58  <= I55ee374c21e5aee6b0ada78409b18bdefed20abbf3dc5716c62daa87b418dcfa ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26 != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[6] ) begin
                    I1b0f11f3bca53713a53e2ed18fb81f5a25c7151c874be612677f5204bca28093  <=  ~I4285be4ac50db4da7f720fe115c342ad8ecefdf6dbace4af4c9714009ae31e86 + 1;
                end else begin
                    I1b0f11f3bca53713a53e2ed18fb81f5a25c7151c874be612677f5204bca28093  <= I4285be4ac50db4da7f720fe115c342ad8ecefdf6dbace4af4c9714009ae31e86 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26 != I2b70416e96231188e62b7bcf0300c4a5b2d2139449150d31414b92ae075aa0e7[0] ) begin
                    I8153d6f17d832da24daaba2909a88f1609e523ad3b6eac7ad42521979aae96da  <=  ~If37e3544f587a047696dc53e30f6031f848e27a13e2328b2c38a4f51421954db + 1;
                end else begin
                    I8153d6f17d832da24daaba2909a88f1609e523ad3b6eac7ad42521979aae96da  <= If37e3544f587a047696dc53e30f6031f848e27a13e2328b2c38a4f51421954db ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[7] ) begin
                    I4c0096e7bbf30db97520f824e05dbc28e6d1db344202349993fc68cbc95d6585  <=  ~Id9067d2f353cbef30dc828f16a97436418af2bf3e5fd19300471de394f710fff + 1;
                end else begin
                    I4c0096e7bbf30db97520f824e05dbc28e6d1db344202349993fc68cbc95d6585  <= Id9067d2f353cbef30dc828f16a97436418af2bf3e5fd19300471de394f710fff ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[10] ) begin
                    I73ecf8ab6430c6343bf7596e671ce01a3e3e7499813ed75c583a7103147b0bb7  <=  ~I93150066a1cfdd9e59edd1d42cd2611eac0df4fdfbea33d913804f52dbd895a5 + 1;
                end else begin
                    I73ecf8ab6430c6343bf7596e671ce01a3e3e7499813ed75c583a7103147b0bb7  <= I93150066a1cfdd9e59edd1d42cd2611eac0df4fdfbea33d913804f52dbd895a5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67 != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[6] ) begin
                    Iea7b69c43ca4b3707d3bfddf19b27616b8686df915734ba86d3685127bfbf39a  <=  ~Ie296c1317a499d9d35191ae9de6c681e2b521a2966b8837ffa470e3de6c8530d + 1;
                end else begin
                    Iea7b69c43ca4b3707d3bfddf19b27616b8686df915734ba86d3685127bfbf39a  <= Ie296c1317a499d9d35191ae9de6c681e2b521a2966b8837ffa470e3de6c8530d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67 != I29599a1dac362c87f4780a94478787a718f63401d2051ccbfe543b44e49b35bb[0] ) begin
                    Ic10ea001dcd0b864b987bc3080e95b338c1e91247bb90e884e161c926183fd2b  <=  ~I0aecd8795e3571b4b428903758f7dac78966a9a928f64c26a3e6f00fd61872ab + 1;
                end else begin
                    Ic10ea001dcd0b864b987bc3080e95b338c1e91247bb90e884e161c926183fd2b  <= I0aecd8795e3571b4b428903758f7dac78966a9a928f64c26a3e6f00fd61872ab ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[7] ) begin
                    If692b993dc571ec401ce86f38a18ea4f96a797b00c04699ce83ce875b7c31730  <=  ~I0bc6fa0d581c2d2fcce482d2821bf87f00bc84606afa8b56d7f4cd88bead4a3d + 1;
                end else begin
                    If692b993dc571ec401ce86f38a18ea4f96a797b00c04699ce83ce875b7c31730  <= I0bc6fa0d581c2d2fcce482d2821bf87f00bc84606afa8b56d7f4cd88bead4a3d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[10] ) begin
                    I5dfc39b913b8e0d00491e3f7f45b6b467a517b5e87baa065097e28e6d695500a  <=  ~Idfee0ad9592b445c7afa92c1099d49c458d1eda5605ad06e6ec975e2d9103e11 + 1;
                end else begin
                    I5dfc39b913b8e0d00491e3f7f45b6b467a517b5e87baa065097e28e6d695500a  <= Idfee0ad9592b445c7afa92c1099d49c458d1eda5605ad06e6ec975e2d9103e11 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[6] ) begin
                    I9ede22dbb56f48c045a1b5a05945124fb97b6ca7e355dd8d9dcfdef6e623b953  <=  ~Ic700c1c29d2fbb8e2e85fd9871082303e3dada09845afca88fd7c35f9d41affe + 1;
                end else begin
                    I9ede22dbb56f48c045a1b5a05945124fb97b6ca7e355dd8d9dcfdef6e623b953  <= Ic700c1c29d2fbb8e2e85fd9871082303e3dada09845afca88fd7c35f9d41affe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d != I5ff7defb023005e77164f9f3b852fa60ce897922c6b814015d3436fe1d1b4a44[0] ) begin
                    I61efe7187a1aaa28235dacf68eb1e1dd97e7cb5900862790bb4d5872d7adbd67  <=  ~Ie1342b74cd710b1a52ba3de5ca28ee42d03eaf53a42a6cedab9ecb6d987d7b55 + 1;
                end else begin
                    I61efe7187a1aaa28235dacf68eb1e1dd97e7cb5900862790bb4d5872d7adbd67  <= Ie1342b74cd710b1a52ba3de5ca28ee42d03eaf53a42a6cedab9ecb6d987d7b55 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[19] ) begin
                    I2c635a0b11af3be4774428af79ff5cbe6a32ede6ad03ac197ecbb3ca2ba78f8f  <=  ~I69f8afa3d9aea957a3c1a9f3dbfd8ef8dc6370b228a7f67f0a27113c094992ed + 1;
                end else begin
                    I2c635a0b11af3be4774428af79ff5cbe6a32ede6ad03ac197ecbb3ca2ba78f8f  <= I69f8afa3d9aea957a3c1a9f3dbfd8ef8dc6370b228a7f67f0a27113c094992ed ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[7] ) begin
                    If6e953221a61b86b1fc339b69af853f6ad538b60770f2f7b880d7aa15bd625b3  <=  ~I3b017b72afccffaac4ff923e52843d312e1cd5e1123575d6daf4692f81cfe748 + 1;
                end else begin
                    If6e953221a61b86b1fc339b69af853f6ad538b60770f2f7b880d7aa15bd625b3  <= I3b017b72afccffaac4ff923e52843d312e1cd5e1123575d6daf4692f81cfe748 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[9] ) begin
                    I295da244d8dab1563a5947230e49171eb905c3758c289526ff6d3e0c3efcebbb  <=  ~I100b4afda393740a5fcf563e8e5fe34d5d7bfc439f2eedd77966bc9b37b3d602 + 1;
                end else begin
                    I295da244d8dab1563a5947230e49171eb905c3758c289526ff6d3e0c3efcebbb  <= I100b4afda393740a5fcf563e8e5fe34d5d7bfc439f2eedd77966bc9b37b3d602 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d != Ie132a24e667376de85b8fff9a639698df164043422122a8058c968bb7996d3a7[0] ) begin
                    I3c710fbd5e4dce0c97eb9da2d8e526f9d44d87fa75088c0421353614e6ef5da9  <=  ~Ieeaf4fb83c3c92f18b21f65ff2a951f74693fa6da2ec322ae6a4873d26729f51 + 1;
                end else begin
                    I3c710fbd5e4dce0c97eb9da2d8e526f9d44d87fa75088c0421353614e6ef5da9  <= Ieeaf4fb83c3c92f18b21f65ff2a951f74693fa6da2ec322ae6a4873d26729f51 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[19] ) begin
                    Id4bcb557769f043a7275ab01d6d9794d4cbbd9309be38f58acc307a1e693f347  <=  ~I27ac039dc48350ce90d2a8a3953936d5f7c97ec1098fb20d853cd062f2d4a6f9 + 1;
                end else begin
                    Id4bcb557769f043a7275ab01d6d9794d4cbbd9309be38f58acc307a1e693f347  <= I27ac039dc48350ce90d2a8a3953936d5f7c97ec1098fb20d853cd062f2d4a6f9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[7] ) begin
                    Id39c55c4f0df8a0d8ee4f8b47f3de8cebf5343bf75521edfe38a695565eea926  <=  ~I224433de24984b12aa905ae86eeaa53ec459acd68fefdba7aa1e8778abb89408 + 1;
                end else begin
                    Id39c55c4f0df8a0d8ee4f8b47f3de8cebf5343bf75521edfe38a695565eea926  <= I224433de24984b12aa905ae86eeaa53ec459acd68fefdba7aa1e8778abb89408 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70 != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[9] ) begin
                    I1e7e130607ec849c80f9e687f0215ceb767a2650626f20ee44a6fe677fde2299  <=  ~Ice1b30668532ff63b6ead40f37366b805ea21a65f6fb7067bf9d3b5d08eced46 + 1;
                end else begin
                    I1e7e130607ec849c80f9e687f0215ceb767a2650626f20ee44a6fe677fde2299  <= Ice1b30668532ff63b6ead40f37366b805ea21a65f6fb7067bf9d3b5d08eced46 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70 != Ie8d5dfc9a77dc01055a551c5f37416d0b13ef83428bf751fb9f95c7d10442697[0] ) begin
                    Ie02f677979058dda2291ddb93acd64f4461f6d75f3a33c21dac97129344f7055  <=  ~I2b6551d9c8b14c787afa552e23234fdbb63c8fdb8fb285416ff1b72a38e7d898 + 1;
                end else begin
                    Ie02f677979058dda2291ddb93acd64f4461f6d75f3a33c21dac97129344f7055  <= I2b6551d9c8b14c787afa552e23234fdbb63c8fdb8fb285416ff1b72a38e7d898 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[19] ) begin
                    Ia00cd24df6e6b22b466e1492500f1948b3ba3d70bdca407d1c22b4dfaf374eb7  <=  ~I24ade58e2190b73f141a858e6812d93a49203181d6d427a29415d014a9cceec6 + 1;
                end else begin
                    Ia00cd24df6e6b22b466e1492500f1948b3ba3d70bdca407d1c22b4dfaf374eb7  <= I24ade58e2190b73f141a858e6812d93a49203181d6d427a29415d014a9cceec6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[7] ) begin
                    I5b0da0701e7399ca2e668c1602f494f41127e4c90e6fa91632da0016e7b395e9  <=  ~I55affee832ae4e480ffb916ce8a5e3b12fb6429f1ccee3a8f9a668aeb8352f7e + 1;
                end else begin
                    I5b0da0701e7399ca2e668c1602f494f41127e4c90e6fa91632da0016e7b395e9  <= I55affee832ae4e480ffb916ce8a5e3b12fb6429f1ccee3a8f9a668aeb8352f7e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[9] ) begin
                    I83d70d4886f48dce0888e203c2c333c76d35f0c73767dd9443ec8fa4790ecb09  <=  ~I3f2f052f1d132cf1a83172a044968741665a7b85e421658976109057a3d00ba1 + 1;
                end else begin
                    I83d70d4886f48dce0888e203c2c333c76d35f0c73767dd9443ec8fa4790ecb09  <= I3f2f052f1d132cf1a83172a044968741665a7b85e421658976109057a3d00ba1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d != Ic94f2b10208cb23bb5f5b1a46c11c3bbae038308b385373cfaad9a18e09ccb90[0] ) begin
                    I2b78100b50f7334d563daa27cab8078fa374dca0c438157d1ad44ed3fd9e3456  <=  ~Ibbe3cd91dfae5930a6ae5799a27b045ce6e0c59fe00a38b5fb4b1691949847f2 + 1;
                end else begin
                    I2b78100b50f7334d563daa27cab8078fa374dca0c438157d1ad44ed3fd9e3456  <= Ibbe3cd91dfae5930a6ae5799a27b045ce6e0c59fe00a38b5fb4b1691949847f2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[19] ) begin
                    I0847713503570d7ab3efee12577ba27aa81869a22b14ec8a244fbd4665d566f4  <=  ~Icbbfd81a7f066da629076f9f7c26eb457be34298a6518cf45e67bb39e74f5f2a + 1;
                end else begin
                    I0847713503570d7ab3efee12577ba27aa81869a22b14ec8a244fbd4665d566f4  <= Icbbfd81a7f066da629076f9f7c26eb457be34298a6518cf45e67bb39e74f5f2a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[7] ) begin
                    I65afc937c55081dabf16dbfd02eb03c97204efbdcfbb523609571bb32d537d5e  <=  ~I762a7e10d310500a1080b7b46a9a30bb003c7a7d48011e96501a647e1de0cb66 + 1;
                end else begin
                    I65afc937c55081dabf16dbfd02eb03c97204efbdcfbb523609571bb32d537d5e  <= I762a7e10d310500a1080b7b46a9a30bb003c7a7d48011e96501a647e1de0cb66 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[9] ) begin
                    Ie42f89c20abd223240a9f93a89ce650ed2f581e1ceab0587a4fea2ddf9f4f98f  <=  ~Idc9ce24f8fd9ca7372ef25d9e2b8414a4c8051c796f9ce64b91a6f3e70faeec6 + 1;
                end else begin
                    Ie42f89c20abd223240a9f93a89ce650ed2f581e1ceab0587a4fea2ddf9f4f98f  <= Idc9ce24f8fd9ca7372ef25d9e2b8414a4c8051c796f9ce64b91a6f3e70faeec6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf != I3b79a6c69be124aeea9d1444f9f985201b55ad0d7a4767a01f612eee12a6ad73[0] ) begin
                    Icdfa68bdad11213dbaa576cbf43ca9deeb1f9f24225264eaeeede7d1aba5fd8a  <=  ~Iffe887b6857424a57f7b7bec156197556dd869c44a2eaa660fa66760cd88888a + 1;
                end else begin
                    Icdfa68bdad11213dbaa576cbf43ca9deeb1f9f24225264eaeeede7d1aba5fd8a  <= Iffe887b6857424a57f7b7bec156197556dd869c44a2eaa660fa66760cd88888a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[20] ) begin
                    I4d032ff7482be75de7d2b816ddb2bebfa9e896e45fdade2b5f81b35c003a59ac  <=  ~Ie7328907da6b377ef494c54a5e6fc2f90992a99258967af4bc2205d0d42e9db1 + 1;
                end else begin
                    I4d032ff7482be75de7d2b816ddb2bebfa9e896e45fdade2b5f81b35c003a59ac  <= Ie7328907da6b377ef494c54a5e6fc2f90992a99258967af4bc2205d0d42e9db1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[11] ) begin
                    I2e15c5739b990462c8a17b590fb7d60ac9c7e6648b79e75697139f55221fbcc5  <=  ~I98616ac468624d04fcf2487684bc23bd20a87b719be4d4533f987ecb1bcc8d5c + 1;
                end else begin
                    I2e15c5739b990462c8a17b590fb7d60ac9c7e6648b79e75697139f55221fbcc5  <= I98616ac468624d04fcf2487684bc23bd20a87b719be4d4533f987ecb1bcc8d5c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[13] ) begin
                    I717aab2686adb8a0688009c23d92aa4475e240ec0747735e6fee5e196a50c444  <=  ~Ieb0d5850e57aa2cd83ee69ba71c85e9e047a9cc5b195da367a9f042a39559f47 + 1;
                end else begin
                    I717aab2686adb8a0688009c23d92aa4475e240ec0747735e6fee5e196a50c444  <= Ieb0d5850e57aa2cd83ee69ba71c85e9e047a9cc5b195da367a9f042a39559f47 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb != Id3ac4bf805d3981ac1eb1b396b3da5c0dbc68754d89668f0a4cf7c6f2a44ddfa[0] ) begin
                    Idb39db95234cbfdbbc89fdee230784c703e170b9e932643a5e1b811b24ae021a  <=  ~If6bf4d8f739928e726bca59f6307a2b78966853a5aeae6bb7dc4786660382ad9 + 1;
                end else begin
                    Idb39db95234cbfdbbc89fdee230784c703e170b9e932643a5e1b811b24ae021a  <= If6bf4d8f739928e726bca59f6307a2b78966853a5aeae6bb7dc4786660382ad9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[20] ) begin
                    I448065f71638c5abddd1eba1fcf567566281d5b4b23ec4ff2d2208d32a506fbf  <=  ~I3fc232b4e4ad45bd25aaed0b1306112944d63174fc4f473899349954e94895cd + 1;
                end else begin
                    I448065f71638c5abddd1eba1fcf567566281d5b4b23ec4ff2d2208d32a506fbf  <= I3fc232b4e4ad45bd25aaed0b1306112944d63174fc4f473899349954e94895cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[11] ) begin
                    Iaef8ec1714d2faf3d3b947db31b7975161077ca31fee04842efc1f7159104d30  <=  ~I07c430087a2a880f756db41ba39cef794ad6d3b28723a7c22df5aa719bf585c2 + 1;
                end else begin
                    Iaef8ec1714d2faf3d3b947db31b7975161077ca31fee04842efc1f7159104d30  <= I07c430087a2a880f756db41ba39cef794ad6d3b28723a7c22df5aa719bf585c2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[13] ) begin
                    I58d2fcb7085fddc9250ca075b010afdc2d019c4091f5d115d9520586224a1ae8  <=  ~Iff963f656b33e8c5d0b4155f3d4ce0be5ec1c056727223d45af4ae070b006272 + 1;
                end else begin
                    I58d2fcb7085fddc9250ca075b010afdc2d019c4091f5d115d9520586224a1ae8  <= Iff963f656b33e8c5d0b4155f3d4ce0be5ec1c056727223d45af4ae070b006272 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02 != Id77fd99c6146776bfc20804c67ae41b88cb0441eecba4f40b87828956b7158b6[0] ) begin
                    I7141b42fce475b5502fd33035bf37addde06271b2259e158ba03a66843b66075  <=  ~I44d78165b52487e966d2063495d2b76b8086031f3d3f0bac7713717f1e56b721 + 1;
                end else begin
                    I7141b42fce475b5502fd33035bf37addde06271b2259e158ba03a66843b66075  <= I44d78165b52487e966d2063495d2b76b8086031f3d3f0bac7713717f1e56b721 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[20] ) begin
                    Ifc8302f040679d23faab1ed8387a8a3aec85aba86ba9a78d3ca903126266af4e  <=  ~I6e5de0450866fddb6d15781d26a3df126ea57faea36d172ff9c08fbed711ea47 + 1;
                end else begin
                    Ifc8302f040679d23faab1ed8387a8a3aec85aba86ba9a78d3ca903126266af4e  <= I6e5de0450866fddb6d15781d26a3df126ea57faea36d172ff9c08fbed711ea47 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[11] ) begin
                    I734136c95a40c62745d684fc7e8cd1114b883c6209df11cfe01b9174cffc720a  <=  ~Ie4db811b4d839e478783694d956589c702666e122689ec06c5fcd299c782b1a7 + 1;
                end else begin
                    I734136c95a40c62745d684fc7e8cd1114b883c6209df11cfe01b9174cffc720a  <= Ie4db811b4d839e478783694d956589c702666e122689ec06c5fcd299c782b1a7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8 != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[13] ) begin
                    If4fa37977e1db59d1bd7a30b2b0919c997b6e25e0438e01b62dc273d10497867  <=  ~I23072d2753b8750a9cd8da42f6ec9fdce24f0ccf4c201e983c3aa96963421ed3 + 1;
                end else begin
                    If4fa37977e1db59d1bd7a30b2b0919c997b6e25e0438e01b62dc273d10497867  <= I23072d2753b8750a9cd8da42f6ec9fdce24f0ccf4c201e983c3aa96963421ed3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8 != I650a7220fd4eb743f652c6c1f9431191621f9fb1a5b5d64bb9649b43bad5b8bf[0] ) begin
                    I245e922da0aa5470370db389d5bc9db33327c905528a1740aa015b7ccdfcc29e  <=  ~I96d2ff73be5717714513ef2406648446833f53abe34481e91be763d63d3f2d09 + 1;
                end else begin
                    I245e922da0aa5470370db389d5bc9db33327c905528a1740aa015b7ccdfcc29e  <= I96d2ff73be5717714513ef2406648446833f53abe34481e91be763d63d3f2d09 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436 != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[20] ) begin
                    I0f4ede6017039c42f04051822cfc539cbcacd77427efe92d393ade1c10a46462  <=  ~If7d7e9843a2eed7a0478c5991a13e140b1ab83460cc8ea6a3bf24a85b8d8ae49 + 1;
                end else begin
                    I0f4ede6017039c42f04051822cfc539cbcacd77427efe92d393ade1c10a46462  <= If7d7e9843a2eed7a0478c5991a13e140b1ab83460cc8ea6a3bf24a85b8d8ae49 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[11] ) begin
                    Idfa7c6c8248be1a2f8a95c6c74a71be3126e039a31f4e16e0b964476c6d47953  <=  ~I61ea75f5f583a43e3691ab2462210c213f53492dd6a4a0a41abc406a7a828bd8 + 1;
                end else begin
                    Idfa7c6c8248be1a2f8a95c6c74a71be3126e039a31f4e16e0b964476c6d47953  <= I61ea75f5f583a43e3691ab2462210c213f53492dd6a4a0a41abc406a7a828bd8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[13] ) begin
                    I0568efb50e0bb85c39c9ac6d2ab3474ab38799257dac5693085eeb0d74859ade  <=  ~I2668038e4b55b5d2fbdfcb8fdc56d43beaf4546ba92b39940b8f055a51d7013f + 1;
                end else begin
                    I0568efb50e0bb85c39c9ac6d2ab3474ab38799257dac5693085eeb0d74859ade  <= I2668038e4b55b5d2fbdfcb8fdc56d43beaf4546ba92b39940b8f055a51d7013f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436 != Ib7417e90e9dc35367f110c364878657dbbf66b1a714d5807e6347095b833c62d[0] ) begin
                    Ia2ff4d61c4f4fdf29be87b50e206c308cf970cbad2638e86ba8c2be8d025b534  <=  ~Ia29b333453d0a00fb718748060cc9eb198035cf24697fefdcc6b75b450e5fa6c + 1;
                end else begin
                    Ia2ff4d61c4f4fdf29be87b50e206c308cf970cbad2638e86ba8c2be8d025b534  <= Ia29b333453d0a00fb718748060cc9eb198035cf24697fefdcc6b75b450e5fa6c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[20] ) begin
                    Id1bb830ea0f92a1c0ed0addc915fc85198e4744c4bf7369b4ee1f7131f5f8542  <=  ~I9c17b85d3c4d97f0a7093e8007d812455859adb691cd79d2e41e78f95c44d2d4 + 1;
                end else begin
                    Id1bb830ea0f92a1c0ed0addc915fc85198e4744c4bf7369b4ee1f7131f5f8542  <= I9c17b85d3c4d97f0a7093e8007d812455859adb691cd79d2e41e78f95c44d2d4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[8] ) begin
                    I75c796f56576dfba821e867b0de1a871ef35851371c3aa422532bd287f02ee11  <=  ~Idb9949cbe1d38f86e61e1cce9211aa264e0abfb2ea1afa05be251144a4a081b1 + 1;
                end else begin
                    I75c796f56576dfba821e867b0de1a871ef35851371c3aa422532bd287f02ee11  <= Idb9949cbe1d38f86e61e1cce9211aa264e0abfb2ea1afa05be251144a4a081b1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2 != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[11] ) begin
                    Ib7f659da098e577e33fc0f5da1c03f6d3e68b3883ad7888152d2e8684a6177f3  <=  ~I18216dc1eb7be60021a2be1d64303e6b9838aaaa2a9b1e6bdffd2a3789661432 + 1;
                end else begin
                    Ib7f659da098e577e33fc0f5da1c03f6d3e68b3883ad7888152d2e8684a6177f3  <= I18216dc1eb7be60021a2be1d64303e6b9838aaaa2a9b1e6bdffd2a3789661432 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2 != Ie59a4afbd0d65de2149e8c60229bce12b77f8f1b2b232a11fb9714371eced2b9[0] ) begin
                    Idd383630385363471e1b17ea946a61194a3cb287d833af386876c3b4ee66e406  <=  ~Id8f0e532c3fc4af615d6cf0967f8a54e6971c1f3572b4383c25360f5f8204ac3 + 1;
                end else begin
                    Idd383630385363471e1b17ea946a61194a3cb287d833af386876c3b4ee66e406  <= Id8f0e532c3fc4af615d6cf0967f8a54e6971c1f3572b4383c25360f5f8204ac3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431 != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[20] ) begin
                    I8b41f817a4008df0994e2efa6b33eb847e82b031082f90a767467ffc03cfdb93  <=  ~Ia59883b6b96f3bbe38c2326bfca00e25d3b596e7ddf9287bbf70107666855849 + 1;
                end else begin
                    I8b41f817a4008df0994e2efa6b33eb847e82b031082f90a767467ffc03cfdb93  <= Ia59883b6b96f3bbe38c2326bfca00e25d3b596e7ddf9287bbf70107666855849 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431 != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[8] ) begin
                    Id5a74d0be90678a7b69691c10e4ab75b47914e213e67eae2f20d4b58e8a8d9ac  <=  ~Ied4edbf18ed0371b7d1ffd53ca5d98f1344d1640b4ca9733d97af5ba5c1c2a5a + 1;
                end else begin
                    Id5a74d0be90678a7b69691c10e4ab75b47914e213e67eae2f20d4b58e8a8d9ac  <= Ied4edbf18ed0371b7d1ffd53ca5d98f1344d1640b4ca9733d97af5ba5c1c2a5a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[11] ) begin
                    Ie538f6d2c778992e2324a9adbde215acaf7b8dc3a72a9230d4fba2332f3cab67  <=  ~If9a4d7f44a518a3ab1ecc6bd5d4e05d8e8f78615ebada754f1ef1e7b13a0e956 + 1;
                end else begin
                    Ie538f6d2c778992e2324a9adbde215acaf7b8dc3a72a9230d4fba2332f3cab67  <= If9a4d7f44a518a3ab1ecc6bd5d4e05d8e8f78615ebada754f1ef1e7b13a0e956 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431 != Iad3f7ae48f752d3ee71320875a2d1d170e879dd5ff51cdfd662241e6a30fca6d[0] ) begin
                    I3daa8702e9dbd047a05e5ea044d14b670c2ae3849526cc514be6a511c5c45c35  <=  ~I53fa59c42044794f03f617ff512486e58e173121f75b8dc3eb292e9246f7740f + 1;
                end else begin
                    I3daa8702e9dbd047a05e5ea044d14b670c2ae3849526cc514be6a511c5c45c35  <= I53fa59c42044794f03f617ff512486e58e173121f75b8dc3eb292e9246f7740f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[20] ) begin
                    I7b529f16d1499766369f75cde5a356cb12c06d21f42a10932edc6d54146735a0  <=  ~I9ae27a7b654a36e4265449d861213978965e4cc3bc7f36b77c6a77cde5e24f77 + 1;
                end else begin
                    I7b529f16d1499766369f75cde5a356cb12c06d21f42a10932edc6d54146735a0  <= I9ae27a7b654a36e4265449d861213978965e4cc3bc7f36b77c6a77cde5e24f77 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[8] ) begin
                    I119a98150511650722429eab31b5785e99128641bad59a3cb31e42158a648c48  <=  ~I9dd84c850b5e32710685c595cad935e3249afc0132b04ad8dec94cf13e16faf5 + 1;
                end else begin
                    I119a98150511650722429eab31b5785e99128641bad59a3cb31e42158a648c48  <= I9dd84c850b5e32710685c595cad935e3249afc0132b04ad8dec94cf13e16faf5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[11] ) begin
                    I6e418efd4b385b2a298c1c53d344e35f593e8380d1c27d7cb62cfe35223121c8  <=  ~Id59c354fd382f5bb1b276d565cfc2a0d55444ebe928c144c3d0b5513d53e3787 + 1;
                end else begin
                    I6e418efd4b385b2a298c1c53d344e35f593e8380d1c27d7cb62cfe35223121c8  <= Id59c354fd382f5bb1b276d565cfc2a0d55444ebe928c144c3d0b5513d53e3787 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5 != I4e9c85ad6975994daf65df213a2d2fa5a6a2abd91e66d9c9a6f540caf4c2afe2[0] ) begin
                    Ia695c63ae87e9a6742c6fecea648a214f5b24ea2b652bb5d83f35d9a59b94f72  <=  ~Idab4a7def7105c2e615a9138bf503482df9a2c434aa1ee7c4937acf6d0e6bac1 + 1;
                end else begin
                    Ia695c63ae87e9a6742c6fecea648a214f5b24ea2b652bb5d83f35d9a59b94f72  <= Idab4a7def7105c2e615a9138bf503482df9a2c434aa1ee7c4937acf6d0e6bac1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[20] ) begin
                    I34a89a8aa68b1657dc7137437574877b170659ebdbcc93a772989e2b8b5be31f  <=  ~I0d0ba52491ed5f98c69d74967cefc454cb2be9dc40bbc5bfe16c8ace0231dd70 + 1;
                end else begin
                    I34a89a8aa68b1657dc7137437574877b170659ebdbcc93a772989e2b8b5be31f  <= I0d0ba52491ed5f98c69d74967cefc454cb2be9dc40bbc5bfe16c8ace0231dd70 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[8] ) begin
                    I08e50de7e2aae48cc03a9959d08cab30d3c1c2ba8c4ef0799645787b0c09473c  <=  ~I05291a3275d232592dd880dda626cf60a03a62c655a2cf4b811f5325a07eb5e1 + 1;
                end else begin
                    I08e50de7e2aae48cc03a9959d08cab30d3c1c2ba8c4ef0799645787b0c09473c  <= I05291a3275d232592dd880dda626cf60a03a62c655a2cf4b811f5325a07eb5e1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[11] ) begin
                    I6f7aa66db409365eac05a200d0a0f1d2b25e9c37ba4a7db3b58a7298af0fd6e6  <=  ~I141f0199ad8f1dcd707f6b0553ebd7fd04217fb960f13cf25e98511ed91bc7aa + 1;
                end else begin
                    I6f7aa66db409365eac05a200d0a0f1d2b25e9c37ba4a7db3b58a7298af0fd6e6  <= I141f0199ad8f1dcd707f6b0553ebd7fd04217fb960f13cf25e98511ed91bc7aa ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f != Ic8f9966a2711f4810086d09b86e16ccf0d31339d146ad5c38d34c973c757947d[0] ) begin
                    Ifc31b600cbbf26e78cee82cd354c17b872586c1a53ddd132edbd25ce87d8aa9a  <=  ~I11a01802ccb6a01458a2cb2be3dea2f663acc531821edd809b95e10fb5a2def7 + 1;
                end else begin
                    Ifc31b600cbbf26e78cee82cd354c17b872586c1a53ddd132edbd25ce87d8aa9a  <= I11a01802ccb6a01458a2cb2be3dea2f663acc531821edd809b95e10fb5a2def7 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I99fb6dd2fc4414a231a70d23f26ed6b852ea4a563b41d3d8aa364e16d953eeb3 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[7] ) begin
                    I8600d4c5861319be0efba19d9b66ad483aa7bf648f2132c1a339157c43920c18  <=  ~Id76b3104f5a076b0f43f85da8b35a62b36a68d76bf8f26ff0667e085b37ce0e1 + 1;
                end else begin
                    I8600d4c5861319be0efba19d9b66ad483aa7bf648f2132c1a339157c43920c18  <= Id76b3104f5a076b0f43f85da8b35a62b36a68d76bf8f26ff0667e085b37ce0e1 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I99fb6dd2fc4414a231a70d23f26ed6b852ea4a563b41d3d8aa364e16d953eeb3 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[10] ) begin
                    I44ba42cf2460fce5fde6d8a9fba799517336268d29b5817597d819a9eb83df0e  <=  ~If5b73982b4248c4d2cc32bc28f0df8b37553ac0b034c0ebe3009bdfee069f642 + 1;
                end else begin
                    I44ba42cf2460fce5fde6d8a9fba799517336268d29b5817597d819a9eb83df0e  <= If5b73982b4248c4d2cc32bc28f0df8b37553ac0b034c0ebe3009bdfee069f642 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I99fb6dd2fc4414a231a70d23f26ed6b852ea4a563b41d3d8aa364e16d953eeb3 != Ic1385b7aee4e3b643e13733b56157e3e92e638da28cd1234e275fc9263709f04[0] ) begin
                    I261e70e693cdbc572e40e81c594f3dac624febb03465bfd0fb864d337e753499  <=  ~I9e3cbc961652bd76ec24ad12037b6384d8690af30372a8e0e5a93c57e4fb7b70 + 1;
                end else begin
                    I261e70e693cdbc572e40e81c594f3dac624febb03465bfd0fb864d337e753499  <= I9e3cbc961652bd76ec24ad12037b6384d8690af30372a8e0e5a93c57e4fb7b70 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If0e6db2779536df3835ac1e3c316bb7d9cf2e88aa7cb70f5b05563886cb4f3bb != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[7] ) begin
                    I434991f7c09dac3a7bd42fce3073dcbcf8b1c6579822074548ea94fdf1ef4eaa  <=  ~I7107302bbea73f0e5ff5ea2791a6d536cb04a165b68ef03ebeab0c0bfffe92cd + 1;
                end else begin
                    I434991f7c09dac3a7bd42fce3073dcbcf8b1c6579822074548ea94fdf1ef4eaa  <= I7107302bbea73f0e5ff5ea2791a6d536cb04a165b68ef03ebeab0c0bfffe92cd ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If0e6db2779536df3835ac1e3c316bb7d9cf2e88aa7cb70f5b05563886cb4f3bb != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[10] ) begin
                    I89cf2ce418b6d96c0e2b9c8e82167a47d40ade45a8f08255a1b849a9df9e6d06  <=  ~I561f05c657c3171c43fdfbb59215727da59d919f424597533b1890f7afe7cf07 + 1;
                end else begin
                    I89cf2ce418b6d96c0e2b9c8e82167a47d40ade45a8f08255a1b849a9df9e6d06  <= I561f05c657c3171c43fdfbb59215727da59d919f424597533b1890f7afe7cf07 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If0e6db2779536df3835ac1e3c316bb7d9cf2e88aa7cb70f5b05563886cb4f3bb != I3a173e6b224a6415ad442ae28a0af62756975427859bbcfc0af6c8e5effd62a6[0] ) begin
                    Ia6f7ae0adde8136c7a25f4fed69bbcaa376b5f28cbb4990afabb57a87ec03019  <=  ~I81789766f2008122a36b608dce3f08425ac203a154b4e43f915e0e3ef19fa022 + 1;
                end else begin
                    Ia6f7ae0adde8136c7a25f4fed69bbcaa376b5f28cbb4990afabb57a87ec03019  <= I81789766f2008122a36b608dce3f08425ac203a154b4e43f915e0e3ef19fa022 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I32eb2fcd88eff04a6295199db748b576fc1d585c2ae058acbf3150711574dd5d != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[7] ) begin
                    Id36acaa2c9161668c95e2cc3e6e852e9243ca7f486ca6c2ae4d124b1a8ddb522  <=  ~I678953f2ad317e167eea663eef2246d68cc67776d905877573ebcc39188a9a4d + 1;
                end else begin
                    Id36acaa2c9161668c95e2cc3e6e852e9243ca7f486ca6c2ae4d124b1a8ddb522  <= I678953f2ad317e167eea663eef2246d68cc67776d905877573ebcc39188a9a4d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I32eb2fcd88eff04a6295199db748b576fc1d585c2ae058acbf3150711574dd5d != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[10] ) begin
                    I4c02563233638e273f05bac3e277c702b38c204fda200dc5ac163662c77a429b  <=  ~I048fdd325368b2b72c83a32e9ac2c0208f392416f178445db74ceeafe56c8408 + 1;
                end else begin
                    I4c02563233638e273f05bac3e277c702b38c204fda200dc5ac163662c77a429b  <= I048fdd325368b2b72c83a32e9ac2c0208f392416f178445db74ceeafe56c8408 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I32eb2fcd88eff04a6295199db748b576fc1d585c2ae058acbf3150711574dd5d != Ia5580120af4590da8aed890f81ca17929e4c998617df957686c095e891649c83[0] ) begin
                    Ic40e94217a2d2c13f4b1ad2766ab1ae4e8ded0b5e0a3522dd51ec806c3e9feef  <=  ~I16b1a9836d7b38707938eb48bf60f17f049403d2fd29d5245798fd1ade1c2531 + 1;
                end else begin
                    Ic40e94217a2d2c13f4b1ad2766ab1ae4e8ded0b5e0a3522dd51ec806c3e9feef  <= I16b1a9836d7b38707938eb48bf60f17f049403d2fd29d5245798fd1ade1c2531 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I244e0f2c03df982bd121a8a0240f862b4e0212ab54dbec0984f987577faebeb2 != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[7] ) begin
                    I30e30c2bee3bac86dd68fe8364f818ab63e91d65c4fa1ef45fcfd03c9df87cc5  <=  ~I48c21b6fc24c93dae3a01b55b280508297e0ff5101c7fbc7d17e823d9a31fb07 + 1;
                end else begin
                    I30e30c2bee3bac86dd68fe8364f818ab63e91d65c4fa1ef45fcfd03c9df87cc5  <= I48c21b6fc24c93dae3a01b55b280508297e0ff5101c7fbc7d17e823d9a31fb07 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I244e0f2c03df982bd121a8a0240f862b4e0212ab54dbec0984f987577faebeb2 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[10] ) begin
                    I3f92074e96f2c2711248b1d770b4ad718a565a323e6fe4ebb379e6494039af47  <=  ~I9d5c1ef1f35b4d40b4f20dcd2c33691152683bf308c95aa53adbf785defb75ef + 1;
                end else begin
                    I3f92074e96f2c2711248b1d770b4ad718a565a323e6fe4ebb379e6494039af47  <= I9d5c1ef1f35b4d40b4f20dcd2c33691152683bf308c95aa53adbf785defb75ef ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I244e0f2c03df982bd121a8a0240f862b4e0212ab54dbec0984f987577faebeb2 != I58a3910d475757bccbde2da0e6b5dd5723cbe44e1f4d3e71ac2973fd2a03b3a8[0] ) begin
                    I78602c68a4a00f530bda7ba1dfa4820b7faeb0edabc636d6a2d8bf97005755d1  <=  ~Iec1baa5364573d0a9866494a039a3409a32b4665d4a79e2a729b54d370ecad97 + 1;
                end else begin
                    I78602c68a4a00f530bda7ba1dfa4820b7faeb0edabc636d6a2d8bf97005755d1  <= Iec1baa5364573d0a9866494a039a3409a32b4665d4a79e2a729b54d370ecad97 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[21] ) begin
                    I2747ce9b7349ed89e3265df62bb0d0e612706d8c1b61e30a2878094662da8ff1  <=  ~I508c79d6f4d56ea0e8100825c438214e4b5087004f8a5041b4beb900509cfde8 + 1;
                end else begin
                    I2747ce9b7349ed89e3265df62bb0d0e612706d8c1b61e30a2878094662da8ff1  <= I508c79d6f4d56ea0e8100825c438214e4b5087004f8a5041b4beb900509cfde8 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[12] ) begin
                    Ibae97ff31fce14dd0506fdfe7407fd6260f7cf8584a01da77312b1aa48594be0  <=  ~Id55510ec558d15440325660ab2ac2cd9d4dd682c082479a742118c9ba1923cae + 1;
                end else begin
                    Ibae97ff31fce14dd0506fdfe7407fd6260f7cf8584a01da77312b1aa48594be0  <= Id55510ec558d15440325660ab2ac2cd9d4dd682c082479a742118c9ba1923cae ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[14] ) begin
                    If072f43c0b06c41c30d9bc40dae674ad9052e5533b1308adb97cff2e03821bab  <=  ~I000c117a768755741005775b84eb6e4c406d2e29765ca9bbab991217963de8d2 + 1;
                end else begin
                    If072f43c0b06c41c30d9bc40dae674ad9052e5533b1308adb97cff2e03821bab  <= I000c117a768755741005775b84eb6e4c406d2e29765ca9bbab991217963de8d2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027 != I1b76b0f61e714e21a844e429806d641f6a24f0eb19c23a3c2fcfb76baaf3e72a[0] ) begin
                    Id8e684d92e6d0b6e10b5e7f7ff9656e6fc67c99edaa59b49e453844ae33d23f6  <=  ~I95d510e99cd368229106d7ef60f9438bc186adb5359c9483b645b255a769df90 + 1;
                end else begin
                    Id8e684d92e6d0b6e10b5e7f7ff9656e6fc67c99edaa59b49e453844ae33d23f6  <= I95d510e99cd368229106d7ef60f9438bc186adb5359c9483b645b255a769df90 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[21] ) begin
                    I23e0423ae4012d108a4e6a495814e0e6f920fa6dcab900bb35cba7b95f590c9b  <=  ~I4cb9b54295972404ff2984e0b2a225773e067803925fc434674a5ef2439df4c3 + 1;
                end else begin
                    I23e0423ae4012d108a4e6a495814e0e6f920fa6dcab900bb35cba7b95f590c9b  <= I4cb9b54295972404ff2984e0b2a225773e067803925fc434674a5ef2439df4c3 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[12] ) begin
                    I5c43417b1bd96dfedeb36f6d3405fc7f6b73c11a55f21ebe6ffd675e991a13c3  <=  ~Ied36baf05b90f7d785653eb1e7f699cfa84cd0a1eb3a985047f57e2885dad2ef + 1;
                end else begin
                    I5c43417b1bd96dfedeb36f6d3405fc7f6b73c11a55f21ebe6ffd675e991a13c3  <= Ied36baf05b90f7d785653eb1e7f699cfa84cd0a1eb3a985047f57e2885dad2ef ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[14] ) begin
                    I13a54b612481fe0fdfe8b52909179bb82298c2bff4f10adc4f41215fa4396311  <=  ~Id3947617c14deada0b43f71b47e700dbd8a1ac15820eed783d58774c249d5f24 + 1;
                end else begin
                    I13a54b612481fe0fdfe8b52909179bb82298c2bff4f10adc4f41215fa4396311  <= Id3947617c14deada0b43f71b47e700dbd8a1ac15820eed783d58774c249d5f24 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f != If0211848e6cda136970069df5b6156d4ac213717491c68ed49ab39d2cffe9999[0] ) begin
                    Ic9d9001a209401fca8a3f28e39c4b89adc8f4e9d225aeffbb5d30893bea1a7b2  <=  ~I846f9754b91cbdf37fc2662d5851bfffa4926c1ef01f4a23f20b02d9588ff3d4 + 1;
                end else begin
                    Ic9d9001a209401fca8a3f28e39c4b89adc8f4e9d225aeffbb5d30893bea1a7b2  <= I846f9754b91cbdf37fc2662d5851bfffa4926c1ef01f4a23f20b02d9588ff3d4 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[21] ) begin
                    I6b4d2a32c92c22b1cfe81ee6620c69af1850621deea406d75f098da0542843e8  <=  ~I7485137b6eb30fbd6f06453139f9cd1ebeec411e566936bc598f0aefde881251 + 1;
                end else begin
                    I6b4d2a32c92c22b1cfe81ee6620c69af1850621deea406d75f098da0542843e8  <= I7485137b6eb30fbd6f06453139f9cd1ebeec411e566936bc598f0aefde881251 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66 != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[12] ) begin
                    I294ca1e2c287bbe18783f7043149078d4fcc1c59e24792d75655fb29a36e33d4  <=  ~I152ada5197e26088aadb2058a128099d201dc6e91d564b80b8e3930567a1a929 + 1;
                end else begin
                    I294ca1e2c287bbe18783f7043149078d4fcc1c59e24792d75655fb29a36e33d4  <= I152ada5197e26088aadb2058a128099d201dc6e91d564b80b8e3930567a1a929 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[14] ) begin
                    I4e5dfe1c7112e24769a5e6aa86584c09ed659fa5d05af38d18183db31189a3a7  <=  ~Ic86eed327a12ce5bd475a6b82a5bdc31777526455fb541a8f4e842605bb34ddf + 1;
                end else begin
                    I4e5dfe1c7112e24769a5e6aa86584c09ed659fa5d05af38d18183db31189a3a7  <= Ic86eed327a12ce5bd475a6b82a5bdc31777526455fb541a8f4e842605bb34ddf ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66 != Id23ae21f713f4f452abcb1c1839b5524c452bb8bb0b6c35683f9bde212bc5f96[0] ) begin
                    I97f666707f6afacfc6156ef498941fe5feeb7424834b4a283139aefb5f50a68f  <=  ~Ic1a3e7a14eff1a6da9e96ddbd750086b011cdc44e8aa1189879b056fc48b3a27 + 1;
                end else begin
                    I97f666707f6afacfc6156ef498941fe5feeb7424834b4a283139aefb5f50a68f  <= Ic1a3e7a14eff1a6da9e96ddbd750086b011cdc44e8aa1189879b056fc48b3a27 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[21] ) begin
                    I6ed6ee11f6983e96e7ccc4e4be6ed8c4ed166ca9075b9cd218f26f018ad2140f  <=  ~I215ee2b19d3ea96eedc62d8cb097051dad2d917dfb2eb2b0e1ed0ff697955765 + 1;
                end else begin
                    I6ed6ee11f6983e96e7ccc4e4be6ed8c4ed166ca9075b9cd218f26f018ad2140f  <= I215ee2b19d3ea96eedc62d8cb097051dad2d917dfb2eb2b0e1ed0ff697955765 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[12] ) begin
                    Id8da43222903044cc48243a7bcce7864e66d151673396879258ee4af7008a706  <=  ~Ibbfd537ee459654bacd89b68f7d66565efcbdaa3838dc0847f83ba17c49b404b + 1;
                end else begin
                    Id8da43222903044cc48243a7bcce7864e66d151673396879258ee4af7008a706  <= Ibbfd537ee459654bacd89b68f7d66565efcbdaa3838dc0847f83ba17c49b404b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[14] ) begin
                    I66291192ca8d81c8e3f667651d5201cb41b6872f73283d13c6718159b008d8cf  <=  ~Iccf845c102c65fc97a1244cb2c0182925c72e95fb4a9b0dc97379f5a32837612 + 1;
                end else begin
                    I66291192ca8d81c8e3f667651d5201cb41b6872f73283d13c6718159b008d8cf  <= Iccf845c102c65fc97a1244cb2c0182925c72e95fb4a9b0dc97379f5a32837612 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a != Id5bdb0f5a920710b1af7cc3abade245196df9d1ab4b7f26277fd93e1bbee5556[0] ) begin
                    Ibdaeb96b71f9ccccfe79b1b3bab77122aa32217b58037d80a3183bf888b60c72  <=  ~I32562e9f1cb6c7224d2efbd29f393e04c0d655e4bef402c2689cb946013f5d1f + 1;
                end else begin
                    Ibdaeb96b71f9ccccfe79b1b3bab77122aa32217b58037d80a3183bf888b60c72  <= I32562e9f1cb6c7224d2efbd29f393e04c0d655e4bef402c2689cb946013f5d1f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228 != Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[21] ) begin
                    I9f9d895211b42c2c9d491349dbe7aafbad775942920197105c34837dba6563a0  <=  ~I8ee1c7843334dc659003797fc7ec177037e184855e8e80063c6e490425de9446 + 1;
                end else begin
                    I9f9d895211b42c2c9d491349dbe7aafbad775942920197105c34837dba6563a0  <= I8ee1c7843334dc659003797fc7ec177037e184855e8e80063c6e490425de9446 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228 != I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[12] ) begin
                    Ifd66abca1532f04fc777617d91cd2d5f4d4fee35c3f075e91639a196780168d8  <=  ~I5c6a9cfeb6a0354276fa86b65ea21b018e71d37b366f907012b41156aa22bfcb + 1;
                end else begin
                    Ifd66abca1532f04fc777617d91cd2d5f4d4fee35c3f075e91639a196780168d8  <= I5c6a9cfeb6a0354276fa86b65ea21b018e71d37b366f907012b41156aa22bfcb ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228 != I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[8] ) begin
                    I06a5cdf2e430e40b5c08ab617356f6b4b0389236041b77e2a57d9d314bfe77f3  <=  ~I76041755b112a333460289875673d3f2b054918770d3a2cc46ab7a9f92b50eb5 + 1;
                end else begin
                    I06a5cdf2e430e40b5c08ab617356f6b4b0389236041b77e2a57d9d314bfe77f3  <= I76041755b112a333460289875673d3f2b054918770d3a2cc46ab7a9f92b50eb5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228 != Ic72616171e7fb8489fa12cc29be1f74602ff8e4bd28ea085e938da615238a0fa[0] ) begin
                    I574e4843ab81be7ad95cb7027fc3284a8780b07fb8a194a9c991997988d7ff8f  <=  ~I30843beae9ebf34c0f73f773e1af0422e40b3ced201574b6f87f400cb37a7175 + 1;
                end else begin
                    I574e4843ab81be7ad95cb7027fc3284a8780b07fb8a194a9c991997988d7ff8f  <= I30843beae9ebf34c0f73f773e1af0422e40b3ced201574b6f87f400cb37a7175 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40 != Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[21] ) begin
                    I31009872a3e84f78bbf1f12a7da708c45e3b708bd943b6f4561ad436164b12d8  <=  ~I7f99ba04346760d4ee2589662be79b19673e741f07d1b9c0c35b54d4bcd3cfc0 + 1;
                end else begin
                    I31009872a3e84f78bbf1f12a7da708c45e3b708bd943b6f4561ad436164b12d8  <= I7f99ba04346760d4ee2589662be79b19673e741f07d1b9c0c35b54d4bcd3cfc0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40 != I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[12] ) begin
                    Ib1e319af12dcd98c09841e8b06e7af86f2569bd7afeb1718bbbd26e30f65c464  <=  ~I311c88c2854536dbb8f578bdf98823eaf5888a7c772bc2c6f0cb49c9c9c79500 + 1;
                end else begin
                    Ib1e319af12dcd98c09841e8b06e7af86f2569bd7afeb1718bbbd26e30f65c464  <= I311c88c2854536dbb8f578bdf98823eaf5888a7c772bc2c6f0cb49c9c9c79500 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40 != I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[8] ) begin
                    I6106f96669a63f337b78a6bad5894881230f0ab6467c23ec877cf27a5bc76cb6  <=  ~I073f480ce57215d8a9930ab34bbed6bcf5e631613fced0e782749a390615672c + 1;
                end else begin
                    I6106f96669a63f337b78a6bad5894881230f0ab6467c23ec877cf27a5bc76cb6  <= I073f480ce57215d8a9930ab34bbed6bcf5e631613fced0e782749a390615672c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40 != Ia09db6bd7cba6c6e15cac4c6ad0d4c98235a7437beeabca1388fb1b4dece5d67[0] ) begin
                    Iaa4463f258ed92a2c85fef0790c47e725c555f37c80dbe366d973c9599a5484d  <=  ~Iaef86ab80a38f09821c64eb7b93cf066c0ba40a4b315075fd4652eb82b687bff + 1;
                end else begin
                    Iaa4463f258ed92a2c85fef0790c47e725c555f37c80dbe366d973c9599a5484d  <= Iaef86ab80a38f09821c64eb7b93cf066c0ba40a4b315075fd4652eb82b687bff ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b != I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[21] ) begin
                    I8d91c857f2c8154bb09d456ff73ebdf81e3b7d9bd1c57c2e6b8c2de74e55cf48  <=  ~Id523ce79d9f7a6b24c5979c58855211eb2bde238c81e549064c23ec62a5c7a3d + 1;
                end else begin
                    I8d91c857f2c8154bb09d456ff73ebdf81e3b7d9bd1c57c2e6b8c2de74e55cf48  <= Id523ce79d9f7a6b24c5979c58855211eb2bde238c81e549064c23ec62a5c7a3d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b != Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[12] ) begin
                    I3386ee46348e8c4359b1ea2153bc64afbe76f2b6bc9a312629b8c52762a22873  <=  ~Id27c2a1647e08c46fba102b41eceb3513a697df9876d76b23fc4118f16b479a0 + 1;
                end else begin
                    I3386ee46348e8c4359b1ea2153bc64afbe76f2b6bc9a312629b8c52762a22873  <= Id27c2a1647e08c46fba102b41eceb3513a697df9876d76b23fc4118f16b479a0 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b != I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[8] ) begin
                    I45a11cd2f581121ac03fe112ec78bd07c070673712fe6112a3e4fb4eba298e27  <=  ~I54a09dd4115c1f70cff7fd7921120216494997fbc08a7e9eb8e59152ef12a9e6 + 1;
                end else begin
                    I45a11cd2f581121ac03fe112ec78bd07c070673712fe6112a3e4fb4eba298e27  <= I54a09dd4115c1f70cff7fd7921120216494997fbc08a7e9eb8e59152ef12a9e6 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b != I15ab76f6e4824af9b3b4f5062e8dd3c426e1ff0c5f68e4733828c710eb7bca54[0] ) begin
                    I7102386e760e34e2d0fc4563b497acec7222bd171333a2169fac800df94ea27c  <=  ~I5a2063e62c2c96b172ecad9fa950c0b42c413214e30d94796ca9c2b8c6bbe522 + 1;
                end else begin
                    I7102386e760e34e2d0fc4563b497acec7222bd171333a2169fac800df94ea27c  <= I5a2063e62c2c96b172ecad9fa950c0b42c413214e30d94796ca9c2b8c6bbe522 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6 != I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[21] ) begin
                    I1b93b1b2c5f55e2267a4deb4f75ca91039d6893af8e082ea85b7a5e9354117e6  <=  ~If0c2c0785586996991da246fc01722deded4e3ca8550290626324c5908d770a5 + 1;
                end else begin
                    I1b93b1b2c5f55e2267a4deb4f75ca91039d6893af8e082ea85b7a5e9354117e6  <= If0c2c0785586996991da246fc01722deded4e3ca8550290626324c5908d770a5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6 != I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[12] ) begin
                    I03929e638a59a35fc0168772ca06f7a502352e03525042ce6d49cf9ecb671093  <=  ~Icb2218fe2214af22ea6fff2b9ff3c8d1772fd9318efa83c7655b0dfee2f6ab4d + 1;
                end else begin
                    I03929e638a59a35fc0168772ca06f7a502352e03525042ce6d49cf9ecb671093  <= Icb2218fe2214af22ea6fff2b9ff3c8d1772fd9318efa83c7655b0dfee2f6ab4d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6 != I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[8] ) begin
                    I6c6885b180013a16955ddefa0dc75c25ac85fb76059df9bf8b63af72c8c1fb4d  <=  ~I0c567cd54c6fded476f507a4a35d7d93fdbd2cd1c555e10edf313ddaf4b0d64f + 1;
                end else begin
                    I6c6885b180013a16955ddefa0dc75c25ac85fb76059df9bf8b63af72c8c1fb4d  <= I0c567cd54c6fded476f507a4a35d7d93fdbd2cd1c555e10edf313ddaf4b0d64f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6 != I12b276cd6b0aa86ca2e28dbb1f4008ab140668e16e4ef96604a6d1741c7f2f95[0] ) begin
                    Iee34d958bf4feec1e5bde8a866a9919f29edd54f1bc51cc9c8216b71101d640b  <=  ~Ic49fb172f5523a522e94efd83b5827b8f63c2d8fd7c76263249d96a00a0e25ad + 1;
                end else begin
                    Iee34d958bf4feec1e5bde8a866a9919f29edd54f1bc51cc9c8216b71101d640b  <= Ic49fb172f5523a522e94efd83b5827b8f63c2d8fd7c76263249d96a00a0e25ad ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50 != I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[9] ) begin
                    I28a2b1ada19dc69ebe4949a75633b2f543159d2d1cc169f3bb6070c1419878e0  <=  ~Ibef81155a593cc991eb8f0da7ea8dbc27f3c935dc1fdf7b857110407ef449718 + 1;
                end else begin
                    I28a2b1ada19dc69ebe4949a75633b2f543159d2d1cc169f3bb6070c1419878e0  <= Ibef81155a593cc991eb8f0da7ea8dbc27f3c935dc1fdf7b857110407ef449718 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50 != I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[8] ) begin
                    Ic551d228c593c4304b4ef79a965ac1d9081774282af09d79cd587ef9abcd6003  <=  ~Id1c35604f896316440f1deadc55ea39d16307edf0e2ddea1d7d450c41dbbc705 + 1;
                end else begin
                    Ic551d228c593c4304b4ef79a965ac1d9081774282af09d79cd587ef9abcd6003  <= Id1c35604f896316440f1deadc55ea39d16307edf0e2ddea1d7d450c41dbbc705 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50 != Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[11] ) begin
                    I47ba4d6ad7b1889cb52ff7a1d42176e166270e39a1d2875f3a0cd260a1fc92ab  <=  ~Ic00c95647ac3595e199e62c4d3e75956755ac952e4cea464b27066ad8f09415f + 1;
                end else begin
                    I47ba4d6ad7b1889cb52ff7a1d42176e166270e39a1d2875f3a0cd260a1fc92ab  <= Ic00c95647ac3595e199e62c4d3e75956755ac952e4cea464b27066ad8f09415f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50 != I01577c8c0e65ca47449450a8b2455ee84cf5c48bb26a0799b5523258a039ae40[0] ) begin
                    I64b0ef6642050de0690c95be2af9606797be36c1656f1306b87ce3e8131c4629  <=  ~I4d89a637472e8c4d071c44792883afdac1fe1c6ffa9d08f7259525884000b34e + 1;
                end else begin
                    I64b0ef6642050de0690c95be2af9606797be36c1656f1306b87ce3e8131c4629  <= I4d89a637472e8c4d071c44792883afdac1fe1c6ffa9d08f7259525884000b34e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f != Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[9] ) begin
                    Ibf22dd3f14f19c3fc769966f72e8ec980dc79c2991f69d03ca2defb7f720f880  <=  ~I081fd1385ec974da04b64bc5764efd6db252fefa40f518ed0ed4b01ce630064a + 1;
                end else begin
                    Ibf22dd3f14f19c3fc769966f72e8ec980dc79c2991f69d03ca2defb7f720f880  <= I081fd1385ec974da04b64bc5764efd6db252fefa40f518ed0ed4b01ce630064a ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f != Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[8] ) begin
                    I7fec897140c79264b7b7b7f3ae228ed090ff69351985c07d317ff9c0cab1e58c  <=  ~I57c394b657ecd32691fcef200ba361abaffca7d8ddbc7bea22502a9f7bff9f5f + 1;
                end else begin
                    I7fec897140c79264b7b7b7f3ae228ed090ff69351985c07d317ff9c0cab1e58c  <= I57c394b657ecd32691fcef200ba361abaffca7d8ddbc7bea22502a9f7bff9f5f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f != I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[11] ) begin
                    I85d8f259f770b22a380d6eb5ace0281c57f0952506152be05f38482c47334988  <=  ~Ia14c31a81641330844c0c48e155c6f7630695ccf3e7238ad6eca01c8a45a104e + 1;
                end else begin
                    I85d8f259f770b22a380d6eb5ace0281c57f0952506152be05f38482c47334988  <= Ia14c31a81641330844c0c48e155c6f7630695ccf3e7238ad6eca01c8a45a104e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f != I63ba87cd2daa7c3c625d3ff5bdaca7f2115fc2d65e13972a22b2c2ae5b746d4a[0] ) begin
                    I23f31ebee34c7f4f9c46fba41d41df176a7465c074ad8527205a5782edab6524  <=  ~Iffdff1b757352d5f1174deb338f337fd8841ce8d132c2e0a16f18fc1a97313a2 + 1;
                end else begin
                    I23f31ebee34c7f4f9c46fba41d41df176a7465c074ad8527205a5782edab6524  <= Iffdff1b757352d5f1174deb338f337fd8841ce8d132c2e0a16f18fc1a97313a2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5 != I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[9] ) begin
                    Ieee1d2436dbda6f58f19df70b691a4ff28d37db8ccc12e04413e45f80d7124e0  <=  ~If8c3dafd18d6fabac3e4ec4dce257aba397ab0d341e25a1bb88f9e32909deb17 + 1;
                end else begin
                    Ieee1d2436dbda6f58f19df70b691a4ff28d37db8ccc12e04413e45f80d7124e0  <= If8c3dafd18d6fabac3e4ec4dce257aba397ab0d341e25a1bb88f9e32909deb17 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5 != Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[8] ) begin
                    I325ec6d7bab5ccd6e9c4a7e9b02a3b8c30072df123bf6318bd97f1e8766457c8  <=  ~Ie4b741e2c3f5dbd43bba89fbaeb4cc6b309042b53629f8db67121eb22a656ee9 + 1;
                end else begin
                    I325ec6d7bab5ccd6e9c4a7e9b02a3b8c30072df123bf6318bd97f1e8766457c8  <= Ie4b741e2c3f5dbd43bba89fbaeb4cc6b309042b53629f8db67121eb22a656ee9 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5 != I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[11] ) begin
                    Ia478acf4034b69d392277c3d5c6683346547ff26d418b3a6c36a3f9a56e3cfe0  <=  ~Ib1a3877a6c9f5b87fd3c2104782a0699748b68ef73a12291b34e914344db9d25 + 1;
                end else begin
                    Ia478acf4034b69d392277c3d5c6683346547ff26d418b3a6c36a3f9a56e3cfe0  <= Ib1a3877a6c9f5b87fd3c2104782a0699748b68ef73a12291b34e914344db9d25 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5 != I576afeb6020cc0a8e35837b4b96968ed04cd444999558626adac849848fe7c6c[0] ) begin
                    I628b9674d7d6caaa70c54539241df2e7a4be0441dde1739b442513c6e4ded8a4  <=  ~Ieab221c067f0649e88f307dd8c46981653088853874e2a256b99f7b7a8bf93d5 + 1;
                end else begin
                    I628b9674d7d6caaa70c54539241df2e7a4be0441dde1739b442513c6e4ded8a4  <= Ieab221c067f0649e88f307dd8c46981653088853874e2a256b99f7b7a8bf93d5 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18 != I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[9] ) begin
                    I47b54f01ac82a9eb80a681633a06c4e1d432d358091e9d079f74484f40ab3e09  <=  ~Ic80161feee5be9576086dd9d1ed8adca369a841f0052af01b2fe93d46af669b2 + 1;
                end else begin
                    I47b54f01ac82a9eb80a681633a06c4e1d432d358091e9d079f74484f40ab3e09  <= Ic80161feee5be9576086dd9d1ed8adca369a841f0052af01b2fe93d46af669b2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18 != I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[8] ) begin
                    Ic0bef9008769fe36d726cf80506004d66e7c843a046653201c9bc2c816115c28  <=  ~Iac4628a0a7bdc975990c2664a736112cdb2bf1b1b30f89ae1e6827a44bdb4474 + 1;
                end else begin
                    Ic0bef9008769fe36d726cf80506004d66e7c843a046653201c9bc2c816115c28  <= Iac4628a0a7bdc975990c2664a736112cdb2bf1b1b30f89ae1e6827a44bdb4474 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18 != Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[11] ) begin
                    Ie4fafd34aeca2efbfd3bfd3bf45f73ceea27b613ed242a43666d85f3680ada44  <=  ~I7da6920e7bb85e837e61b04ba09453237164470bf2eb7607af94194e05407bfe + 1;
                end else begin
                    Ie4fafd34aeca2efbfd3bfd3bf45f73ceea27b613ed242a43666d85f3680ada44  <= I7da6920e7bb85e837e61b04ba09453237164470bf2eb7607af94194e05407bfe ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18 != I3b8769ce28405c0bb978c458bd6272f10cea5338af4170ce4e93a8932ae8dcaf[0] ) begin
                    Ib066c9d790586949b27c4cf09dc957e7d28161ab00e8dc6920e4e0cc5ac665d9  <=  ~Ie3ca82b8d601f023d408833c7b5445539ebf8f17bb678e486fb3f650b2e01d9d + 1;
                end else begin
                    Ib066c9d790586949b27c4cf09dc957e7d28161ab00e8dc6920e4e0cc5ac665d9  <= Ie3ca82b8d601f023d408833c7b5445539ebf8f17bb678e486fb3f650b2e01d9d ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728 != Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[22] ) begin
                    Ia0964979ac559942d1da1c41ecb3d9e94c6c7c0da3d16177cf2379db8f37aa65  <=  ~Ifc8ba6aad04e3418146443a14c520552e32ac2f43fabe430ef0d640b4262337e + 1;
                end else begin
                    Ia0964979ac559942d1da1c41ecb3d9e94c6c7c0da3d16177cf2379db8f37aa65  <= Ifc8ba6aad04e3418146443a14c520552e32ac2f43fabe430ef0d640b4262337e ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728 != Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[13] ) begin
                    I8eb86c8d64d83d4ac46667af42b6383e4d165459475ec6be9d547a70ef0248af  <=  ~If1aa1bf1d7206ef9c00f8c1aafd738c03603858f9757a3f671242af1b139cc64 + 1;
                end else begin
                    I8eb86c8d64d83d4ac46667af42b6383e4d165459475ec6be9d547a70ef0248af  <= If1aa1bf1d7206ef9c00f8c1aafd738c03603858f9757a3f671242af1b139cc64 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728 != If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[15] ) begin
                    I2f05dd0209278c1e661998552da73728c1521c024a7d26f4652d4f151c6e5f80  <=  ~I97205d95f7ff115112b2b1a7eb32bf70ff7c1e2fb431785547ed7f98d5fea0af + 1;
                end else begin
                    I2f05dd0209278c1e661998552da73728c1521c024a7d26f4652d4f151c6e5f80  <= I97205d95f7ff115112b2b1a7eb32bf70ff7c1e2fb431785547ed7f98d5fea0af ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728 != Ib4638612fcabc0a2c2f2bba5a2b9eb71cdea23575641b3f81fb6220fcaf284f4[0] ) begin
                    I57419941b1979cd06c4fa0e6be943f004dd80da502425ee5b6dabd2239139cd7  <=  ~Ia6232cf34275276641c494e4f4cbd7a8796f1f946733ed0fe15d9e11cd8c740f + 1;
                end else begin
                    I57419941b1979cd06c4fa0e6be943f004dd80da502425ee5b6dabd2239139cd7  <= Ia6232cf34275276641c494e4f4cbd7a8796f1f946733ed0fe15d9e11cd8c740f ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6 != I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[22] ) begin
                    I0678dba3dc1a3400ab26e223257bf71c03f0e8d284810653b5e507fe964427f4  <=  ~I24883a74ba0e0eaf8efff93301dd4d714667c28020ff65d73e4056b2d014e287 + 1;
                end else begin
                    I0678dba3dc1a3400ab26e223257bf71c03f0e8d284810653b5e507fe964427f4  <= I24883a74ba0e0eaf8efff93301dd4d714667c28020ff65d73e4056b2d014e287 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6 != Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[13] ) begin
                    Iea011619fa5b0fb7d22dc4bb4ce3fcc4856dfc7286ff393fb329ac0d7e348207  <=  ~Ibdd97caada239a1152f2155c8cb9e25402600931810f6bafe34159894246d962 + 1;
                end else begin
                    Iea011619fa5b0fb7d22dc4bb4ce3fcc4856dfc7286ff393fb329ac0d7e348207  <= Ibdd97caada239a1152f2155c8cb9e25402600931810f6bafe34159894246d962 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6 != Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[15] ) begin
                    I26a27b64a7aafdbcf4a6d058181fb84e0e16767f4bd7a9c45211c4c1246d3b9e  <=  ~I4ba3a78d1129b6b95ec4421b8dc75b90921b67ed09cc636c1fe08c778c9a4c87 + 1;
                end else begin
                    I26a27b64a7aafdbcf4a6d058181fb84e0e16767f4bd7a9c45211c4c1246d3b9e  <= I4ba3a78d1129b6b95ec4421b8dc75b90921b67ed09cc636c1fe08c778c9a4c87 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6 != I16ea389c88e4591f7686eae3f1988dd5361bf893895697c0ade8627986a9fc5e[0] ) begin
                    Iabb5703a54942b1bdcfe2213d2011c659ec812f751dc75943b2ce511c81ffaf9  <=  ~Ia8fe4e59fc4b364c711cdef5a6718ae33543de2e35744d9cda4cf33f340d7add + 1;
                end else begin
                    Iabb5703a54942b1bdcfe2213d2011c659ec812f751dc75943b2ce511c81ffaf9  <= Ia8fe4e59fc4b364c711cdef5a6718ae33543de2e35744d9cda4cf33f340d7add ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205 != I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[22] ) begin
                    I3619e836fee4be75d6700a0e72e84df3a5a61003227363b8c4d348b8353075e0  <=  ~Ib0319b3fbdfab7c4df3ba7c1d710d7ca176cf8cd4223ea11fe12102cb5ac7f12 + 1;
                end else begin
                    I3619e836fee4be75d6700a0e72e84df3a5a61003227363b8c4d348b8353075e0  <= Ib0319b3fbdfab7c4df3ba7c1d710d7ca176cf8cd4223ea11fe12102cb5ac7f12 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205 != I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[13] ) begin
                    I71f31c9a9943d9fd422d00aa01888aac32dd8b34236bdd9bdf3e660413a3512a  <=  ~Ice9d3685b31919d1cfe76a96ac6e1738ef6c66e069de55830f61665cb5bc0ca2 + 1;
                end else begin
                    I71f31c9a9943d9fd422d00aa01888aac32dd8b34236bdd9bdf3e660413a3512a  <= Ice9d3685b31919d1cfe76a96ac6e1738ef6c66e069de55830f61665cb5bc0ca2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205 != Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[15] ) begin
                    Iff97998b0778cb649d03228ed3acc81c1b3a97f6bc47041c423120b1311112d0  <=  ~I36a3a77efd095e4c91274958f1ed4b9fc929f2b6794e4b879b8275f3a01ae48c + 1;
                end else begin
                    Iff97998b0778cb649d03228ed3acc81c1b3a97f6bc47041c423120b1311112d0  <= I36a3a77efd095e4c91274958f1ed4b9fc929f2b6794e4b879b8275f3a01ae48c ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205 != Ia17edf214ab782c25bbab97f6bb4e04b2fc46d41f9a97fcf617418d54ab76a7e[0] ) begin
                    I798a6a6074b50fc61bd4e1b4696560abd2e515c86d47f85e9a3077cf6672acc8  <=  ~I0643791cd1c7ee5c205da45ee4720229c6f7b61e98a7f642afc47506f6e10210 + 1;
                end else begin
                    I798a6a6074b50fc61bd4e1b4696560abd2e515c86d47f85e9a3077cf6672acc8  <= I0643791cd1c7ee5c205da45ee4720229c6f7b61e98a7f642afc47506f6e10210 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d != I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[22] ) begin
                    I571233769cc63838bcc3d61e7a5e95805c3f4116c0053dfe86831eafff7c32fe  <=  ~I485c81ca3402c9b70ad8a10b749c0ee5e81569d1a64231a5fb25e3af8cc4abba + 1;
                end else begin
                    I571233769cc63838bcc3d61e7a5e95805c3f4116c0053dfe86831eafff7c32fe  <= I485c81ca3402c9b70ad8a10b749c0ee5e81569d1a64231a5fb25e3af8cc4abba ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d != I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[13] ) begin
                    Ideae854591637828f033505e4fc9dee34d82369d02f7680ef6887c597ac1ac82  <=  ~Ief695bef8a02a4f5e89c14ac6b89f84678cc7d7a9d71bf2a5e3c1abd44d1cbb2 + 1;
                end else begin
                    Ideae854591637828f033505e4fc9dee34d82369d02f7680ef6887c597ac1ac82  <= Ief695bef8a02a4f5e89c14ac6b89f84678cc7d7a9d71bf2a5e3c1abd44d1cbb2 ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d != I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[15] ) begin
                    I4bfef3f43cb1a77ce8b2bf4b26160a161e7f28308b8d2817e6e2840f09463e37  <=  ~I0ce015383446aeba50b7677c9060a1e18dab91eb8040a718fcb7e104a700c29b + 1;
                end else begin
                    I4bfef3f43cb1a77ce8b2bf4b26160a161e7f28308b8d2817e6e2840f09463e37  <= I0ce015383446aeba50b7677c9060a1e18dab91eb8040a718fcb7e104a700c29b ;
                end
             end
             if (If95958c4bb278a7461a73692815e09d6e0ade514cfbee5da62532d1e8a371458) begin
                if (Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d != Ibcfba9f1fb81d976955a1fa7101f0b0db16c344c82cc5ce81f50dd3aa2928d37[0] ) begin
                    I3f4a8ec7c554b1f0b9d3d2963b0e3dec4654bf07c5b836f8fd07c639cd19d588  <=  ~I9f790cf09f0d8b1c047cd0df401052898d374d930d5ccd784d142c544d8b54b6 + 1;
                end else begin
                    I3f4a8ec7c554b1f0b9d3d2963b0e3dec4654bf07c5b836f8fd07c639cd19d588  <= I9f790cf09f0d8b1c047cd0df401052898d374d930d5ccd784d142c544d8b54b6 ;
                end
             end
       end
   end


   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[0]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[1]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[2]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[3]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[4]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[5]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[6]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[7]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[8]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[9]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[10]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[11]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[12]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[13]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[14]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[15]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[16]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[17]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[18]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[19]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[20]  <= 1'b0;
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[21]  <= 1'b0;
            Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[0]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[1]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[2]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[3]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[4]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[5]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[6]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[7]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[8]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[9]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[10]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[11]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[12]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[13]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[14]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[15]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[16]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[17]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[18]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[19]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[20]  <= 1'b0;
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[21]  <= 1'b0;
            I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[0]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[1]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[2]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[3]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[4]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[5]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[6]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[7]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[8]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[9]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[10]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[11]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[12]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[13]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[14]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[15]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[16]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[17]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[18]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[19]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[20]  <= 1'b0;
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[21]  <= 1'b0;
            Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[0]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[1]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[2]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[3]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[4]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[5]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[6]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[7]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[8]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[9]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[10]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[11]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[12]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[13]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[14]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[15]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[16]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[17]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[18]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[19]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[20]  <= 1'b0;
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[21]  <= 1'b0;
            I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[0]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[1]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[2]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[3]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[4]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[5]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[6]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[7]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[8]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[9]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[10]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[11]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[12]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[13]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[14]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[15]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[16]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[17]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[18]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[19]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[20]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[21]  <= 1'b0;
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[22]  <= 1'b0;
            If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[0]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[1]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[2]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[3]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[4]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[5]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[6]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[7]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[8]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[9]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[10]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[11]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[12]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[13]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[14]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[15]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[16]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[17]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[18]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[19]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[20]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[21]  <= 1'b0;
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[22]  <= 1'b0;
            Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[0]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[1]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[2]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[3]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[4]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[5]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[6]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[7]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[8]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[9]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[10]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[11]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[12]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[13]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[14]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[15]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[16]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[17]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[18]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[19]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[20]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[21]  <= 1'b0;
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[22]  <= 1'b0;
            If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[0]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[1]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[2]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[3]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[4]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[5]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[6]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[7]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[8]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[9]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[10]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[11]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[12]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[13]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[14]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[15]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[16]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[16]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[17]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[17]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[18]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[18]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[19]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[19]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[20]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[20]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[21]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[21]  <= 1'b0;
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[22]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[22]  <= 1'b0;
            I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[0]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[1]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[2]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[3]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[4]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[5]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[6]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[7]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[8]  <= 1'b0;
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[9]  <= 1'b0;
            Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[0]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[1]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[2]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[3]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[4]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[5]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[6]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[7]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[8]  <= 1'b0;
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[9]  <= 1'b0;
            I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[0]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[1]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[2]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[3]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[4]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[5]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[6]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[7]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[8]  <= 1'b0;
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[9]  <= 1'b0;
            I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[0]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[1]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[2]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[3]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[4]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[5]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[6]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[7]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[8]  <= 1'b0;
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[9]  <= 1'b0;
            I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[0]  <= 1'b0;
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[1]  <= 1'b0;
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[2]  <= 1'b0;
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[3]  <= 1'b0;
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[4]  <= 1'b0;
            I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[0]  <= 1'b0;
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[1]  <= 1'b0;
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[2]  <= 1'b0;
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[3]  <= 1'b0;
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[4]  <= 1'b0;
            Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[0]  <= 1'b0;
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[1]  <= 1'b0;
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[2]  <= 1'b0;
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[3]  <= 1'b0;
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[4]  <= 1'b0;
            Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[0]  <= 1'b0;
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[1]  <= 1'b0;
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[2]  <= 1'b0;
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[3]  <= 1'b0;
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[4]  <= 1'b0;
            I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[0]  <= 1'b0;
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[1]  <= 1'b0;
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[2]  <= 1'b0;
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[3]  <= 1'b0;
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[4]  <= 1'b0;
            I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[0]  <= 1'b0;
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[1]  <= 1'b0;
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[2]  <= 1'b0;
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[3]  <= 1'b0;
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[4]  <= 1'b0;
            I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[0]  <= 1'b0;
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[1]  <= 1'b0;
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[2]  <= 1'b0;
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[3]  <= 1'b0;
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[4]  <= 1'b0;
            If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[0]  <= 1'b0;
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[1]  <= 1'b0;
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[2]  <= 1'b0;
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[3]  <= 1'b0;
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[4]  <= 1'b0;
            Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[0]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[1]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[2]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[3]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[4]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[5]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[6]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[7]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[8]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[9]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[10]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[11]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[12]  <= 1'b0;
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[13]  <= 1'b0;
            I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[0]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[1]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[2]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[3]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[4]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[5]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[6]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[7]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[8]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[9]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[10]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[11]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[12]  <= 1'b0;
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[13]  <= 1'b0;
            I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[0]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[1]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[2]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[3]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[4]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[5]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[6]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[7]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[8]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[9]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[10]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[11]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[12]  <= 1'b0;
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[13]  <= 1'b0;
            I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[0]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[1]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[2]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[3]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[4]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[5]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[6]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[7]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[8]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[9]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[10]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[11]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[12]  <= 1'b0;
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[13]  <= 1'b0;
            I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[0]  <= 1'b0;
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[1]  <= 1'b0;
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[2]  <= 1'b0;
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[3]  <= 1'b0;
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[4]  <= 1'b0;
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[5]  <= 1'b0;
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[6]  <= 1'b0;
            I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[0]  <= 1'b0;
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[1]  <= 1'b0;
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[2]  <= 1'b0;
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[3]  <= 1'b0;
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[4]  <= 1'b0;
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[5]  <= 1'b0;
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[6]  <= 1'b0;
            I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[0]  <= 1'b0;
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[1]  <= 1'b0;
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[2]  <= 1'b0;
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[3]  <= 1'b0;
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[4]  <= 1'b0;
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[5]  <= 1'b0;
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[6]  <= 1'b0;
            Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[0]  <= 1'b0;
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[1]  <= 1'b0;
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[2]  <= 1'b0;
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[3]  <= 1'b0;
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[4]  <= 1'b0;
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[5]  <= 1'b0;
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[6]  <= 1'b0;
            I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[0]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[1]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[2]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[3]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[4]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[5]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[6]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[7]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[8]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[9]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[10]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[11]  <= 1'b0;
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[12]  <= 1'b0;
            I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[0]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[1]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[2]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[3]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[4]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[5]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[6]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[7]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[8]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[9]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[10]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[11]  <= 1'b0;
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[12]  <= 1'b0;
            I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[0]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[1]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[2]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[3]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[4]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[5]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[6]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[7]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[8]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[9]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[10]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[11]  <= 1'b0;
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[12]  <= 1'b0;
            I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[0]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[1]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[2]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[3]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[4]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[5]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[6]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[7]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[8]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[9]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[10]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[11]  <= 1'b0;
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[12]  <= 1'b0;
            I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[0]  <= 1'b0;
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[1]  <= 1'b0;
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[2]  <= 1'b0;
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[3]  <= 1'b0;
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[4]  <= 1'b0;
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[5]  <= 1'b0;
            Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[0]  <= 1'b0;
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[1]  <= 1'b0;
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[2]  <= 1'b0;
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[3]  <= 1'b0;
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[4]  <= 1'b0;
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[5]  <= 1'b0;
            I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[0]  <= 1'b0;
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[1]  <= 1'b0;
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[2]  <= 1'b0;
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[3]  <= 1'b0;
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[4]  <= 1'b0;
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[5]  <= 1'b0;
            I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[0]  <= 1'b0;
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[1]  <= 1'b0;
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[2]  <= 1'b0;
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[3]  <= 1'b0;
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[4]  <= 1'b0;
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[5]  <= 1'b0;
            I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[0]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[1]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[2]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[3]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[4]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[5]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[6]  <= 1'b0;
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[7]  <= 1'b0;
            If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[0]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[1]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[2]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[3]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[4]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[5]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[6]  <= 1'b0;
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[7]  <= 1'b0;
            Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[0]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[1]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[2]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[3]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[4]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[5]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[6]  <= 1'b0;
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[7]  <= 1'b0;
            I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[0]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[1]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[2]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[3]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[4]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[5]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[6]  <= 1'b0;
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[7]  <= 1'b0;
            Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[0]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[1]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[2]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[3]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[4]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[5]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[6]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[7]  <= 1'b0;
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[8]  <= 1'b0;
            I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[0]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[1]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[2]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[3]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[4]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[5]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[6]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[7]  <= 1'b0;
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[8]  <= 1'b0;
            I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[0]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[1]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[2]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[3]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[4]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[5]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[6]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[7]  <= 1'b0;
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[8]  <= 1'b0;
            Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[0]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[1]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[2]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[3]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[4]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[5]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[6]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[7]  <= 1'b0;
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[8]  <= 1'b0;
            I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[0]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[1]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[2]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[3]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[4]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[5]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[6]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[7]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[8]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[9]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[10]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[11]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[12]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[13]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[14]  <= 1'b0;
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[15]  <= 1'b0;
            I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[0]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[1]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[2]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[3]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[4]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[5]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[6]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[7]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[8]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[9]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[10]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[11]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[12]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[13]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[14]  <= 1'b0;
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[15]  <= 1'b0;
            Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[0]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[1]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[2]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[3]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[4]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[5]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[6]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[7]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[8]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[9]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[10]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[11]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[12]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[13]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[14]  <= 1'b0;
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[15]  <= 1'b0;
            I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[0]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[1]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[2]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[3]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[4]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[5]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[6]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[7]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[8]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[9]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[10]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[11]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[12]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[12]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[13]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[13]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[14]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[14]  <= 1'b0;
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[15]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[15]  <= 1'b0;
            I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[0]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[1]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[2]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[3]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[4]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[5]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[6]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[7]  <= 1'b0;
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[8]  <= 1'b0;
            I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[0]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[1]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[2]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[3]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[4]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[5]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[6]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[7]  <= 1'b0;
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[8]  <= 1'b0;
            I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[0]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[1]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[2]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[3]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[4]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[5]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[6]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[7]  <= 1'b0;
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[8]  <= 1'b0;
            Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[0]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[1]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[2]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[3]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[4]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[5]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[6]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[7]  <= 1'b0;
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[8]  <= 1'b0;
            I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[0]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[1]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[2]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[3]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[4]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[5]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[6]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[7]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[8]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[9]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[10]  <= 1'b0;
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[11]  <= 1'b0;
            I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[0]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[1]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[2]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[3]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[4]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[5]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[6]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[7]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[8]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[9]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[10]  <= 1'b0;
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[11]  <= 1'b0;
            I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[0]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[1]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[2]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[3]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[4]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[5]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[6]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[7]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[8]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[9]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[10]  <= 1'b0;
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[11]  <= 1'b0;
            I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[0]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[1]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[1]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[2]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[2]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[3]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[3]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[4]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[4]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[5]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[5]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[6]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[6]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[7]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[7]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[8]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[8]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[9]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[9]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[10]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[10]  <= 1'b0;
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[11]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[11]  <= 1'b0;
            I7689b1f287170d28fc72712f5ff2fd209108b000a63e268b12da08dfed6d60b0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9aea0703810e5cd52352d3b0ede17aa0ccb943f1e0507585e4cccd0d0c427e98[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iea53e5522afe762dd4185f0262512abbb94b905893974c13e954df5553942b1d[0]  <= 1'b0;
            Ic114200c11d550dcee2bd668ffd91dbdd193a00571dda2d6f99b4985ef999f83                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I42c6c1d7cfb81335f01807b1d1c6b77c109482d338e81eda1ed174f739a6bf1b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If481e9fd41cf8181d432f397381b8376d9da7ddfba17b52e65e301e74c3b9b0d[0]  <= 1'b0;
            I2090cbe74e266e4385d5075f2913013cc38b26c5332d982cabead5dbe52d7775                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I839de42c6f3369ef5c6200c12baee8c9e698b3108fd6dcd58a71351d9bedae54[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If2e4ac195be838db9dd7b062319aba299887896862f1a340013226fa025b18fc[0]  <= 1'b0;
            I7802f219761d40fb4b24650bdbbc6faea69cf01618fbddae575028e96aa7c627                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0a1e88a592eeec68c060dd84ca2d75809b8fd80dd97a01a8d12cd9869bf94532[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I40914301545dfe0b6673f76e0dc0d1ab3968ca3b18fe8f4ff63d5623c31bafa7[0]  <= 1'b0;
            I9e11bb32c337ed1d87274c3040deee6d8813fd3f6795de87aeab9f93686ee409                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9114e17d37b4346674c23a6ef3a2aee35426292fbf73d7f30c895090bb749034[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Idf30e1a70a723113d32f621f0375dd85270da2f7386cff5ef4ff88cfca78b848[0]  <= 1'b0;
            I08382faacfb31fa012c97cbde6527792abbdf2c9124d886540d385dbf39e24a7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ife5225eb20e50e3cc959d9080f6faa318b4977bc9d04a67414a6cdf16c98e295[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic246bc24fb918b7c4a32727a332df57bfb205adc05150ae8d944a77cbdc62822[0]  <= 1'b0;
            I5c8ffe997fea9d77126fb36c6deb4f9b9c9b38e6aa562b574011ee5915a00857                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I28dfde2c443cd84194231fc87b8a1c6382ff3c2ff9b6d43e31e3a7116be41169[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6cac9957a16e7cfa8a125b40d8ce42cb7f502078a791b177d9bbe9589b612426[0]  <= 1'b0;
            I6f9b56f1fa7e83cc6acf75b74037938bcd08ba89ac2cb3dbf4df512fc9d521f8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I55da00c15261d3abb33c69ecc3f2090fb2bb3c29a3653fd999f6232982cf31ac[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iee4ad1e7709a56d53cd8b97f587f1f791fb88bf278fcfef32a29fa05247ca13d[0]  <= 1'b0;
            I3ea241ea179029fe0c486fead3909ff2c05b2d47e4484549d1d521a4f891a9a8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I05ca033870ef7adc8ce911a962bbd120591a1fe3b3044782b7e569e2b94ac629[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16a4499c48e5c24fd8a6d49ec3bf63c20c85f440c0c897cdb840e9f28fa2e68a[0]  <= 1'b0;
            I6f9fd1c4756d8d1250b0ed96355e2739d3bcdaa3603b7e1cb5cb0dd0ad5985e5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4ef4ed6e15f48f289815b7e00b2454a26e076b8dc9b8903e118507c9688e905d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibed209db0bc502e3fceb4ab86ac20a2ebf87c43391a546d592e5aa32709aa8bd[0]  <= 1'b0;
            If084c3e6863c87018f76e95d715c83cc83dd85ddf7664f98c6ff35e8a0ea40d9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I25e57b538f9a08a355a5ff8d26d94f81bbf2ebd0039881e74aec76ffb1dd48aa[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I05dc9e8db597a2123632b2934d864ae64cab5192401d8f66ebebd95618590ba2[0]  <= 1'b0;
            I7fcd9ade547e48c042200e4bae7d4699b326df8a285204b7e23eee2a019cb01d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I070ee6bd21603d58d3243ac556db2ca3c0476c64fde6d32aff54e0577b0472f0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib309786164a7d646c17533008b3aaf0fd86eda3c5ee167efc2080ef5b26a9ddf[0]  <= 1'b0;
            I9207b21b45d4265cc52ef02ed257ea78cc5a269d98165b2a7714a25b1c477521                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id2ede5f3d3ce0652bc9ceeadf1de91fb99234718893eea8cc1779cf900284e88[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id9bbd0f5c16ba0ffae6a0e5304e1726b97df06f06feaccbb1bbcaf0e01be3823[0]  <= 1'b0;
            I4322d4cf469c3caa560e48f6eb1fea264c42dd76b65977c24c676681518691f8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie251294e2cb883a913e91485cecfa90bbd107955ceb6d60d4a9b1808aaadb2d4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4294b001f220e009c2a65fbf8b36ce1d8961c317ae8ded31cbe5aa288191e009[0]  <= 1'b0;
            I924625bbe810db6c8d5cca4407571d5819d0f7361e2d7f1906bbeb822457aae4                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I983e8c64c323025590663edf53b0666d93d838f15879b5e3df245a8e9ac6fb80[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id1fe66d1340965020f513e73a4f77d18f4703c194c3954d40a7f1bc37fc1342b[0]  <= 1'b0;
            I3a01e4ea96fcd387a6bda68d7d07cd6b4e89ca653c798f08ac8402696b42a371                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I46e5ca785f6f4304dbc4fbbf3816d83106047f0eceea77717a1ad5c41a9ca441[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie95c9af987f352eca30c8546d306af7cdada8d2a8037200d303e6afbd5a4f448[0]  <= 1'b0;
            I96114d8145aafde7f8f5666ca2f6dcea9ddfe9796f2e3a54556fb1b23fb1a331                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibefeb67be2754ad6b9a6cda09c66529a7ca51536f5c6ca6b05e6ac1de34ae514[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id34d005cdd89bf304f95101c6fbfdd40d6c0b1742b5f3bee3bf043bf88c3d063[0]  <= 1'b0;
            I006672e4b2c9c693fe5b05655ebb6f31e96ca8e2c92eb488cd28e5a940e49766                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0dd45b65c82498edff9ac44b5b07ed30818dc1ea2af48e5c1394466865f36adf[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I79d61ad4114817a49b1dc8e9314d9e3be9758d861974ead362ff0ac862d1d77f[0]  <= 1'b0;
            I408f22a4a77906024a2e6ceb970b39ba9ca76300fb2584bff35e37da452c6613                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ica92be8c7303e09b9f549ec558e655816c1d23a39b8d5324060f64a391984c1b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icfe1fffea36cf64044389903be9550fe283d4dbb7f1b47aff2005e70765a6045[0]  <= 1'b0;
            Ie84e7eb709edc06e55ae27284cb93a0c656ce8559679c49a47c7f03f0d64fce2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I726b6a7ed2ab76b049762263a08d5121a597f30ce25a6880b51d6b01aff801d7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib08cf17b2065d04f587d1a8231ec1e4bbb6b2b15819de8a7efe18b477515ccf8[0]  <= 1'b0;
            I84fb24aeaf533382e57c00dd73683ce0e4f5f33a0e7a3b36f2ab00732891682f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I89362accf0644c192f06b113020d2071f1389e8ddd8d4fee492205db15b25b66[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I21832b7270210e1bb6a23930ad9ced36d3da201d80310263e26eb96bebd23612[0]  <= 1'b0;
            Ifc8b49d8467101e2eedcab4b6ad6a73e4f657c0e995ccaee5dee276a5ae916b2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4473c0cfd2d569bc671ba814a524058946271eb49a04fc384e9373185e1f4a6b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5dcc76c47f3c9129431152fa6f7047be203fc556198b45db15a9991647bb8c85[0]  <= 1'b0;
            I001fd8ecbe068f57df7498db3f519cbb5a65bc5af187f1d34b5eab3df45447d9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2ba73f603d9cb767572f2b2f2a9732e2ebc066392aa85888df87da4dd8b84113[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I450f5b0f5d2b96636ae010048040ebd744fc4ca164cd764bb33615741ecaa62f[0]  <= 1'b0;
            I11745815606a2dcec9059a24625e93a31b0f15d9b81c97403905e00d3fd64f43                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I82f10eef14d4ad82b1f7f8c5d056c398386a6cf790095113a615a8bb6cfba233[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I35d64df6881fde0d4836aa408258db7cc1bfb2f066abf8c9345670b78c466b9e[0]  <= 1'b0;
            I37a341bca6a12362e49dae8435798cd8e7550a16cd506a7f852f4223088bdb4d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2fd5dd69a5f551c26d9970d09ab0e26ac5183a0022af58e2bec1dd1efefb139c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I11944fb91fa1b1d5f076cc36db77f0f8434f0edbb1236c7a9bcb45f79432ea9f[0]  <= 1'b0;
            I8ab2f0a2c9cf1f1e0401a67f3749b106fac7d45293bb9648325f330e3230517e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2fd258374a5bda5c58c1fdc6e305789a598fbe70657d6dc18e8878b6c2b0441a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I49642204473312df5a3bcab2692aa7558f44f21416226675a4ec10b0543cc5e9[0]  <= 1'b0;
            Ic6ce7ef3f9390c17ef23e718bce985f168504ddff0d66e2babddf08b37dd2819                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I76942d3b012aef2097112a1c1adfa2bf986414df19a633b87d2f3c2a61d27351[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I24e0d361a2679430549932a968d7cc25f980275fea5554e3453ed0a652d31caa[0]  <= 1'b0;
            I26c16ba52eb0f661ca599263265d1d0d7e1f155b4afec85407f3ece6fff3c391                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ida428d199205588ecd8cc963ceb39e24bf6f2d004b675f3cb883960e0f089842[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I386015f8daacd2ac9cfed376d3418b56ac13f075a43dde939e4056c29565a926[0]  <= 1'b0;
            I31afedbc324d4ddcd04b3ef766154a6414cc6e31eedb0ff24b40698430e84927                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I91f0247d07693c53d716345c810ffa0ee8d3f4b793ca8831763f5465db649c89[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I32832b039ae7e6f4b1e38cfdf680e5044e383b921a76189054511ebe5b8c0d7c[0]  <= 1'b0;
            I807fdac75cca555b8d81d1b4d7e53ae7cfa0e4b83bcb260cadae218faed4f781                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I754c4c2dda64bb938ac60db8cd469c6f3ee0831a3a6b6b98e902c1b72663ff28[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I09fff9b84a38f3d19685f9627d01a7183cf65d72110802f11e8da0e01194bf88[0]  <= 1'b0;
            I0f8a9c8deb02bf990a6ac2ac0569f9d0ad9f167d7c18dc70ba544912aed4bf78                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I567c2801d5598a057d5773ea5045f594de038bab88d554ad2c713cf56ef632b4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib82c65f09934744abbba984b6e375bd69ce7231a5085bb00ba4e673cfd3aba38[0]  <= 1'b0;
            Ib3e6663aab02fdb649843c552944b6e325240f5010acb414c311ae56e78f8459                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic9f57a4a1184139b219a3a5e3c554705469b79d3ab175ddc74512ccbfd5898b0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8ec5727130bf67c04580aa1b5b46cdf964db65750f2fc9ce55025b1c117b2bef[0]  <= 1'b0;
            I41339bac55a76a05186d632423b1fef8173940f0cbddfb64c83282af5cd04cf6                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2dc38e534505cf47f391eb9f4b090e16136d12619b4fe91cc8029bb5a050689d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I862dddc300df692e8bbf4ca45a24d840e51ac1e975631cf4ebb8337ceefc2eb1[0]  <= 1'b0;
            I28fb4df9f762474ad496e8689f21d13bcc5bd4fd79190892b78409a06720e2f3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib83aabc196c7633dfb4a9bcb4b8d06959130620de297f9dff77b1454a8f2f96d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id08a37df0c5095196e2d760938c4d0b7e8716c25b55d9a9656d86c2c473f9c2f[0]  <= 1'b0;
            I84ce9c6711b257cb8cf2f09bcc02e0f03490605e543ba12942207df6fabed5ac                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia23743e423f143b75923bc7b1a4363323d46ace080c8ee9d15ff687afd4bef65[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I40204cd18eb803f82fc3ef933553c6ec41331f6d4a15538c287b8f57adebb89e[0]  <= 1'b0;
            I8f3d31b6843ca54e80e8f61be651cb7788b43302b001d791357fad349785eb1d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id49eabe82a09acf1b3a3aa3be9bfbc0ff958b96b44ada842e892c587fbddb8fc[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I677f733f4e801d99dc2fd1987683a7ac6c8609d84da6c95b8a7056ce07845665[0]  <= 1'b0;
            I6fb6112b591f6f1495935e422361833f041f7231996d88a3936b5da186e4c48d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I93584fe5ab7128b24b2372bfeea00f7a2bf09d50b1fb535d01cc141c6d6fc377[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifeb10787a88bae5943b616e3bf751faff5e7eea80e45e24d60a760f4d6b0154c[0]  <= 1'b0;
            I959de6064e6c31bf0d18c2d6b4c274ebd5e9fadd996fcb32e695047831716951                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I44142c70d3ba4660f5b85d895710afc623ed3470ba85eab3dee5e49a59e1b124[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iecc97eedc286cd1c3d301e35036e81a10d164d59da9252a92ca5f355a828367b[0]  <= 1'b0;
            I0f46fb1c05f0f882ae878e86285077da38a459201c305e13fb4925ba34eaef8e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id8b538e6a6c4a147c7000388923f1d89a193f8ec53ef214556e005218d2c240e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia9a21e6f22a6cc828e041980ab142b418938a92bf8e868216402a46b8c614a19[0]  <= 1'b0;
            I99e249a8eaee9127d347ab629dc27a21d5b55d2826c354eaffd9e6fec47b1043                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I658f9399a929745b4ba467a1e019fdbe214acd543dd4f5f51a95292420281401[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I355f4f82732333ae56692d1c7ee89b368d938d9ce1d5f806be7e46482c10e19c[0]  <= 1'b0;
            I2f779bcb2996facec77594ce5efd7c78acaa443f2b6ab3a5506ae96dcb986b23                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id1ba70174cf019078c719d1d50a82a61fbfdeea2a13e21a1247e567b9266365f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9b2ce64b97ca55921bacb9b6aa4cdc8da5c1e33db4215a2470b7cfab3693576c[0]  <= 1'b0;
            Ia765277dd8a5fbb2a65aedce2934fd6c4dc9daa4e0b316604f6f137f19fd5d25                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I797dfd66b521bd680024b6e46455d624aa58b4271f5e6ca19fc7abf520f26222[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2d78ac4a4125ec25a02df6484c0ae640a37f915383b72f33b91e87cdf376fdf7[0]  <= 1'b0;
            I1a47d1294e98ebbb0493fe3cf7743d1932eac70fe9d2754367a51d9a49448d12                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I74f49d84817f2467b8ccdf03acbd7372c58f1a4fddcce45cb882431b2be20b39[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id727bdc545af53e8f89be0ac5627d0c0c0f0bd7d75030bcb41f198a4fe9c7d64[0]  <= 1'b0;
            I71c11e07942c42d17f5b85b1da8857e91f789966944c1e0948bf5f0285c91079                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib756dd9d8d9a5233fcd368ffa91f5d7d9c8825b01bc26140e5a717d3ce263e64[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7661c17a1c73dbca82a6d3bfba2ab85ebb0131c1e513f093e1b0aec54907595d[0]  <= 1'b0;
            Id810b154e951f2b2d0b8ae826f31effa4f39b3a0396d446ebcceedd7225c5018                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1bb2be29dd44258b24a36ad9b1625ead1cf965856f1d9695c62ae80de142169d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I553a83634252c50164bdde3576d7e1552a147490d02eac6dfd1140a46b813d08[0]  <= 1'b0;
            I2a96d9fee197ec3bcdd50abe43ee0d3992f5b03db5cdc958771ed812bf3a0b4e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icbff209e6c8353c58f46c0688f06da0cdf71a95defd8937f2d52d63d387d74b5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib450c1ee41d04516060a410bbdfb605f0ce13cd8781596ce5218928ed207de8a[0]  <= 1'b0;
            I280a4a7c5231cbfe245c071a856f7d1560c4154e9f9a4c5fb6895baa2f4f5871                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia628bc749f04b3d12509effbd4e0bc5ac0fadf48a2cd5663e4c2094593870a42[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ica745abd4de790f1cd3e2a5a32a9d0b5edf1b64e85759c49f3b4e51779443709[0]  <= 1'b0;
            I01562027a6c7a542ae356bb1d0db0dc55b2094f3470a1894e67a3b7fee9e4361                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5ac2c7b61022af9bd2550f824b8e129ca1c336b1ff900b0af785d86e33cf3358[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6399b29558311ea40cda1388848ce13bb7593bfed01ca2a10fa5d8ed6700df56[0]  <= 1'b0;
            Ie3eb1aebcdf48fc8f41590f0e9524e989193fd14fae379a200c20d1fd3755db3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie511320217185f90f1e4a23ab51ae9686801b09657c714a5bdd9c4e26f070bff[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6f529a4dd77f75d9af4350baf53ba61c1e9c5ea6227c26690987d244dfe71528[0]  <= 1'b0;
            Ic585c7a7014e8bff08f28b2d432e9783bea57ff5b456d851503a2c3eee80a768                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I032b833c683eaf0c1c4c60ad831278ab0ed11ed856361be3be59dae656141fb0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7a94e46f1351801c2edf76bf3b70e3b5100b8e6108d60d9341591aa59f4e95d1[0]  <= 1'b0;
            I4f0a460fa116f5a45cd0c435e594ccc7597b449cf5205391a2dc6e977f4bdeb1                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib41d86b318a3004b648c9a1b0ad00bbb144511fd63b1c7648cf3ccfb996686d3[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I0b761d71a88d70e6228dcf7325206f840d9da85892ba151c317e06079291fc2e[0]  <= 1'b0;
            Ib7f3bef766d8e66cc9002dbcf3538dbe974b70de4d7a8a3d9cc3bfbe815841d5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icc4bebb1db4145f9cce0fd4c250f7501f300b6cde1f31327d80b844adeeca1c7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic2ae521a3a6fef956f28a89da365b0838d535c9f7801a405cf60cc776ba0af2a[0]  <= 1'b0;
            I027d6136f1b64e5e2f94af338f8fbc0ef9fdf8dd0a2d58aa0eb6879557361681                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Idead9dbad4283dce602c05f81e98610ab7f65f9911342174ceff7c95dfa9ddb0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I01d9f8a8900be1981c601c0ccb45c1f39a0fdc16179245d80fbb2ad6d7060899[0]  <= 1'b0;
            Ic62f1d181b6452f30ab2146b4e43113b2ca1bf21962f686be46f59084d39fa0e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If7060467d2fac9aee8d69c5ebdc24d515a657bedea3da55d13ed6ed4e3c8e79b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icdfc2f0ce24f01af7df8a99b58de3a74e1dda0eea5b41ff2c342106cb226abdc[0]  <= 1'b0;
            Iecddbb8ccabf830117fa8836a6eafc8dda6fa463d9c907ea25d298249bd066dc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6aefe769159bdc69fee8e09e46357993c13dd8ec9f059cd51d43944ecd7ce3ff[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I929ef5474f10c76c4686fb044b2833b6ba1571f2e1c82b6d92cfaadfa44946e6[0]  <= 1'b0;
            I5a2b6e5bff0ffadb36a7f02dbb3cf48ffd37e6e29ef09200db12ccf9fa9d8450                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icac3a5cc88034cf8211c158a1bee2a04c228afd4eace1b50c7460ad5331ae02d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I55312932ff9d69c8ffa1e42efdb5e775ccb21a8f9e8791b080b67654462e537a[0]  <= 1'b0;
            I3a9d955359963dadbc16853d82bc2495f84c37d8cabb868a144c5f24d9edb2c9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ifa5d23491b028cbdcfd79fdea2e0784f068c1fd381dda7ebfb5d457800e510cd[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Icbdbaf4eb2f30bb78db34a582e06dc91689b9eab2f8fdfe4fbfb41a8cce93ca5[0]  <= 1'b0;
            Idaf457dba6ceb8f056ac34d3bd84bb9e9554c0d55db8928b9b48692c316e6fc5                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic27b23bf87ceb2ec2d6460321286d798980f966c89d0f8ea42a79a0549b2128e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ifa4cbbd5c3ab5e47a7d5135e4dbaf365e79c4c6a806bfae88c9c0e1c9ffe2fa5[0]  <= 1'b0;
            Iec8531839aeb35f1c356e474abfc871d1ce889c4aaee1b37b272dd9650fb6981                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I01500dbf2528609729acf26a24c11bab0adf8cdbc0633527f21644816cfa0dc0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2341907334935e19ef0e392216e39bb35c215730c464a85c0e1b804b364b492c[0]  <= 1'b0;
            I6a320bd601e721d94d7ac0aeb59e2c81a0a9737d2f7b49d668369336dec2ebfe                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6db96717b6fe00f1f87347adf69ce2d4b4464faa472ca989bb272b36454e868b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic0bbaf8314688690b5a15a5613ab149f604a8bfb92a2b9ed014e7ce2757d0743[0]  <= 1'b0;
            Icd9be4d5172c268eba385d2cf858caf3450d81a87bb90fde24fccae0d1637d99                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia8cd57b3b123e08e2bc00f82da941eb4431cc816928254135dd13ef52eb9c03a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I19ff0bebf62a994a2b5814ea41289f72cd62a38d2f37dc0027beb0f488926d4f[0]  <= 1'b0;
            I64227cc72d5c6450ebded626fdcdfd149c8e29dcd6839ad76b2b9a932817fdf0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4fa8db615d84b02196afb2ad926769bcbfffb7c81170387b4d460c7403f0dfab[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4f9435bbcce379d6d591547481382ab188003b97877c0f32462ef9e33aa8bc1a[0]  <= 1'b0;
            Ic754b281b704937ea08e702dcb74b7175f8901b29809052424f867a6685c1d41                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie81813a1836449254acfcf7674552545d2cbc852ee2bd2f37378345ccdfc61b4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9e497e3ee797c274b82ecca58218c47f9b663bcac21b1431b45c17d5e54e5a4a[0]  <= 1'b0;
            I861b39dacbc8ae1c9cb21a407a53608f0d5adf148148ddb8c3ab1cbce25e2497                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id9fde3ad430d66c92a5aa6797b76ce147e39e4245ea761e36d81214e7a02b4d8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib929181cef39d751d2726a054cd0478d309e58350ecd11d3363ecba8bd4cb7fa[0]  <= 1'b0;
            I994137ceebfa9f1bfb6f3342c02ef25b1a5e881f6fcf6c2e7f274663b5b4a3ba                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8f2cae5483691fdf6ea64a4ccb2372967aa676835ffd4f562269bac888840d17[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I64fa7f4fa09b7909840d8edb83f29f6a2379419e65b80f592b37d8ea00e59475[0]  <= 1'b0;
            I5193db4e129f33dd7cd8691b74f52f030a066b583bbe2d9a4a6e9962f1c43280                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icd8572ba29de1a399bc077f53730492f4e89deb95b9136608da0d029ba60ddd1[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I35beac843abd6268c39acb691d3105a5c386f05461bca8c63b951ce1c2ed07bc[0]  <= 1'b0;
            Iecd0fbf7643812e36e8d17ed6782ecf4b181df9d284988b1f416de07cdfe6095                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6eab6bb656dc82d656eea6da9dea574b230f56c6ab898a7f80973183896d8347[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9d8fbde44d35c50f5f24ceae6f2e16ca2f280573caeb8a3021b6f69dec3d04b4[0]  <= 1'b0;
            I390b2f0e16e0de51443f9cbf8ae301009d17581f5e20ec4956a8e95ede2c0822                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Id802e388c3b33f7d0a0960e0e51da02e7128da423d518a916f761a16b73c17d7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I507d851a78a765c18af6d529292384fb4cbb06cfec0e22d516adc79b8ea13c7f[0]  <= 1'b0;
            Ia733b3c17807a98828719894627b0a1fb161ffee86fb28c11d92f5b185a6284e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I47507e717446a9ca85cec7e5fa382cfe435affddcbf5b25d4e74f23a143b02b0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I80fb8d450dd144ffade989cc2cec363cf6bbcdc267f5372163fde38313387499[0]  <= 1'b0;
            I6b87b44befe3363656697619cf3dd967526646ced0f90813c24c960ad4d57d5f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0d76ba051f3db8c1efd9a8f0bd0ca77cb28c7dfd68cf4c290ab00edfedb15237[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7844074cddcce1b95a010729a9e4ce2bfc4f7e1962b84af0e0a3cbb2c2c08206[0]  <= 1'b0;
            I29ee4a3cefb214cdfe60e6907e63799323eec92930d4a48797c96a7c1f3e3a15                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I39dc59000bb2e3fcdebec08ddd22a460fad0c09e8b68adc7e72a6e4c3025da49[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I88be0c0499713ce396832a79853e9918ecdfed2519fba6fd7c0bae51450478e7[0]  <= 1'b0;
            I748cf7beef2ac47341c77503d0042b6e1570248031f1d9880d0bf14969378379                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6db1df05e1ea3d8011bbd6e08c9d50d91e672a20aa2448167343b839e8f6f888[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib585733bf4c3eb59a772866965420fc7397b01272410cdb701f289daf9549fc9[0]  <= 1'b0;
            I559b90a32f7cfdeb35bcf30683787c6357460614330553ffd4f5732cc03507ed                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I0d11d2b76d26d33ebe0c7577f5d7bc68ab8f4840deb765b17f4f7fde0a4b2fae[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ida673298c761bab46fb26d4e73caa99f5b3ade7f924d99fcedae4e47c70b5b67[0]  <= 1'b0;
            Ie6d770decdaac3d75cd6c9eba7edc89898bd152a7c75f43a464a47c9994c9a87                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ifbbf33f600185eab85dd2c0dc5ab2f5e0e2cce52373cc2acf5e466a2e27ded58[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I60bb81cc7cd9a6212f7b4261a21655accd6cd09e7aaf5f78f7f1f4dec0e8489b[0]  <= 1'b0;
            I6541e01880f3c658b3404a81e96fd03b861ba4a26ec927e9c2c64aa9973dafc2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia38b628fe0740039fd44aa0a75c751e1a9e176bfc305a978377c1fc9525c00e4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I85d3c885ce504524ab43daed7bbcb599cd7e5d6d3635cf46e278345134e97e22[0]  <= 1'b0;
            I184fea1e133f0a5b9b8a88926ebceffbb79cf7816941eaf9a326764d876c924f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Iaeb5b860946e41cde629a762ab6e6ea4a0f177083c9ac84d90ca99fcb90e7c9a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iaa08a49e0ca4f92f38c7f4d115ae1b275e45c42dfa6fd4b6a2ff40536b7f5f15[0]  <= 1'b0;
            I78d3ad872172f1089358c601e00c98f526455a961f30bfd6a966e8d8bb6bd098                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibc0b2c21012904530a727f0c5643b5187d7bb8706a308bdd0de67a80147db974[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I197b3231cb1da107c5001075809e9fa75e4089871d473490981a8b44d3ff5e4c[0]  <= 1'b0;
            Ibe18bd1138dcd8295a35b807d811d5b05b07df9efd2326d0cae0cac6589e7bbb                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I008d6180d4774d2472158544239ee654e73570389873b54b695946cb78ddb7e8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I384c04b75344f97c691f70965d7e08266ab9cd8862e04ba73b502a0f36ac5ea7[0]  <= 1'b0;
            I68fb3ebbcbcaf18cb81eeae19529cbcf7fe4175df44bd847d87ba9675ffa862c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Idaea720265ed96d87e8852c36eebd63e2be5b9768c7803f13fe85e7532b75ea2[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibf95afb3941a2272d76cd7256d0789f11fb35a3020c3ccca5b099d335d4a2330[0]  <= 1'b0;
            Id2154e04af88ba8cccdbe100e1c4e4bccbffee35bebd3d43f9229d2915bc1deb                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia7bf8296bff6d2322977b0a31ba519bca04a1d6c6f6c0cb5a47e3408bdfac573[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I885622bb1c7371f4afa3e9966f870d2bf7750c2d2280a2a993a5bd9854187994[0]  <= 1'b0;
            Ic95be152c428a61c5e57fa5a5e776b9341efe9f2d08c73fe0a9d2663b0a974e0                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2a69131c92e4454ec846c7528679731db69a2aa63420f0f22289d5c0be743be9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I719a3e78d6a298f7db920bf7e355f6fca2c46135abb8ccd1cc3ea470912d05c1[0]  <= 1'b0;
            I6e7d06d6c6a765e6994847af070c889f9c7059754ed634122e0204f750919234                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia5fc094477d9d66d7fab491b73a00f50abec21827f63372fc1b7e0bd31ccf375[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1729b841d155c32b617727459f01aa9a9a6af56de5f464e20e900e3a4da30dba[0]  <= 1'b0;
            If0343bdeee565245554859329a0188f1267cab02c325fbe93d4df18606760025                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I41d88c1cdef0448f878686d88600bd254e722761979a244cb1d00724fc1d35d8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I96affe6d042e09b07278ae45744977fd3719a31fa5d578adaa2b3a66b2c3ebd0[0]  <= 1'b0;
            Ie090cc0a910baacb33f7e858eddac0b221b9a5c567ebde9bba44380b06e8dc29                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I85e825a905ae7dd292f400406048736ce90fa7d47b6dc5507254283662fc7564[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I12e1e01b28d2d443785fac1d0314b477b221b17b715f1153c5379a85b4b5e3aa[0]  <= 1'b0;
            Ia0e41f1ae6bbe04c95f97b4d03e31d86b4399463bbd9fb5bd714b9c2b58bb23f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I80cf17357df8073b050d80de366bbb919c5f6c8983ca87f6606a84df1b92c549[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie244ea5cb57e0b4c14c0c8c22592347d1389a6b0f53b821335b821ca5130ad6e[0]  <= 1'b0;
            If4a86cc5d7bf6b2552861b330822e6bf86fa60debb5d503d86e081b720f3432e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I68a074e808119d0f33d54d3863c907dd5d761b3f6b144b9283e67f956d5932ef[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5a07f349b1fd7d668d35583c50dfa3ceda070e5dc241bff1ecdddace6624bd57[0]  <= 1'b0;
            I0d2ad8151436f1c3336aae018a92e8bd400452c12972fef401e7ab55030d285b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4aab61ec97ec8dfc8da6d2ab5898bcdfdaebb0f024fea498a6ecbf0bd15fd1c5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6e5f194e3acb27a7fdd060e05aff00bb9fcd0904b3f920d7db0fee84c1534558[0]  <= 1'b0;
            Id2881f7fc5d7a68a4583d24b1a8a9e09928ea1e5e3ec22fff19d4d59e12a201e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I26395ccf79a44d582b559acac5845eae4a01464019f7739b7d52d8c8a4c11154[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I09780397509ca78f4b4aed5b08cf22d8eae797d1d1864cdba4a951ac8d583c91[0]  <= 1'b0;
            I8733749031c60ed31e2867dedeae4f9ddd4da169ff086c567288ece5da43decd                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie9c493e499f4b2aa598c54d5a5afdf39447612225daf7f9f5b3c2a23b5ee0ff0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iefcb9b5b2f238005d0f37bc519349bbbc130e3e072814ec48b4edf9c853a6913[0]  <= 1'b0;
            I9180b03e001160fe9a51818e7641c427a35e0b2cbeda9e6bc0e32878bca05815                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4368873c6f3e3d6ba5e7e83747fb90120e80de634655a9d2a97bbee88a9d8501[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9835f6f38580d8765566723f5a9adbfb4935af8bf719b3e4918e1b746cf12241[0]  <= 1'b0;
            I2f00eb344711414f5f6efe7eee64b5690b4610385673a7186711075eeb319cf9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I082b315a51a6a180909ea4f576a9a3c8b0550e64aa222610c2e6906ca78aebad[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2266ca44e019a30bb553f955a158a5b075035c4b20a0b3fca6a3675ec79b9997[0]  <= 1'b0;
            Iea8f3fa357088442ab8048febba14f1e6ae367c6b1a854ce0b2c4861c4a2ed27                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I23872b1af6db7e455f25a7ddcc050167bb10de0afd16973c0a90804349210372[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I684ec077e37638f022f10b5eb31403e6f9117a83a606f2a5013c2c33b8d1a8ab[0]  <= 1'b0;
            I0d3923859952e0ab6d926924645383b83904ee287f1783cdaa7f314b171f4171                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9796589e7a8535d47d56f792d80838aa402e3c235035b517765096d2a6843215[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9331428911b817ea45d1b5ae75eb3ee6e05c189785c995e5d2625f12ce4e0846[0]  <= 1'b0;
            I45f444d890e00116a19e16e3c50c555419e910e2413c0277f62032d6ff66ca15                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I46d39260d96216c08b7940ea3bfe542bdbd0966f5e798321bc90a2a00f64360f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7769e8ceb72790c37b351c32983860280aef172974d19a2e99348607863a97d4[0]  <= 1'b0;
            Ic67dc4f0898ca883d489eab901e11caae2adbe1c1c502ab57f5366cc26d4d335                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1033817563ce88e3b26188a88303cc6703f47afdaae4d5457fab8b73bade5274[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If09c36408407b246848b29df63e789fd1041815243beb4f27db0e774e853f1cd[0]  <= 1'b0;
            I89150482cc550af995633308cb14fc4aac6984b8c5bb09ed4018e5692f8866e4                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I343bc73eaaf00a82b2674c8cdfbbc5c6ea52d10fbb9e9453cf4fcf2421b97e47[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I533b63eedc528cb36abc0a469b66b144a6ae5122c038eef85d8d0557c3dff3ea[0]  <= 1'b0;
            Id4c7f10c8e46d38df8e36571905e342a0b283e8badd00d3e4081890010c25f34                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1af6f4d00567aa1e302e7d8830d761e7a9a616f5e4e958b264701c476216de4f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I051e3b709db2e7861d31165ec1e5ee679f1e6dffa5a951072831ce479c16f27f[0]  <= 1'b0;
            I3c6ebb6c57609827961bfb1e39059b0805cec40a48787adfc9b2b138a5012c9b                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1682f44d820722e2566b0d6c02fbf3dc72547221d519ed071e7c7d77728ba21e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2fa018ce903921d0a174a63dbbb29eea8d5700b376335b2ba9bd448e8782018a[0]  <= 1'b0;
            Ic8177ee86d033bd8ab95b63937a4f80b02ebbb66d4c16d84c8822d133e7cdd0d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If0095cd5e911c91331d2ef6ab3866101080b3cabe8d1ba9104b6b5ae5d18c713[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I36e06c1d77080ff75778f3dfa4ed60e66f9a3bedc39b214e3fdb5b6c21f1cd3e[0]  <= 1'b0;
            I65cdf21d7c52f9a1fd2d4bb265a678e8b543e0dedd9fdc5cf9e12ecf756e66ae                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If7f60dea1e83c3f86ff8ce3adda8214324b2064d06d69ca68477288522ad9de0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id647e3bd88fdc7a3642092d071f66f74657c8364937caf63c723f1e027c157bc[0]  <= 1'b0;
            Ib047d12eab2012f21895617ed9bff57a0678c2c85235301fa1276f99ecc8625f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I3b1abc53d350b3b39e60c3a5725e5a21632e7f0275988b98c1fdaeed5342f9c0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I015b73e7e4bc4c2a3073a304e58d24f5c8c32e90299f004bc0f75eb9e18e6d41[0]  <= 1'b0;
            I4864402239c958072b187da428e64688ab13cd5a3ba940785ac5086f81c50e92                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7943272afdae80761f8b673788c92e4461bf3de3229f7addec1e54743b11beca[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7c211cef6a581c5a6871d4c9a2b7ba29a9d05d36b0a758106e006caebfc592e5[0]  <= 1'b0;
            I8d03bb3beaf84d3f94a15648cd5536d5f14020daffea4160bbd12426018140e3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I8417f8f367de885ebb86571786bd964d4a81d6712a88c3a8071c08d13cc7cf58[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3f2014435aac47a3c807e9ad3f0829179f9285582b7ff2e3bae250a25e800aee[0]  <= 1'b0;
            Id3b64ab87f29683b9210364e13398a54c486d0b8b8a7a5ec6f15c29cf752b5cf                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I653822ee3643c81b817be0d9c3f682d0c806ae17dedb0cae5b1aa0ca914e6857[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib27fb4891a6edd486a99f23a750057de12a5a3e3fc6a5fad7976aa7e961e0c54[0]  <= 1'b0;
            I2f3b819fb1f865426e38d2b39a1a4a8ea0560e0888f19913e2393d416205f3b3                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ieb917f5db48f3d352eb252f6ce309bd972cab47f09ba1c140f66192b260f3925[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib58cd067e009a5f4b72af8cfb1e5c49c18f51a2ad8880f65aee683bf8ecd40ad[0]  <= 1'b0;
            I23e7ddde350dba3f41b08c523c29dae580b57e09b8fd9d35af6ba3bd4b104b6e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I313a01d9fe403e838310c49dc37a50b738025400e99faefbd9b8cbd426edcfaa[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I7e40bd6625b1d7deff82f67d46817c7af70f1da57561ab528b553b3d244b3f1d[0]  <= 1'b0;
            Ifbd6430f8434621a650f4942f3be3669bfaa802cd912188e4139542d2a64a511                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1b81a8a827bd2222ea6820d80d13e537868e0157970625d628f0c062733ec3d4[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I01949f24f74578cb63dd095e8ce639ce0d273c14da81e75d00097535e391aa4c[0]  <= 1'b0;
            I1cb9b876fadc25322c3f466b101084a68e5a283260303beb238d55ca788523c7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5615438871373f7ad838fb5e8c24b9517fb94ecf6627c803e66a78f778fe9c42[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id8f2a0d3524b27621ca5a576bf16e15789e6257060225da04da2a5fcc8cf751e[0]  <= 1'b0;
            I9bd2fc6de34fc3d410b3d5e30c2e9e811c7063afaa6888afd119cdc02e39afae                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I07f9ecb15d2696b2cacc35c935b497b2f8cedc55e2a661fa57f2d0783e6a1001[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6020dcffd9e047c03740cffcdfe790eaf614ea1036a50fefcec9e13e5b5ac4bc[0]  <= 1'b0;
            I9e9c82e0f8d919f8e2e03046a1654698592da05002140ff69fdd551598618d59                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7fbeac90b85dfc78e20281021fc1d7cc90f9deacb2091ab55ed07f51fbdbcc11[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I815f772d86db329f78fa75c3326c129ccf0f6c5f383b42ef18033e48d11525d2[0]  <= 1'b0;
            Ic9fded9a702f4299431ec45bc00c9111907d62279133f1a5f62e5f6527823aaf                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I46dfb75396740f84b7758552420a7ba8693bb1ca5259a67530c588585de1c337[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2c8a33831a21c4c21dd58a300467abcc82d52e7636a73a12a003a4144d43e0dc[0]  <= 1'b0;
            Ib95adef89f659c6d98e43f4a9c43340a0acdf273ea6bfea0b8e99f0751c250e2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I60e36bd866a477c35110e2688e7fbb13b0303d210e014c9e151b313d130101a8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I8c7b9ead4ab28ae2c2aa5185a0746c9cfe9fd90bdd68f2ba05291045a296d566[0]  <= 1'b0;
            I2f3612471464f3108bd427b6427c8fe79dce2b8e23dc4bb74cecb7e89a3b64a1                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ibb36dcaba8439f48b18ad2dc8399df26b940f7cd815996635da092d41ee5b106[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I32ed4ecd4363760151c1accda085c9afa3efe63daf7a312feefc00b804401c27[0]  <= 1'b0;
            Iccedefdcae7039447a6901e1cac8bf962a9f520d3b343c2b00e654c7e11a24f2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I387a4fa48a52a029d2bb0c8e5163f15c4cd55d570db8d89e5f73d7bd6e21ae5b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I6aa6d6c6213348ea0cc3e8b207bca2c1db81499441e4ed721ca0ee01ae831291[0]  <= 1'b0;
            I8252bcef404ae08a2a748c98d672c368fbe4187f26e788e54d93af9077f92a20                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie2ad7096c10eafa6e451ff7793b2dda562b6623b1eaeed56bbad4019662851ac[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib4f23d2e5f8c73110ae24212c4ec0e7ef29c09c8178ec3850f061a5b0386feca[0]  <= 1'b0;
            Iaa2493521eb50d228c5b0619dca5c86b89a165f9855552ce98021778cc196f8d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9de97cb2569312c40a541c0038e02c03024581050590e5677dcde888f4c6c3ac[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If2be986b27ce8aa2117f87e9a144015a10acf0a07847f83acec2804b9e987e8b[0]  <= 1'b0;
            I69d7f0497be77c5b1457ccdc35789d454bbe83f7d9eb458527d737a2222c7796                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7a55e4af3d00a3684ba08ac52c3dc7dd0188efbb684b859ecf017f783fce247a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I9f17331c6a9858b60705d889b5b77078042cffe9e956de20eb067ad7e70626b7[0]  <= 1'b0;
            I2c40224a96616b7749f39d78a0c07514232a019bf2c9ecd7340560f5aa5ce6bd                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib1644713e1c2c63d093c8af3a2be146dabd70cfe25a1a6ac062174576477b113[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I2b70416e96231188e62b7bcf0300c4a5b2d2139449150d31414b92ae075aa0e7[0]  <= 1'b0;
            Id95e503df18410329be5e7761b6857182c75f7d2b0268d0fc377a415c89cad3f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie907506d9949011db3e41c72b9581fb832dfb29f82249768fd9893a3de358b35[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I29599a1dac362c87f4780a94478787a718f63401d2051ccbfe543b44e49b35bb[0]  <= 1'b0;
            I5cca65d1f11141b49a1136898dac8226cb1ec1654c8b8846471f1e4c36bcf3fc                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I678204e14a0213dfa7135814f07e5f6c4d12452a503ed555ca2c20c10f047d5d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I5ff7defb023005e77164f9f3b852fa60ce897922c6b814015d3436fe1d1b4a44[0]  <= 1'b0;
            I6abf4748a0be2d4365fd1d9b53a44c3183015e1bdfb9a3f671eb5beed231eda1                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ice68b876a3b3943637914d8d12aec7fd37cb867f7a7c20be11a66dd85803827d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie132a24e667376de85b8fff9a639698df164043422122a8058c968bb7996d3a7[0]  <= 1'b0;
            I56bb103437d88864c0ecd5bea1ab5a0313fef2b904c52adb559e19bef8f716bb                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I35e112474e97e65f8e8aa9a4dcce274c7ffda9cdef901ba31801b4daa68888fe[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie8d5dfc9a77dc01055a551c5f37416d0b13ef83428bf751fb9f95c7d10442697[0]  <= 1'b0;
            I5596d8fa3572e105a1618deba542906f0ba5acef8d7b0a48d0fe2e4eb3cf7481                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I84992c3714fef30f928dc3330821045f20e176826278d42a9606f2dfadfcb9c8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic94f2b10208cb23bb5f5b1a46c11c3bbae038308b385373cfaad9a18e09ccb90[0]  <= 1'b0;
            Ic00f466513895a54a6974af570c7bd5aba8c0ecab5612798bf512ca88f27081d                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I011fbcda61a4f528c38920d0077565c4592c5f6d1a2f5a1a7dcb6a4a734e0c83[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3b79a6c69be124aeea9d1444f9f985201b55ad0d7a4767a01f612eee12a6ad73[0]  <= 1'b0;
            I456f1fae558de9875bb1f76cfbb1840945f61ea1bce9c9bbcd0ead15d4b2803e                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6d2154a30adb0faf296cf58ca9229eb1a298767fccc4a1214092a2b977f7442f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id3ac4bf805d3981ac1eb1b396b3da5c0dbc68754d89668f0a4cf7c6f2a44ddfa[0]  <= 1'b0;
            I7b2c627cf9d530af8ad8ebc0d3dbc53988ea1819d98b5e36e1517e21cc954782                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie500f9b1405b49a263908c145ee4a337f2ba4cd2d4d784a2acb77068d09d1662[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id77fd99c6146776bfc20804c67ae41b88cb0441eecba4f40b87828956b7158b6[0]  <= 1'b0;
            Ic61cceb25c811577024c75e771c53089a2adb9f80e6a622eb82f9d8e5bbb6c16                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I26997f7f737ba99dcbde55d67661cf9e4efecf397b1ab3ec59e0cc5d8654a75c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I650a7220fd4eb743f652c6c1f9431191621f9fb1a5b5d64bb9649b43bad5b8bf[0]  <= 1'b0;
            Id8edf0b11a998a6c5737c8877c9b203e44c777ca9ee01cce63f046a6bd375c13                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            If6181a32c0ba3cb93e47ed1f1279bd4e739882c2905d6d64d0149f26d052f0d0[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib7417e90e9dc35367f110c364878657dbbf66b1a714d5807e6347095b833c62d[0]  <= 1'b0;
            I2813295228131e78d6af31808dc1d9a6f712ddc60b2629d5329dc6ee2d07c9d9                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Idb4bd19284288df2a5b701cedcd57347e4f7c37947ec1588daedf3c9ede0a12e[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ie59a4afbd0d65de2149e8c60229bce12b77f8f1b2b232a11fb9714371eced2b9[0]  <= 1'b0;
            I6736fca4e33cbc58b4658d91a401b558b1fbf9b3496e1830a8d7b4237d0ef125                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I4be880e4f25fc41932b9ab9295794ffa2f334ee5338ef0d59894d18918d3e0be[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Iad3f7ae48f752d3ee71320875a2d1d170e879dd5ff51cdfd662241e6a30fca6d[0]  <= 1'b0;
            Id66c49fe8c0d931dab1b901945cc3926c6e7e3d220480a28e0099a0656241a03                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2dacf26260c042fa148fa6c4e97bf878ad2e89e221acc0616141e1841b0c320f[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I4e9c85ad6975994daf65df213a2d2fa5a6a2abd91e66d9c9a6f540caf4c2afe2[0]  <= 1'b0;
            I1d8a87a805073dbe04ce0f76953a234bceb3e6027b2a187071b492f644843715                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6cc3662b07a43d62f870bc24d55a9e5675a0e50d923f3b293d7004c2c62ad31b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic8f9966a2711f4810086d09b86e16ccf0d31339d146ad5c38d34c973c757947d[0]  <= 1'b0;
            Ieb9ae0dc5ee16583e8d05536052b61089e8004344fa0e3fdbc88c5af5119f293                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I670beb5586ec69af20e65eeaa49be81826908f01db21d27643e2561621962b87[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic1385b7aee4e3b643e13733b56157e3e92e638da28cd1234e275fc9263709f04[0]  <= 1'b0;
            Iff41f572ab79a4cc8e83538b32d4861e88ebdd0a9ce51555053943225158c5af                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I88ba583883fb596ad6cc6716008143d6b643816e8e694ea5f32ba95f3cfffe48[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3a173e6b224a6415ad442ae28a0af62756975427859bbcfc0af6c8e5effd62a6[0]  <= 1'b0;
            I7f8fe2415810e04fccd129edfe956981aea020e4b24dd85d59991f4ef0131380                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia8545410ad46518007f6812cf6132f4f4482933818a0fe103dae14b1530518d7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia5580120af4590da8aed890f81ca17929e4c998617df957686c095e891649c83[0]  <= 1'b0;
            I5eafefae338dc0fdd7610a7cc3093d323fbd397263d3c8b7546bf540e77d60de                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7018895fda9af57bf39b18e9edc144f8854067ef25800ef8eabe76015fc207b5[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I58a3910d475757bccbde2da0e6b5dd5723cbe44e1f4d3e71ac2973fd2a03b3a8[0]  <= 1'b0;
            Ie5d6a774e706204102b6a2d413e41c538f5e61284a19c7a47c42e356ea77d072                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ib57f995d569a522f5562976385f777cd6cc39ed15491d0ad8f88cc0e908c326a[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I1b76b0f61e714e21a844e429806d641f6a24f0eb19c23a3c2fcfb76baaf3e72a[0]  <= 1'b0;
            Iab62db2e5fab6a7735067ea4afe23d7904f71c5b92219a1ea7848fa358da3cdd                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I35636bd5c56cd95d41880b5c936108a3ab7c1517a8e09f76731b2154d39c87f8[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            If0211848e6cda136970069df5b6156d4ac213717491c68ed49ab39d2cffe9999[0]  <= 1'b0;
            Icdf027acf32cc766a4ab1f19373a58cad87f74c1ca1791f66e958de6f18803ab                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I84280195e0f72492aadcce8eda907d5de2e05dc16b9c5ba1fc2f345192ade355[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id23ae21f713f4f452abcb1c1839b5524c452bb8bb0b6c35683f9bde212bc5f96[0]  <= 1'b0;
            Ib087093eca2530f923f55a4b4cddc83869730b169ab16bf26f6378b580da58f2                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6532aae67414dd9e03b874fd4b6a321437892a7d89bab17ec2d5a684aa9ad55d[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Id5bdb0f5a920710b1af7cc3abade245196df9d1ab4b7f26277fd93e1bbee5556[0]  <= 1'b0;
            Ice19f7340dbb41a6b126bdae27e69b813b5d6f73ba4db6ee79715328be678511                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I7032c41ce2651dbb03999e2120193d71ed608e40ac2d51329837f3abc0a976b9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ic72616171e7fb8489fa12cc29be1f74602ff8e4bd28ea085e938da615238a0fa[0]  <= 1'b0;
            I575538bdc858fc8c843bc6b68625f1ba5fd33a904937071914caccc65f324a49                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I9a800fae8c9498d12065155e7e781ba817ee2b03ea6540813400bbe438f4691c[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia09db6bd7cba6c6e15cac4c6ad0d4c98235a7437beeabca1388fb1b4dece5d67[0]  <= 1'b0;
            Idea12ce0edfa5df65e47f6496f2a457a03907e9d62de2cb3797ec2cc6c5adf07                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I1dca7dc76f83994b077209eb2742069045e743b6eb763805cbddf87e6a8fcc34[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I15ab76f6e4824af9b3b4f5062e8dd3c426e1ff0c5f68e4733828c710eb7bca54[0]  <= 1'b0;
            Ib368839377e69cd28a997a22724c32efdc8820a04f9b5f93d9877bf398ec6e61                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic16409f8fa42d6ac05643c3943352c03f19cfee0c3068e96d6ca3630b8f2cacf[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I12b276cd6b0aa86ca2e28dbb1f4008ab140668e16e4ef96604a6d1741c7f2f95[0]  <= 1'b0;
            I67be614a904dd4d47457ba0dc7a19b2e9f8e4231797917ef3610aea55d5ba3a8                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ic66f776d5d728142606f048e3cf27e927f094082fe1dd31f90e757beebd5b5e9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I01577c8c0e65ca47449450a8b2455ee84cf5c48bb26a0799b5523258a039ae40[0]  <= 1'b0;
            I7cd598a52037f986959ad3f02b4b2783a613170f53a7e49573c5da74f1cbf614                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Icfe7c47d401f26676f3f8f13e34894792fff7a3881d754de5b4ac1130cfad989[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I63ba87cd2daa7c3c625d3ff5bdaca7f2115fc2d65e13972a22b2c2ae5b746d4a[0]  <= 1'b0;
            Ide70b17967ff52e323b4a51db51e71445ad3c5483c745b2cec2cc338e5f42f6f                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ia6852c630d3d698cbe47da7b990ed04d4e0b995b3d765ff6a8146da11e42dea9[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I576afeb6020cc0a8e35837b4b96968ed04cd444999558626adac849848fe7c6c[0]  <= 1'b0;
            Ib28a3a83a3be0baf561a184b6de18de0c4847ff892c403bb9da441f017dd5efb                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I5e5d78a5f1d49833052eb3e84c516dea9f05d6d49879c593f5e0b9745f84fde7[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I3b8769ce28405c0bb978c458bd6272f10cea5338af4170ce4e93a8932ae8dcaf[0]  <= 1'b0;
            I2416ae27b898336a36264980b371003c06275245f514135d0adac28d88379cf7                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I6454add174b2968c545e831c5bacd6b95b351b7d68448b3fa9c2e5476a8cca35[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ib4638612fcabc0a2c2f2bba5a2b9eb71cdea23575641b3f81fb6220fcaf284f4[0]  <= 1'b0;
            I2d58b3296656a43e75a58883e59a576c0bf73dcd6bc28a939582be7ce0a0ffbd                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            Ie062df11427db764a0e09705579e134d08f4ed2a027e913a43495db5d5fb9051[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            I16ea389c88e4591f7686eae3f1988dd5361bf893895697c0ade8627986a9fc5e[0]  <= 1'b0;
            I3f548241255df4c4a5a8b71a4352ffad6c3e5278c73de2b1afd1a1f1f1f94684                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I2a2245385398379002074dfa174bde148f97bb3bd83073505b550c0c0bbd1e65[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ia17edf214ab782c25bbab97f6bb4e04b2fc46d41f9a97fcf617418d54ab76a7e[0]  <= 1'b0;
            Ic3ef9d69272fb936b5ada08c6eb60ccaa6acf7b139689e5cb44e0ab76c0ee24c                   <= {MAX_SUM_WDTH_LONG    {1'b0}};
            I862f2564a9e7f99bc8370fe12c1a5e57612d564f1606a21f6a468d558c23fc5b[0]        <= {(MAX_SUM_WDTH_LONG  ){1'b0}};
            Ibcfba9f1fb81d976955a1fa7101f0b0db16c344c82cc5ce81f50dd3aa2928d37[0]  <= 1'b0;
       end else begin
           if (start_dec || Ie6f0821795a2d09a9d5d9fee0deb445f74581e2f81076cf0395d62fcc7ecd5c9) begin
               I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75  <=
                      (I96fb06aca6108479f7e21e1835a091a9060c2925cc6320c8ed71a0a0092bdeab) +
                      (Ie000dee1e3953811fe9424588b71a7dbc88f41ec69afd16e17e8fabf141c31ec) +
                      (Ie873b138e19cd7f7e8afa8bd8f8c4610b65d0fcd647e76d880d25f6fe36c54ef) +
                      (I8ab1772a3bc752331b0bf62069643cadb48bc13bbb06ad3eddc68ac603d73654) +
                      (I4bce49360270b653e45b914c493ca8e5b74beb0b6b85838bb3b54f1f39389fe3) +
                      (Ibb4ff9ffdb2771ff640bf958798f8447a0dbcf15ed0ef9f82068826ec621de77) +
                      (Ia4691d32d9e84827a250e0b3d6ea8142c24c9df4ade01c19583e6cfca06cd990) +
                      (I3a1380b85cc7f797ff92d02b7081d1ec3ba069aac74162ca059c399daa10690d) +
                      (I14919dedf2b4d4caae8efa1726435d1946f48e1e9b1052133bebe8affeb3556d) +
                      (I852a201bdaecd968b6f9c9b6bd64dc8035a17fb92ffc806a690781666354b069) +
                      (I345c0aef41ee2863a96a076a78d92c7498f50ef90e82e75565df1d1f38a08161) +
                      (Ifb94a220081758ce91634fef64be084898a662f7c0e8cc9f86859bf3852b3efe) +
                      (I5f1b294a0702ab37f94304ae67fe91abc04c397dd682d371126a7ceacf7c43ec) +
                      (I81aa911c9f6f4bd88314aa3c5310efef6c40219ca93521bbea3c1afcea7bb48f) +
                      (I97f674eaee005fc7a54ccb648f5a0a67cec041e895d62eacbcc9a37068b912a7) +
                      (I7628fd0a5ee3ec547c1b4798a4d76de651807424cd18f0b3b8a3bea849e6fe0d) +
                      (I1d8a992801d3f6a457848578ce286b496d4e2a69937344bdcbab4e8b1af1fe4e) +
                      (Ia28f68b737aaaaa6b98aa5e9696b937e564754edef217740c414c16fe2e485b6) +
                      (I099e314496f03784e5504a35292defa79dc063aa81e6aa8764802f7fe3a47114) +
                      (Id4bcb557769f043a7275ab01d6d9794d4cbbd9309be38f58acc307a1e693f347) +
                      (Id1bb830ea0f92a1c0ed0addc915fc85198e4744c4bf7369b4ee1f7131f5f8542) +
                      (I31009872a3e84f78bbf1f12a7da708c45e3b708bd943b6f4561ad436164b12d8) +
                      (({q0_1[0],q0_0[0]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[0],q0_0[0]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6  <=
                      (Idd9957e5b52c4d33e24910559d8203415afdf467bbe1c9de950145282c7eacf0) +
                      (I6a09910e62aa0cf665f69be80c9ad61f2d31115012314b8188cf79fae365626c) +
                      (I3d6f6b104bd2ffb35ea6782748bb777ec7eceae47ef2e1d18d37d1677d56cb80) +
                      (Id5055b759fe480d476c4bf08c420a5dafe9e65cb03c6d6991c1d225af0a51d7b) +
                      (I93e543ef3d58bc8bd48a279299dadae1d7f4528c3d09d7106b969e15565d3a15) +
                      (Ib6ff050679c6366efde7b9809fcf42051f107c18863bcea79d41b5fee0603e9c) +
                      (Iba81256fd46cc69f1367fc6ed7b712d2695e099c52b476f9b39f0a13404dceaa) +
                      (I608b794037b45c46a29ea01e378b63a1f267c4b489b0866fe2f6090936fa9d44) +
                      (Ic48347f5264e8e479996a8dba0171a108b602be1e1d24b2fcb43cd2bdb82f61d) +
                      (Ib62b5b3c80d193b97bd6b5c0d5678e424026381949c3f24546d367df930cbcae) +
                      (Ia7900b5a01cfc1c4db79ca653f072956c13e2040cbd94cf07de2f1d969222fa8) +
                      (I1aa136009f34c39a8dbc39b4444642cd09c9cd2f01bd6310287d4ddc9bedad85) +
                      (Ic195e053a186bcb0e653c0ddec75c57d1b3210c583162dd90978858c98fa53f2) +
                      (Ic859d34db6baa83e73a8627c251c877e93f15653973d0634c42a8ffc9f628bae) +
                      (Ibeb23788ce301c724494a2852312b38344c27416a5604c0145fa330ccd1f290d) +
                      (I5ccf8e87b0b8e8ce9bdf4b3329e4458a628f2568184f82b998ac62ea28bc0307) +
                      (Iaea7277e745e05f803325e0f19dbc5a54234878a9a3cb2cedcc013e3942e9cc0) +
                      (Ic94e7c887d7f24b573b470820c36fe8a0fef750e2c46675f8867d78f2100f1f9) +
                      (Ifa0b8243f5ab6adb88a70fc1245e3480ea3fb3f3af846fdefd0613ca91d7b122) +
                      (Ia00cd24df6e6b22b466e1492500f1948b3ba3d70bdca407d1c22b4dfaf374eb7) +
                      (I8b41f817a4008df0994e2efa6b33eb847e82b031082f90a767467ffc03cfdb93) +
                      (I8d91c857f2c8154bb09d456ff73ebdf81e3b7d9bd1c57c2e6b8c2de74e55cf48) +
                      (({q0_1[1],q0_0[1]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[1],q0_0[1]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee  <=
                      (Id0f930aa222bd91b8a7d5f80a38d84993a63fa1c6aca3d37ed259294e08869d8) +
                      (I58598429d44ad951f91139a213d3b0bdacac6d71f1b9753886dfe1d39d0024ac) +
                      (I3cca3cf08c967f80e7e255a590bb9c442abc535cd529f7ff304f25d5519dab04) +
                      (I42d1b7202048c81ca3a8bba0dbbce65501cb7a519fde37085c68d01db7edd635) +
                      (I07bdf8f629cfc9c094023be167a717880dc3a42099b01bffb431036521cd6019) +
                      (Ifaa925832248fd0e2f5841096d9618c2fdaa3c63a3130b57f493782f96473088) +
                      (I2c22aed0ed8abb0cb8906a35a4d44cfd7cc68b2924e474680a2eb6cf7caf5582) +
                      (I31ca3705bdc7e063c61023d93193b3ced40cf440afd817d0d730f6c8d37f8b92) +
                      (I789461a909fa4abaf3840dfca4f63bfa63fdab389e149fddb7d8ae2b876dc912) +
                      (I6ff3298d93471156b56cfbbea17c8dc0405bfe8654e9f830bb33bc6c9a649b3e) +
                      (I9eb30c75f8d71ade925633d7c8bc6b948ae519cdff33ddb885761bf72a8b0869) +
                      (I5456c559bdce4d65af540e4c71c19e44227c62e5c129b7de968ac7f311dd76f4) +
                      (I98e4b84e98742d38b206ac059ad123966ee63903c616b9c31b4ba9615edb9f40) +
                      (I40d7eae63827c6efe2ac480c8eb9f8a8f77bbfa845caae02d137397c9da822a9) +
                      (I30a9d5330fac5c3ec7b63cfab0edcef0eda61dddb23d2aabf733b9982c12b4ad) +
                      (Icbdf29918b91006ffdc8b68c707840ee6bb9c27779dabd372e2033888743409f) +
                      (I7f6b89a61d6313029102fc48e92a54ffdece30e9eac1191d840c488be69d8223) +
                      (I9471414594b824d60836981bf4b9931c135520ad1ae7dea177e0bc591c2572c2) +
                      (I0e9135a0817e96971dc8c4fe6eec717a563c44738f7e38d5bfb2f4dda8c77876) +
                      (I0847713503570d7ab3efee12577ba27aa81869a22b14ec8a244fbd4665d566f4) +
                      (I7b529f16d1499766369f75cde5a356cb12c06d21f42a10932edc6d54146735a0) +
                      (I1b93b1b2c5f55e2267a4deb4f75ca91039d6893af8e082ea85b7a5e9354117e6) +
                      (({q0_1[2],q0_0[2]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[2],q0_0[2]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493  <=
                      (I7200758287b0c7ed92552ced989756e1d49b5418181b9e36421da7e2694ed3a2) +
                      (I96e7a523360a0cc0f3abfea09a566658e5e9f3316c3c412f99fd6340d1b64235) +
                      (Ic4839247bb24d460ee6d963d31fc390e8d9d679cd73f058d94ec34a18ceb39c0) +
                      (I23ef4f4232fa0d8813a25ddca38a2745fb660c05dbe9ddc2cc33c47d45b3fecf) +
                      (Id5e78e4ed6db0562ed51d1da1f34242f54def8255088c3a1ccf0221ee8fa153f) +
                      (I17cdc222663e370d6ef2539ad03c45a7949d9606583c17568a24c528a3e8c12f) +
                      (I65e452247faa2c9d6b01dcbbebd5e8c31884c88e70dc8ec76d55aac7e77e2d46) +
                      (Ib0641eb8fe554f69ebb57e8e900f995c07bddadffd25c01781ba234b87af4a94) +
                      (Iee9c2c6a9b8e84402eb1e0de611c1cb8ae1e802226f2c07833bafaba74f1ac15) +
                      (I443435c78145236b927711299e8bedd0d29a743e3784ac22f70b2284b6be11c1) +
                      (I4a86387a3136768ab52d320fae7fe63c7c74bb5541d18889faa263c71b2bfce6) +
                      (Ia0c4bcb29e2939b889fb7a5a7b62b49a3eeb3ee6f4555518c9059cb34dfebc7a) +
                      (I3de9fbe37d08009f5fa66bf7c59debe7da836dc078e212968afdc608b100e3bd) +
                      (I7c6d90cd79e1b85ce9a5452570cfeec8faf9ce3e6bc886f66495ec2a66fc8c7e) +
                      (I57d80f41498f8d7b91410dc02e646a45a3f05d45e9b5871ae95d6432ecd2af56) +
                      (Ief90cf0b0997823c3071eb46b636e384077579beae3d85d29e639a7719763396) +
                      (I295d7aef060ca978805bdf65138e5bf134551eda9c396a22165a77a3091dfd28) +
                      (I73a855a590363c762c34008e77f73f961950c0dd71b795acab3adf40c4540453) +
                      (Ie38c638da580ca7d25fc0754497163d0369f31a6cdb4bd26663a759b74efd588) +
                      (I2c635a0b11af3be4774428af79ff5cbe6a32ede6ad03ac197ecbb3ca2ba78f8f) +
                      (I34a89a8aa68b1657dc7137437574877b170659ebdbcc93a772989e2b8b5be31f) +
                      (I9f9d895211b42c2c9d491349dbe7aafbad775942920197105c34837dba6563a0) +
                      (({q0_1[3],q0_0[3]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[3],q0_0[3]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac  <=
                      (I11c6d693bd6c019722571e1aa6eea0507f351a89cfc6d16f8fc51997981aea81) +
                      (Ib53bac100fd49f57a5185ff4ad973dfe8eaef6de1937bb32d9246dae9459442b) +
                      (I7ce5fe43a760b5a43815388233952e1bfe5d8b5a7c002f26ae2d462129aad434) +
                      (I3a2c9aabb8b064f82bd6f6571bdebdd704abb7526f4977a7b98613f883fdc62a) +
                      (I52f4d169be660862052b60924958cc9a0eb99b1454608fc48d47192452f8b390) +
                      (Iade009d6c5b9e00f5459c53b0c254dda356081e6965366db7b7ac42a992e3ae7) +
                      (I52dd625c97050874c15b1980a389843c4a7a890d73f6efb003c4324c029772aa) +
                      (I11bf8ca77f64484279bd3f36febe1c6869fb79b4585a800449a0e5c683c6aa18) +
                      (I255a6c7b69c31d60711a86b1f0da51040ab60c48952002406e028a200a835049) +
                      (I24bc395a7644f2a2d7702656737c32662f8c2e8a7e2b2d4c1bca200dcdf49219) +
                      (Ia84166c5479fb08b9d5bafbf3446230d231e77cb1a3034b53477e2f0632ca74a) +
                      (I544bba815490c8592dda0fd85cb612828256c09ba1431bc2632b74cc9cd2aa29) +
                      (I7b8225b7ff4972426858a8550dc67a231d85fe94426bf0812906f1aee0e2d097) +
                      (I3358739f5e55263208e661a339d6b29f188f07ef07e2ee7a63a24011a4f8568f) +
                      (I5eff39d324b6a8910fad41786d651086c622d331987e649ba4b3baae11ca40ce) +
                      (I4a5c4f290852b8c1baa90ae00400045825f13c24b546dc4a7848f91824185f7c) +
                      (I9af65d3592633577409561b2069e30c73196d1a4798cb92f4d2f14db8771895c) +
                      (Ie2261f6d4e2c2ce04997cd365593486e02a7d85106b9c3b568ccdfcda7a9c352) +
                      (Icf0b2747a9e17f2d2672f7a17111c6bf54bed7d8fedcb5260f25fdc4280ae727) +
                      (Ifb6bf654293ed3bacd2a4ffc883b8ca5e4dedea39e338bd1a30b21e8f8df2f62) +
                      (I0f4ede6017039c42f04051822cfc539cbcacd77427efe92d393ade1c10a46462) +
                      (I23e0423ae4012d108a4e6a495814e0e6f920fa6dcab900bb35cba7b95f590c9b) +
                      (I571233769cc63838bcc3d61e7a5e95805c3f4116c0053dfe86831eafff7c32fe) +
                      (({q0_1[4],q0_0[4]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[4],q0_0[4]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d  <=
                      (I7fbf7b7f7a1f0155cb188ee4219620cb35a2fcf98d2687cddfa2508273b70154) +
                      (I4f56f225d6fa40e0469f803c2f72ca27e9c45768ad2af9af9ad10e529e249aa0) +
                      (I634dc6f7c843c6e4c63ce6a21b9cd7a386600d1155c0696988403fc1ab790217) +
                      (Ieedfb1902d1f76f95f5f971b578c2440fa5de47dd78e9dc70c35698f813048cb) +
                      (I88272c473a90efa576a83d0c277090f5814599e5aa192b878cde74215909c46b) +
                      (Ia3e877a9f66cb7582b125e56b7c3f79601eb8e700f54e14f967a4d9df9b5725d) +
                      (Ie278ca9a470ffe4ac78bc335aec472b66707cf02bd91256aff2e7c73b5d2c6b6) +
                      (I5ef535b2e573d96fd518cbd837132928a2a0c6a25d4eb3c360f1cc0aed89656c) +
                      (Ic486b9953b158eae95a2d8914f8144e669e056675946d245c8239bfc249a16ac) +
                      (Id89c8a47964d1e4aa4bb9e96a79092cf7fb55eee5808d6323ecbdecf8926adcd) +
                      (Id1e80f29821e7ae727d759f44b21e84843025c938468caf7c8adfba52f1cae43) +
                      (I7530c712ec14c8fe97d1699177ef642847c5c1ce6185d1eab39b8416b562b454) +
                      (I41b365f8c613bf86dc5e2ed41719ec6823046127babf87a083503ebcfd38ae75) +
                      (If9bd4d7f3740f15bdf597de00eecf1cbf2e3b4efdbacbbad889c0946a6b34a24) +
                      (I31c470f2adda0a23b85c3245646a168f2478bfdff11a434c1455be20db703c64) +
                      (I9fa9c98579041b6735eb78f7b3727824dd61991c6a6d91a158c6ac65cb20b05d) +
                      (I9fc6fbd6f2f888b9750fa59a966971aa6ba6fe4eee8c8f3ed4c3ea60141a7d23) +
                      (I8c133563a8b5e359a6a45a7f3b4e939fc84766f9fa09634d18e5d2101d0c0645) +
                      (I84238bd7e53e0dd7ba07efd813661c8cd1648b76c44665dfe51fd07dfaa9b249) +
                      (I6c3a9695a1c1d22809b1378e82cbdbebc1ca78428194df50cce0a69d6a159398) +
                      (I4d032ff7482be75de7d2b816ddb2bebfa9e896e45fdade2b5f81b35c003a59ac) +
                      (I6b4d2a32c92c22b1cfe81ee6620c69af1850621deea406d75f098da0542843e8) +
                      (Ia0964979ac559942d1da1c41ecb3d9e94c6c7c0da3d16177cf2379db8f37aa65) +
                      (({q0_1[5],q0_0[5]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[5],q0_0[5]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e  <=
                      (I236cce67d0aea9f9c8d5ea3c39cb598d55f734b44ad6e3972e7f6b91d56001fe) +
                      (Iceb8741c9680982b02ba9fa2dd76d3b45155ca5f688b70c41d66f3b3690dce42) +
                      (Iac9f4a2fa823ae63e73b655020376580991cd4b2b3123204a757afeefe35a10f) +
                      (Ifb57457918458a6aa9c5df68dbb83243fbc49b3b7037575f43749dfe1bef373a) +
                      (I91589fd8a2ab91f079bb41631c44926b2c6f83b82448d758d97578c314d0b76c) +
                      (Ic20b5a20229313d70c01a5f53e13e96095c1d8695144668e66efdc81efdd8374) +
                      (I53e90d4a2bbfaffcf92f2e9fd80c491e61990aa575337df13d24211a558315a0) +
                      (Ie57b3acbbf1d1593e02ad38bc0e07bb84db2655f9282adb3ac5edc311e882641) +
                      (I632095e999af63661b01bfe8bad0078cfc2e74217253d3971230968c235bc526) +
                      (I6a66a98136fb7fe52fd830d869dc53a3855a545aedc1d16927f76bc12e319060) +
                      (Ifea15bb5031583fe42f92f554866179105e46b1eac3c6b691958a998c26ac2da) +
                      (I8b2c2b27add863ad56639a306f803b656ee8f91170e649d29aedc5321181f857) +
                      (Ie3290070e785df28e64ff4df124d14c370c9edb924d5f35b059a6c82e8373f91) +
                      (I02ed3128371185efeae1e27046aa378006ec78d7c458dcba137f69c29c4363bc) +
                      (I8dcb7a5498da4a9d3e4a76923e84c88a30ec174503cd435864a066ff0ff464ba) +
                      (I94024b61447a332a2c36a75bbf305f3fd80606bfbfcc4ee8c5783e3910e9840b) +
                      (Ibcddbd4e851466c5ff49f13244c2478ab6c089e6d8ad294cdfbdc8451ac6a895) +
                      (I50ff347e89fb452beb071f112e4a51e074cb3d66bd903552db23c17670286e7b) +
                      (I8b5ee5d271abdbdc518ce02f900da21e858d3e2530585fd859690a1a71502434) +
                      (I54e64fd01d9aff7ddfc4babeff6703891da38578bb141d250c4ef5949d818cfb) +
                      (I448065f71638c5abddd1eba1fcf567566281d5b4b23ec4ff2d2208d32a506fbf) +
                      (I6ed6ee11f6983e96e7ccc4e4be6ed8c4ed166ca9075b9cd218f26f018ad2140f) +
                      (I0678dba3dc1a3400ab26e223257bf71c03f0e8d284810653b5e507fe964427f4) +
                      (({q0_1[6],q0_0[6]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[6],q0_0[6]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c  <=
                      (If34d8ceb2732716c923a7f250495970948ae431d5f1e0a025618c1070940ec39) +
                      (I60014273d45dd5019a1b82bdc0a65e44d9a16368d996c8c9ff312fe27e236171) +
                      (If16869134ec7e59b567e29a1125f0d27eff7a3c612240e25462e2ee84a7e0104) +
                      (I8d95c0be0c84d3ee590f8e77065a6ef224e0a75b50aeadea980f9ef4b8d25001) +
                      (I28940d6e8fc5937055f8f50c0d65ac9fd892bdc9f0f2a571808f930c8ad21717) +
                      (Ifbf3cda7e0639ad343a64c5b3d2f45017f1d280bf72c96520cbf272104c90ad9) +
                      (I4aabce2cc01e829bb9c3d6a984cf2b5bf9230cf3913db788c47a932ddf71b869) +
                      (Ic9dc8459f6cd65f223a6386c82f754469ef74fbab59ded4fd1370fb69136c847) +
                      (Ib22de4dadb6e63ea49c52cd8bc86dadfd7b73a002dd8e726a9cf1b7b299a8c46) +
                      (Id6c8c2ebab66fb903f108466c8d15060ed1328fe9a979858569c39069bf050c7) +
                      (I385f4177f3a22b6fa4a6352d164c7d54c94b980806080c51d00a65f030966110) +
                      (Ibcf016cc83d0fcc2c731aa53147c199b32b3dc7a9f1a255e1a0e31615077205f) +
                      (I7e7be31550be1cacb2acdb27d5120769dd7a0a49efb833051ceb83c8cf691e21) +
                      (I26d08096b43367ba37b8f6dcd919bf4ecb9c660a39f2c0ae29f655e42b88887a) +
                      (I2c200a5ade27683d4afd55e06371f9880a7bb99259e2ccda5c368fe46bb385bd) +
                      (I92d28f6c97dab90de260df37f619e0a9000db48e278327a5c5d1528a34bb6dd2) +
                      (Ib053c04dd4e330e6784846706317bb6c8b12f9b36a57ee12807bff7de8ba7f0c) +
                      (I0f71479f871309f1717e7a1a2372ebfff4623c315cc31914588df3896740a074) +
                      (If49d6a59c1d539e369406ee4e8a2ebb30199f46c335584e62921f98fd811001d) +
                      (I051f072f564eefd657cb4d59c1c851b56df2e70861d875f3b4c9b95e8945db08) +
                      (Ifc8302f040679d23faab1ed8387a8a3aec85aba86ba9a78d3ca903126266af4e) +
                      (I2747ce9b7349ed89e3265df62bb0d0e612706d8c1b61e30a2878094662da8ff1) +
                      (I3619e836fee4be75d6700a0e72e84df3a5a61003227363b8c4d348b8353075e0) +
                      (({q0_1[7],q0_0[7]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[7],q0_0[7]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7  <=
                      (Id658b37d70ac8e3a324133f475a77c7948231571aa66ea0dd11b6460fca011a3) +
                      (I737ae96fe290087c8ae686b90b2ac94df2185f7ad8b4252a6ec850278ba5ea9d) +
                      (I18777be7a1745485d18289e0b4a6e43e8a2e6758be0967b8cea04a3b0faf973f) +
                      (I1c30d2957a73fc51bb7044b869e28e0a8f6e0378a6098ee5e244efb43ab6a690) +
                      (I69f7964c2f630ef03f49c2a6cac12420e0998397470245e6afaed2546b33775c) +
                      (I6f63c71eab6c2d7e3eb41fd78c9e18d6362d2dd4100c72b43d3e4b9d06663165) +
                      (I23c91b29deaa2df1f4d96e343f6fb852a2b594937a4f62dc4be1fcbe0347c439) +
                      (I8411087f9f6fa41d454a74dc89e5152e5e8edfa501c8753bd0735cec3789f14b) +
                      (I119a98150511650722429eab31b5785e99128641bad59a3cb31e42158a648c48) +
                      (I28a2b1ada19dc69ebe4949a75633b2f543159d2d1cc169f3bb6070c1419878e0) +
                      (({q0_1[8],q0_0[8]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[8],q0_0[8]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975  <=
                      (Ibbbf3f4aa7f74c37a0e8ac8a675ac9a9fec748ac720e6a78e9cf937dd089b8e3) +
                      (I59a4b1b33d114a1b5bdd708e1f856f4bf729c6b86a4064967ca1faf779189164) +
                      (I9b13cfb3566db96edc7c018b88f158faa57e4db029e3982290989c6fc08163b2) +
                      (I8a1ba53134dcd1141a6f03dbed0f18ff7be9728dd9a6d6b138ff266c5307ba24) +
                      (Ifd2ca31ff3eec501f34892055a36979681d27574ed8007e4df5cc0109b71bd89) +
                      (I6b2620e847ea73b8618ac7bdcd8236c4278de3bef0bf1511ee9779306438fa38) +
                      (Id2cf59876d070e0f34ee834d2691f7fbdb039bc9273329e2ce8eddfe736f0a45) +
                      (Iae213c2ac7729f8efe23deca256bf56f030403ef6ac00a3bc181414b6a3aa75e) +
                      (I08e50de7e2aae48cc03a9959d08cab30d3c1c2ba8c4ef0799645787b0c09473c) +
                      (Ibf22dd3f14f19c3fc769966f72e8ec980dc79c2991f69d03ca2defb7f720f880) +
                      (({q0_1[9],q0_0[9]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[9],q0_0[9]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948  <=
                      (Ibdd37577b403da9aa72ec3f4707379b1151c0b15edbfc4fd304c4e35c1672da6) +
                      (I8e23f89e84e219d5351bdfd4aab58f61c1cb310cc731164c6e0dd2eac37b07af) +
                      (I3baaba73f51f47e6a3f2310f692de9f7b9a871c65605e14d204d6965153ff4f0) +
                      (I82d316ed1475017844ea73f32085b755d17c9fdafd8191df2e363496e1950869) +
                      (Id9e3ea08b52843b4a9426b735967bd4ac3d49bd67ab8fc85688b0f55e6df186a) +
                      (I77e34c24ea46e99b6bfc0f960d428d6ba3ea4f9261d5a183d83c386f259ab431) +
                      (I930ad334ce972f0b5dbddf698f6101a196d8072e90d8144b31ce3f4b48a73e59) +
                      (I4c0096e7bbf30db97520f824e05dbc28e6d1db344202349993fc68cbc95d6585) +
                      (I75c796f56576dfba821e867b0de1a871ef35851371c3aa422532bd287f02ee11) +
                      (Ieee1d2436dbda6f58f19df70b691a4ff28d37db8ccc12e04413e45f80d7124e0) +
                      (({q0_1[10],q0_0[10]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[10],q0_0[10]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f  <=
                      (I65b0824920910c82c7d677c2dcf4216e86940b3edc0b3da85d8f65505f58ad48) +
                      (I169d92aaa7eb4f8516e38745955b91d8f6e0ff43cb212186293bb78884282978) +
                      (I492e47d35231729b266a9f31aba61a3ac2c93a9786a20f6a152d342cd1d0b911) +
                      (I2624a2d841eeb09774127e5d709364f803826266b46f0fc3122fcdcf0aa129e6) +
                      (Ia6414b3aff6031e10856953f6b15ffdb0971aeb680d784a7199386be15624ff6) +
                      (Iaf94ae58c1d9c9206d02651cd03cf2e02bba505f76b849158530a38382396ffa) +
                      (Ia0a40c2a77389cda4a8333aeaecf37a2595fbda87854a43162ad1299544bd9e6) +
                      (If692b993dc571ec401ce86f38a18ea4f96a797b00c04699ce83ce875b7c31730) +
                      (Id5a74d0be90678a7b69691c10e4ab75b47914e213e67eae2f20d4b58e8a8d9ac) +
                      (I47b54f01ac82a9eb80a681633a06c4e1d432d358091e9d079f74484f40ab3e09) +
                      (({q0_1[11],q0_0[11]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[11],q0_0[11]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85  <=
                      (I6201d3c2d85bffa03f368b5862fba1b2e0ce3735fcc8711cb8107adf16ccdeb9) +
                      (Ifcc25cd8dc442c6720ac0f764b432530aa63681953d8ba16b441892ff5966bfa) +
                      (I256cb35fd6d4e6c6e1c1a9b42dcbc307f858e5f9525acee9fa7af42c820664f2) +
                      (I67183da8c2763243a285b7cd41d838337f98eb6e59feaaa0a9150bcd6c29877b) +
                      (I730fa6d01ade8f1439b29b955c5cff62700a90e523a4f4208ca2f9978e59afcd) +
                      (({q0_1[12],q0_0[12]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[12],q0_0[12]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd  <=
                      (I37084afdf6695d3b8fb0530643c8b03deb2499f4f68ead04e3b5b79aa4467f73) +
                      (Iee510842ece3717ba6eefc3ccd844e97a9718788683d4c7ceaefa6ca0030585b) +
                      (I53d3de58d6308b770e4a8884447a5f0b92931c8d83c62c86714b6e539b498894) +
                      (I1e8142c7ece070c02ed90211fbeb423bc2a4ab19fae011793be99c68ff103705) +
                      (I425913b12fc3c865d95f1caead00d8c49de08765b634aa444243f4a03a53d0df) +
                      (({q0_1[13],q0_0[13]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[13],q0_0[13]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03  <=
                      (Ibe0fac26b5e106fc1753aeb842e8a04067fc91c95e358b1caa58db8192381837) +
                      (Ibadfd4f0852067e83ba6f0d57699585ae20eb542d1ad8f2cce3bda0d043ff2e0) +
                      (Ife27bd449bf6acad3f06d6e337bfc29c612ba6b3f06927e6f9699ab24d1e836e) +
                      (Ie130bec82505842b184f5dd86865ab095110bc65e59662767e152f427dd7462c) +
                      (I2abc1178fa35959d8eb41342a7d7289e29054439c7bc06adc61f3a1d2e55bd6f) +
                      (({q0_1[14],q0_0[14]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[14],q0_0[14]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e  <=
                      (Id27dfca888552262f492b81fd23b881938f66eb15f7ab21afb210fc6056fa09f) +
                      (Ia96c921ce4e0590c903d02dc69790c6af52898da90f4766121fa7b31e0ce6190) +
                      (Idf239af48228dc01198fdd7240b8282cf247cbc6969403dd994aeac0e5f81898) +
                      (I6687de5f8cb258492154a67fd3a3d5ee88d97a4db1c6c273ad158d5205ae3b48) +
                      (Ib924c4eaf872874debc3b6ee65921f0381331e1421cbfc3bd17e8caf273049cb) +
                      (({q0_1[15],q0_0[15]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[15],q0_0[15]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5  <=
                      (If53d34fa90e564a24f6e116baa8a7934ec4c51c5f0bce8160f0f389391792fe9) +
                      (If0fe01f34db565bf669e2df82579abb4d3629e8bb001bbf874b9b76f8f780a37) +
                      (I61f7e06790f5516eba113bb79388fb515faa1b3a3bf06598a07f534ce2845618) +
                      (Id6b81456b5d3050b4e1fe80ccc8f992cf56eb0f08a1d29ec1e7cabe1baeb0872) +
                      (Iaa0b6d0f2fe24db548975f410ac5b79f687b7646169247f3891ce9e4644ee0fa) +
                      (({q0_1[16],q0_0[16]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[16],q0_0[16]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c  <=
                      (I45ade5cafdcd254cc640ea8725da6961717fd6c50f747242aab6976ace4e8f10) +
                      (Ie2e727d2073eda2be7642a6a2937cd3c4e553d8bb6ec56d914231b5bfb12405b) +
                      (I1aadd9b378df1ab58a1b1af097539d1407636833d9c2d8b08c8f70be326fe199) +
                      (If83264f9ff9f7b77429559aff8b14fce54040210c6ba3476b77824c28b95bea9) +
                      (I1cf0e3016bbd2d8e5debffedb198273a2d019ce75f2f8352a285d17264d262f0) +
                      (({q0_1[17],q0_0[17]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[17],q0_0[17]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55  <=
                      (If9628510f239b2275efec7ce187b8eb7360beb042a425934ac81632815361368) +
                      (I7d0cbdb63988e88f9f3f69b35029cb2078b97b6cc9008644b2721eda7fb6cfad) +
                      (Iea2bd90043dd35ae24830a90ed10d12869de66637ab0237a1ad459fa916b57af) +
                      (I0f54db0f4bdec3ff62a8f1b5f4974982e3600a906dcfc79789fb9fac058c353c) +
                      (I9a4f77c8ba9a40c1b543070a42451ed37c0f22850a4734cdda393e69c7b54733) +
                      (({q0_1[18],q0_0[18]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[18],q0_0[18]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75  <=
                      (Icdea1f407aaefacb918babc28247d540a8a52d513d26d7fbb5e81a41797e7555) +
                      (I83ec3e2a8ec621acd2afe475255e144f2158e1941ec685a346b75fc471b9cb76) +
                      (I25600d0eb62c066eda0baba4269851387918088406d117377eb8bcc2e080e426) +
                      (If45b8fca9a85788040c10a47569139b44384357512af96ee7bd8cd98d88f8f0f) +
                      (I926233df0c5e8461173cedabbf49fead4b0ab577d82f2585af3a1fb6e3130e21) +
                      (({q0_1[19],q0_0[19]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[19],q0_0[19]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8  <=
                      (I979c6bc2b8486315e3db6888ef068b88396857d05a62470d4f3c33833cfde130) +
                      (If2b1e365b8ee6d4afa8536f5c2f5c80d31e86ab6729b26795614d75a6a18ef42) +
                      (I50e7a3df23a8147b9a87cb5e38d44bce7613b2a717d1e3a8bda1171f9522997f) +
                      (I3d6bb14416567aa7b8883b3d1778b55c251a22ed42b09bb3cbae6a5210cf11f0) +
                      (I54b0a17c9919d856bb3ed7cbbd8e42fd4ffa33ce8c32d45e4be1e28b71426ee5) +
                      (I4a6a17ada186c2bb60e521443c0a5a0248d03242c4ae01b751fcce4abe853065) +
                      (I33d759e40b55a0d83119f5c19cf87e6e3181c7e3eed94eec60fb52f9c376addd) +
                      (I84920b6036437109dbc48865b69f249d82da5c7288a7eb7744ea7ea567e03657) +
                      (I78f0dcc6533ef218ce6959768639c983d2119dd518e988eb3dcd6f0b4de98c82) +
                      (If64a23ad02d1da21fe63cb33f95d37c576739eb181b0fe50d7a5101817b4ede9) +
                      (Id4cd4fdc9fdb1198c2894543e212f665c925298f1c92b4da9c432eca9442963d) +
                      (I2e15c5739b990462c8a17b590fb7d60ac9c7e6648b79e75697139f55221fbcc5) +
                      (I294ca1e2c287bbe18783f7043149078d4fcc1c59e24792d75655fb29a36e33d4) +
                      (Ideae854591637828f033505e4fc9dee34d82369d02f7680ef6887c597ac1ac82) +
                      (({q0_1[20],q0_0[20]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[20],q0_0[20]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68  <=
                      (I597d0e1b64b5d47502804c7ba47fd0c17322bfdbd4d332b11f9742713f76855f) +
                      (Icad68e9babee274d9a5b79cf432d9e2a1938e06f51aeb564af6936972b3f8e54) +
                      (I15b5266ec781a5ae11540d23bf8b1a0b2eb45d94ab6f367a872885ff3207d5a9) +
                      (I5c1a09aa19ef4bb254881dd92543acf840270aa36ad4e0f5f63a6182a4c93a1d) +
                      (I9afcfde9391d485e865b08f9b8ff69cc2ecaace5f5e26e27b7e1775b625722c0) +
                      (Ibe932d914d189b275138de8d6f3ffb914940d4b2bbecb574fba3c6aed885c44e) +
                      (Ie2abebb2c2604e435cea102275e0726254ad91df1973aece477e1e5315f82d0b) +
                      (I8befad7180232073f2f7db5a3f546a5a1af79b21cc9cb00a13e266db4eebba48) +
                      (I3a9293b8f323c7e097a099fa6beb33ca299723796aec9396365d43334eb55e35) +
                      (I52698fa0d5291f0dc20fb5f24c33e968ea63f47765bb7d231720330b624b2fae) +
                      (Id8d0e36ce1faa76feb8cbe0331f2179ddfc066b70e93e990b5d5bce17f505440) +
                      (Iaef8ec1714d2faf3d3b947db31b7975161077ca31fee04842efc1f7159104d30) +
                      (Id8da43222903044cc48243a7bcce7864e66d151673396879258ee4af7008a706) +
                      (I8eb86c8d64d83d4ac46667af42b6383e4d165459475ec6be9d547a70ef0248af) +
                      (({q0_1[21],q0_0[21]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[21],q0_0[21]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b  <=
                      (Iaf205cfa67ea9b2c39d6705da465f081eb75c326c1d80e63e1331a098ca9a4ac) +
                      (I16ffb13aa3dfd9da5da39d9b2246d5ab46fd0fdb7c02781abf4d8bd754bbbdf3) +
                      (I9a15ed1b2fa413056071c97b4f003717902f38d29805752222c45cbb2cf58109) +
                      (I6a10084ceb62d383dbc5871a208fc087b23de418b2c780813ae950bf4e594c96) +
                      (I63f5ecb10fc3ed9bd8bf79403afed8ab1a70600ceb1e755de0d44af98495ea88) +
                      (I377aa224e1817d2ab5cb02a5a290a723621782607fcd59b319d8cec1b092bc1b) +
                      (Ib1310cd21337a1faa061ffd12a2670171f582e03471ab315b90de9f8fc30959a) +
                      (Iabc9fc6e9581216af19559d8e709ea0842cba4f29f3fdfb05bd71d6d9f7594ae) +
                      (Id165331f616d7e8f347cbe46daff955009fef6f8c0310c64c01dd35990231279) +
                      (If17c7df712b5dd40132ac60628bd514bc70092122a0cb89ba7d4559439779fc9) +
                      (I9d7506b5ed3de0e32e821ce6ddd1c28aed177910ccacc4d4aa2a8ee57212d162) +
                      (I734136c95a40c62745d684fc7e8cd1114b883c6209df11cfe01b9174cffc720a) +
                      (Ibae97ff31fce14dd0506fdfe7407fd6260f7cf8584a01da77312b1aa48594be0) +
                      (Iea011619fa5b0fb7d22dc4bb4ce3fcc4856dfc7286ff393fb329ac0d7e348207) +
                      (({q0_1[22],q0_0[22]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[22],q0_0[22]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e  <=
                      (I954e0367a6f3af96a7e033da51e7256543d7eabd37191d4b03f3077567cb629f) +
                      (I1e6d7d9769dc32e1e014951538f1cd1014e9d07b675e6369e88ad5a6fd400787) +
                      (Iac4172f940fcbc93db2047b26fece588f3fa63ef255ef404beb5e6ea016b2ba3) +
                      (I0e9a7c6c53b89ca2685615c270e8ef3d3f51fad8619953972e1037edfe633834) +
                      (Ib99b447a19aa10415461faaa8d8026b0073582bd078930f2cdf0f531259d9c50) +
                      (Icd30277c9d839d833f27f571231dd138497796d3e7818460d836a48b87e34d03) +
                      (I2862bdd9be64c24d98e80e8b662a7c97c70943bab3d49cc8d39443abcd5c2c3c) +
                      (I4f73c51d25db7485bf4a0d63f95f14fc0661431870ce704f70cbb787eb336f09) +
                      (I2647390c3800518f2251794a7ee4aa2d71ca9589534cf73eda0accbd2b3342da) +
                      (Ie05c1da46b594d3c94aac179f6c98334d0d667cea08108719b44541b7b0a2049) +
                      (I1bfa3da571b0e3d943ec7b9a8c641283e080bcc6502fa8317ced3c0a6eb2c4cf) +
                      (Idfa7c6c8248be1a2f8a95c6c74a71be3126e039a31f4e16e0b964476c6d47953) +
                      (I5c43417b1bd96dfedeb36f6d3405fc7f6b73c11a55f21ebe6ffd675e991a13c3) +
                      (I71f31c9a9943d9fd422d00aa01888aac32dd8b34236bdd9bdf3e660413a3512a) +
                      (({q0_1[23],q0_0[23]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[23],q0_0[23]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a  <=
                      (Icc43ea934f0c07465170977b52d2f402fe155ef77f3ca27119fa665a1d918694) +
                      (I78abc91706fec0893eee10a69916f7247b718169155038bdc0bb6f8661ed1c3a) +
                      (Ia428f915c49f84567006696ba3f5c783035325755b4fefcf74d65aaae1f3d3c9) +
                      (If270910122bcee1c18cc592dba9b38c026f792d8d1472400a09edee9d7633e22) +
                      (I1517acf28729695d689aced1c7eb358d9acfc4453fedf95a76fc22c972550c63) +
                      (I8ca8dfb7a3a8ecb9eac34d1d1ef4768d31b86a757cb7b9ce61ef159816ceea7f) +
                      (I2cb1ae23e53b89ca0fd3d1df98b32d5b9e478e9eb579b0875981a6b056e8ef4e) +
                      (({q0_1[24],q0_0[24]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[24],q0_0[24]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0  <=
                      (I1a2646b8251f83855c3fe8f6172f36500201ce43b9b5ba2cf0f25fd5d540e89c) +
                      (I1d9a8ff2514f112838c7e4f568303dfcac3f86d94003ec4f1a40a35b79ee8ef6) +
                      (I83c8ad082be8fe1a71adac4f41a3bd7019d2df299d19f8e5a293367e49b04fa5) +
                      (Idc29625b375c44e890e371217aaa25d5fda337ba8177fcceca881adc72292a3b) +
                      (I6e88f83ef5bc5f950a4bcb904ffede2603201e72e362aedb8db04412f7bc2bd5) +
                      (I7ff25e517e328eda581e7637a2114a7cffe873df520114410c0487e503c01aa6) +
                      (I463662fa980f8a5e4be086aa5f37db53b1d6ea8dfe11725b8c407f779a168998) +
                      (({q0_1[25],q0_0[25]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[25],q0_0[25]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4  <=
                      (I8db02445666e4aa12d7e495ba28ca0eae6ef411094d30330e91eb9eb03b38aa7) +
                      (I8c971b4c1be575fe328c0a4a9ecc5dc75f08d36f65aa58642976d971a6c316d7) +
                      (I09e6d011dacfba2800f9ade6a495076a67e4acc6a944fd649a7c382422e8fa6a) +
                      (I76599c709cdbb3f3cfe4071b96fb7dcdf8e072fe85ad5c8e7bbabd4f6182303a) +
                      (I0d9bc57dbbebd429ee5a5e5dabc1cd0bd9f4de95a920346b9e61cee83969ba0f) +
                      (I91716015389a9d3b1d0cc77327f439e02e54be0d3524b2cdbeed886eea673b10) +
                      (Ibc3e77c4d6cb28599b7a21c7992802beffb168f54d8dfa650750ffdc6730df29) +
                      (({q0_1[26],q0_0[26]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[26],q0_0[26]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e  <=
                      (I34f861f0a748b0ad1550db8ce40149dc638194b0089cf22e2380a39a49f8c902) +
                      (Ibadbb4e272ab1105914763e2790898c8e37a553a1b6726e8818431bf5209b369) +
                      (I308f551a8479d066b2a4b473206e8f407082cf83b37a376e6b0e1454f7ea2635) +
                      (I58c6fbcd5f77398c3514e6a850bb69d9f57880a387f10132aa63079c0a1f4857) +
                      (Ia9d25b6cb880b9a00c9bb27bdb80c08988eee46afccbd578659eb98301fbb8a8) +
                      (Ied710d5ba03554d4103468029a9d895c25c10765b6e3d73bbdebc54d7cc7d8db) +
                      (Id7dcf87d2a40e82e7f01327d834d5207ae5873a7e5133c3dddead9d0cb9703f9) +
                      (({q0_1[27],q0_0[27]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[27],q0_0[27]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a  <=
                      (I982c94b61dff8249f2f3055f60da6e2c2b0b56c403f151168b28a5a211aa6428) +
                      (I710a57e6c5c8e228325430ba2a5fc32ed9da101d76ccf1d8c9f3397859b39ef3) +
                      (I2cb87b14b006ce6a36ee5439eb18a4287c5b9ae79748faee259c0435d0dac81c) +
                      (Ife00518e7b24a5de694b56a32211898b3c23d2dbd2df91a4197216c23fb5aa7b) +
                      (Ica9ef16b19711ccdfe32e34eed347b590635f1ba7983272eb02f980f80642254) +
                      (I9331a9d6610ae5cb77aa3d477fce0c0ad7378a884c86c4872a1573f2d8a90d8c) +
                      (I48d9ec419ebe83e2a5a8281e7beac36acc9e554b86b154736dc51ff940f5348d) +
                      (Iab97067540ba8c9551711cdbff0c6aa3993534d3e8b352bda090a0997c681afa) +
                      (I25c667a6616c9a94f6618166c99298b28d897f9ac8276bb85816e4b42582cdfe) +
                      (I2d2137ac29a7c23160dedc43e9caf010f72f7d08b057e49fcac89984e616fa5a) +
                      (I11775c069ab4acd951a3ca47bfa65c7632a6a8a369bb103d0bb719806dfe0c57) +
                      (I6e418efd4b385b2a298c1c53d344e35f593e8380d1c27d7cb62cfe35223121c8) +
                      (Ifd66abca1532f04fc777617d91cd2d5f4d4fee35c3f075e91639a196780168d8) +
                      (({q0_1[28],q0_0[28]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[28],q0_0[28]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2  <=
                      (I6dcc482b16866339b78b922f9a7ec0f4a0ef311c353e6a4e107dfcc351abbb23) +
                      (I8c8bc477ddc4000dde6459d7cbc4ba665fd4ecd97242d9f9fe97ca6825bb033b) +
                      (I54da11ab334a3942047eb5953935aedd00ef1a24bb5361fba51504632ae61831) +
                      (Ide2ca364c5742f786e5408980fbe12322ebcc2920fd99ed322112d3623d9e372) +
                      (I6024b75d70e3da7df4e532e712df56a8bed06352ba0a545ec355f59473929d41) +
                      (Ia79355adc994f77e150b93a3e38c8bd6f0a5848a212ac64559cf1210ee0d11d7) +
                      (I1b68e82cfc8606d3a9325ff2da047f345e2f34b44eb428bf2a3bdcf42a6e869e) +
                      (Ia1d4bd5d90332afbfaaac3cd0d8f5fcbc626ec4adbb0b0f16fc80923925f703f) +
                      (I87af49f5f04df14686aef62aa27c16723af3ad05398f00e29788666b27784de5) +
                      (Ic1211f3a0703e281ce073a20afbabe9b2a698d1cf74f07f099d21fd89ffc8908) +
                      (I2985f4f17b726f40ab6609b57a796727fe46605944c5e25c594caa8dfbea9f58) +
                      (I6f7aa66db409365eac05a200d0a0f1d2b25e9c37ba4a7db3b58a7298af0fd6e6) +
                      (Ib1e319af12dcd98c09841e8b06e7af86f2569bd7afeb1718bbbd26e30f65c464) +
                      (({q0_1[29],q0_0[29]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[29],q0_0[29]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc  <=
                      (I30e28a0e32497e3137bb689fdbde46389bc490300e15be88612f28eff07976e6) +
                      (I0b525cae7fe005cf25a07cb0b1486152d726fc74aa55f03480f10af97379953b) +
                      (I3df4fc0f2f099890a34d7b376328da6460d429e2516a5f8fd1aee5a8fee835df) +
                      (Ib1b15c9e15e963cc4f2e9caa1b6b132e338947224b705b51ebe710d7e0f661d7) +
                      (Id364040d3b9f1ebf34ae3fdf7465d955b49d7a2f4709219f76229766d6df98a4) +
                      (I7cd9dadb64725f4217f1330c893724a7537a616ef41d9dc49fd2794125e0dc3d) +
                      (Ibdd77bf8b31352e365f7e6440a57247a8ba62e667b000c1347165bb39f3c7c2b) +
                      (I35e7fd3f09acca79a1003b0a4b7ac62c4a2be93bcf333abbfb13a5eefd7d5eaf) +
                      (I7e269b2e2d9ec70c47570bad75bce0ddf53e85e3cb4ba87f784ca520c5ff1084) +
                      (I0c23517b9814053cd1f89a8b80a64fcff6ae65937dc97199c0b79ba8f7a34ff3) +
                      (I73ecf8ab6430c6343bf7596e671ce01a3e3e7499813ed75c583a7103147b0bb7) +
                      (Ib7f659da098e577e33fc0f5da1c03f6d3e68b3883ad7888152d2e8684a6177f3) +
                      (I3386ee46348e8c4359b1ea2153bc64afbe76f2b6bc9a312629b8c52762a22873) +
                      (({q0_1[30],q0_0[30]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[30],q0_0[30]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93  <=
                      (I8c2fe0c8cb55f09e4dcdbaa3960acfd815764161f53c6234273dffe4558644cf) +
                      (Idc64cee034c1ee132335ae593844b2c46e3f1b1b2cda8699940df311735a32a0) +
                      (I1c7699448a10638886eaa021495d4c7cc378fe1e9b0aafccda001c15484b9419) +
                      (I45b03b0185f9efbc11c707a64fda9203cc82ec2fbaee7ff34610c74d7cc1132b) +
                      (I3097f16921e899a99f2a2b013a3f6d339ac9672fa5e17655ceba4de2d506e151) +
                      (If0d62663c8a08719b83a27c76fa62525eb14d452d4ff0f33e94c67f58d7c86f9) +
                      (Ifedfb1db4b16b86149f5eb8b0adf06499331d423c368c0077c738a190a1814f0) +
                      (Ice24cd0bd76a7d12a0199df195b34f41f7f72f037177656693b3154d102ba729) +
                      (I6148a04ce3733485aeb6c4d20b6117eea37a510aba76ac29e82d44980bec0934) +
                      (Ia6391e6b0ad4d9fe4136b90a57d121f2b5f16ed4662429f1b85677591fee37a6) +
                      (I5dfc39b913b8e0d00491e3f7f45b6b467a517b5e87baa065097e28e6d695500a) +
                      (Ie538f6d2c778992e2324a9adbde215acaf7b8dc3a72a9230d4fba2332f3cab67) +
                      (I03929e638a59a35fc0168772ca06f7a502352e03525042ce6d49cf9ecb671093) +
                      (({q0_1[31],q0_0[31]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[31],q0_0[31]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d  <=
                      (Ieb5e001b45961175497657da7a0340c2a15b6d8de1b72ad68ac3aa7f96a47af0) +
                      (I6d58dbbb9b18e4b347b34e548c70a9bc0d819986fb3a6bcc3ff8a67c1fce9c9f) +
                      (I82772b528a8c156f2932a23a720f8446f3062e9605839897b4652bb2936fca1d) +
                      (Idb259e613b71ccde839570ff2e7f21a9cb7bf676ffd4aadfb08d6a963bea9640) +
                      (Ie9b1b4412060f1e9acccc1f3ff897bce33f24fea3bfc91266f9e42c1f38aaaad) +
                      (I259a9b6041f341013e6ea0706c4e9ef9a77148bc003b3f0cf9593ebd915b30c1) +
                      (({q0_1[32],q0_0[32]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[32],q0_0[32]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6  <=
                      (I41a57b30ab1dd9c40a723f99315558a47412465aa3fe967250572e8373aa7180) +
                      (I42968c25ee2870f891f69991ae3ad8bc1c3acde2f8f4d6c0cacc48f562399c37) +
                      (I44103a07ffcd818c0d9280b96ba08c32f96edc83a981ec9748ed3d6e9c061d62) +
                      (I1c886223618a03ba9e18de68462ddcc522338cd26d24b5e126da9da1df1339f4) +
                      (Iac242fc0dcf37a86cc334319d77aaae46dd223017f2a6489c4e33314eabc9874) +
                      (I3225ba7b6d0e0c7a94dfbc8e074ade02b79a66f6aaf97580a451c2d1781a625c) +
                      (({q0_1[33],q0_0[33]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[33],q0_0[33]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab  <=
                      (I25779b63a47c05d4588d4b33fecaff61647609a62fcc90f0f541c6b30ea9342c) +
                      (I05bd9a1d7818f4945ddc448149dee571e80dca8b6eba7ab79b17b6f84d3f35f4) +
                      (I17eff5960d8d41f0832a48fe9a3ae0dfeef1bfc44b73eff506fe1d3813398d15) +
                      (I1b02edd5d00090446500b1dbf66a7e674de978c068b81ff0b0fb7abb9ffb1654) +
                      (I2c865426b0f044469b391bbc13f977fdd19dc89c908574ba289388e382d55cbc) +
                      (I2e557a901de23b8442e8002b3560bbf9cb8592b7bfb7a6e2f8aad12843a5a041) +
                      (({q0_1[34],q0_0[34]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[34],q0_0[34]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727  <=
                      (I469f4965961eacfe3dd0cb82fce4905e19e6695d71bec95956e8209d2ae39ba1) +
                      (I6e148041c3612c795f1eb1513a9eba29e0509f02f94971fed189dd9f03d54a4c) +
                      (I2f687e6270528a72aa2f9f9cc0a5a6368f8eef358270329cc40b56abc0e4a35e) +
                      (I661bc8acd80497efe43e3d6fd92bc4107b1ca63eaf162cff5695b35f8d4a7e26) +
                      (Ic72f2f8a61b8ecf8960d476bcf8fbbfd4389e932377679286e7182cc12c418c8) +
                      (I823e337e6437e5ba36ecaf0b1ac6b7a4e74cd2ed7019dd5447355626a8877d89) +
                      (({q0_1[35],q0_0[35]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[35],q0_0[35]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733  <=
                      (I1622b11941b00f6d2ecd90320158533a66501a6ddb78defb4464a937f132c232) +
                      (I9ab473d34fac3327f03768e14c7bb20056aa8a3dd31520d385552eb6d214f890) +
                      (Iedf1b21de2a0eb04c4a64f9eb34e2b0b3a152d90b1938b61ca45c880eab16ab6) +
                      (Ibe3e6de02f0c30287dd89b07be5254ff70d9683389574d02f1423e792bd2d534) +
                      (Iad8ee4f6cd13a9f415cd3519de0179a66cfc993a840b3101cee554b55c0e7e7a) +
                      (I15123100f4377e14c62cf47fb1fb652badc3bd0e8f0ab4b970a0bece065a6380) +
                      (Ic0a892c18037ef674c8d94cdfc94cfca47d977ca2da9e678303255b96575f022) +
                      (I2c316e8b8cb6b499a7a8fbb513b3067829197cfacee877c35874a2ec686ada4a) +
                      (({q0_1[36],q0_0[36]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[36],q0_0[36]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521  <=
                      (Ib3a2af9bef5f5d8d7228a3b49a5e0d4a37a33117e057078a552588a24d46addc) +
                      (Ia042bc20eb6866de0ab9ca9154f0db63f7d4ad84d553be858a0be88fbb8f7f33) +
                      (I5b4ba308b0fc2946fb11b66aa5c24c7b5cb2a21955116b97f3790de65cd2a064) +
                      (I005ecc3a38317079c7bc5008817e11017c33671f77364ad9a07d0eff1e0ebf0b) +
                      (Ib63856036797d30e60f13453da509ace15e3324c25bdfdea5aa495d592e2006a) +
                      (Ia9bf10fecfe62530ea6be4687ecf78a2ac08c6fc6e38328c2d64a80cb5a3d72b) +
                      (Ie1447c9e1eb4ed110e6b0353bc5dd2cd14ec645355c3cf897df6f6c5808475ad) +
                      (Ic8f640e7a0c71ddb20a985259b5e48746d28d2898383765c3b78c577f281d27f) +
                      (({q0_1[37],q0_0[37]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[37],q0_0[37]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1  <=
                      (I3b1d695a626aefa8e5b146c7f7f26a8da119680783da7afb019209ac9fd719aa) +
                      (I1d91c7e9c2f99df4e0523b7e01b6fa6ea3930382238ccfbc07201b7d3edcc969) +
                      (I7c1e9623dc53c8aa8611b46c0375994510a97c4d49d0b091964cbe4671acf1d6) +
                      (I1b5d096081c0190c0ce6a674de1afee9ccd766a9cfab0637a0aec33199061bbf) +
                      (If145a331c8a8abde8c26d2571cc8b38e1eaf2768a4658d350cb602bf8614a521) +
                      (I86e764dc3320206d9b52013c2d735ff4d27bf6e4a82227486e64b4ceb68dfe8a) +
                      (I4a98524c02346f4b9468666ffaa9d996b9b868a5a8730264d798d7a66b7454bc) +
                      (I1187dbcc72f33b4cc3442982af526be4cfca1b5ac65be943d4ec380421632117) +
                      (({q0_1[38],q0_0[38]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[38],q0_0[38]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709  <=
                      (I73ce2860dd9aa9ca2c0d541a6ae1e5069badd35988d922cffb6aef0038cde662) +
                      (Iea2dd4d33966d53ae739a16876ac2cf04e1d95374a5af68e59a5703dfef2aa79) +
                      (Ic0a386f5301913434a3d6aaea1d56d6acb3484fababb7b8831d09563bd8842cb) +
                      (Ia8a4fca33add1c3c58b04eafe9d023751882f409c5d2905f77aae3fef8c2b008) +
                      (I9cd4ac82c1e6f2dab27efa85314df34a40d8747959eba18330bd424a38debece) +
                      (I9bcd5f3f4630ce7a24ea4479c9ddfce59ed809dfaad9d767e80295c41b332f4a) +
                      (Iac7a05e270cb898af4ba32c16445d0dbdffdafdcc5fae209f09367abcff9d6b7) +
                      (Iad7f008b5f08f3ba94a0832261fb4add17f0897e3c7d54a250377b813e284331) +
                      (({q0_1[39],q0_0[39]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[39],q0_0[39]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d  <=
                      (Ic072a2fb2ce65ca734c05e747f12ad094cc5aaf9267dd94dba345b5c7b11dcdc) +
                      (Ic20328b806ccf89387180fe6d88ba762051c6bc2c7f82494129e8c3600108804) +
                      (I11855780f53e8711f8eca9370af31f472dffd126c02cfce8154a959f33c68af6) +
                      (I39b8420e976cbdf011232d83446a5cb92c2ba58577792c9c61dd71358205e936) +
                      (Ibca01267ba9d7e2fe9f8df34a548836390ba12b9b782f16ba40965c00735213a) +
                      (I105a7d84244a0d9143b9b2a3c64ea6964f7e1f43b7f8f5cb15d579885bbf746f) +
                      (I1b0f11f3bca53713a53e2ed18fb81f5a25c7151c874be612677f5204bca28093) +
                      (I434991f7c09dac3a7bd42fce3073dcbcf8b1c6579822074548ea94fdf1ef4eaa) +
                      (I7fec897140c79264b7b7b7f3ae228ed090ff69351985c07d317ff9c0cab1e58c) +
                      (({q0_1[40],q0_0[40]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[40],q0_0[40]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7  <=
                      (I82bc7aad8e3adf5b7bd03d9fdac6eea60cb800e4502e3af7bdc9d49139563fd0) +
                      (I218ab164221d559f1e8bc2a13f06a7593eb4133134762698eec270be5d4c3906) +
                      (I4135dbaf658fb73b41800cd275824d1c9f410ab1b6e555b6c4c8df12f96c5861) +
                      (Ief38674752576e92e90fbe2a7abcfc952274123875a95657dd42c910133cccde) +
                      (I783b89f0c1e5463646e0fceb976f2b27aac523a677eff6e597e434672b0daac1) +
                      (Ib0ee967a174d7c841ebe71e144d6303bfc80a6083ff6ad745c76d488dea66d9e) +
                      (Iea7b69c43ca4b3707d3bfddf19b27616b8686df915734ba86d3685127bfbf39a) +
                      (Id36acaa2c9161668c95e2cc3e6e852e9243ca7f486ca6c2ae4d124b1a8ddb522) +
                      (I325ec6d7bab5ccd6e9c4a7e9b02a3b8c30072df123bf6318bd97f1e8766457c8) +
                      (({q0_1[41],q0_0[41]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[41],q0_0[41]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499  <=
                      (I07c37e958136be68b3d658649964c73ca78160582248da1d45eb9ee82c1f679b) +
                      (Ie17e17c22c7215d0482ba310638db13a96c0943216f9ebaf53c0c29c69971b23) +
                      (Ie44aa17133d02266160c8fd6f75716f8bc4a3775356cd1ef0f495b13145ba864) +
                      (Idaf1699bc7916d99a2a5ce0174383c189dca6d7537734b19dc379bd634d0d209) +
                      (I64aaf806ebf0ead2a4836251dccd62a394b984823592340be94f4ea02e12d766) +
                      (I152b3a1e710e5a39bac6338591c6597ee2a38fc25555f563beb7a1a967bf4e94) +
                      (I9ede22dbb56f48c045a1b5a05945124fb97b6ca7e355dd8d9dcfdef6e623b953) +
                      (I30e30c2bee3bac86dd68fe8364f818ab63e91d65c4fa1ef45fcfd03c9df87cc5) +
                      (Ic0bef9008769fe36d726cf80506004d66e7c843a046653201c9bc2c816115c28) +
                      (({q0_1[42],q0_0[42]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[42],q0_0[42]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b  <=
                      (I252a77c3eaec2d6accaee6de3ba5d0b354636e2a2aef4992eca0e2a74eb4d25f) +
                      (I5fa628cdc28fdeb96014a4d2c2d06b092136cf2a14a0420bd5d3861b83687413) +
                      (If258ff7e66143201e30b3fd451e1b8e2ec9e46596c2653ec836617c093f28018) +
                      (Id160a3b60a3c7a3ad93044461ade9ccf0b7a627efa4b1bba84a2ea0d4fbdb551) +
                      (Ia42e25bf722566321268c83de181d196619f062381c7fdb381ab5f6aeba6589b) +
                      (I4f96b4022f127e7d965786f2cac8ee6afdbee96980608c876c6b699495f80b0f) +
                      (I6a2505f0de03f3e2d303fd207ee819f5a1777b650930b87a235ab3cca5de6e87) +
                      (I8600d4c5861319be0efba19d9b66ad483aa7bf648f2132c1a339157c43920c18) +
                      (Ic551d228c593c4304b4ef79a965ac1d9081774282af09d79cd587ef9abcd6003) +
                      (({q0_1[43],q0_0[43]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[43],q0_0[43]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29  <=
                      (I01d7d3d20ba0eab63d519ae054b6c22c5be4000c846a6a4883ffbbddee37663e) +
                      (I4177cb2b0a83442a271f59bf4f758851d5146ee00d76a1177c9a34d4208b7c09) +
                      (I5df828301af902c72794032c0e55d8e7548c9b2277b2edc77f53796ff8e04804) +
                      (Id595e96924941a80a6ade8778fcbcef39b07a62fa1d7350fe50182fdae302556) +
                      (Iefbb3d08b0b2fc51d2f6b60b25b8143f3f88a705e770396e2f6d050632ded97e) +
                      (I71c3a88492c33461f93d43680f11eae8ef3e9402a4b931c5d31f959a2f8c147e) +
                      (I7a7bbb1d7d9b77199c0b29fda08f8a63112052ffb0a502a05586ced336e13c62) +
                      (Ie1657c5216d7c6e743a23819c08b7c7f2fc8a56793e1bc67fa5c5f3b37976641) +
                      (Icac36c9706c9e063b771faf556f6699e280687be228aebf6ce71f5ae775a9754) +
                      (I8b3bb7a4701d3ef22c71a9631482e13afc2ff80f40e2f0ae75cb2211af5ce6d9) +
                      (I6a24b9c3ea194d09d619dff007c4c6f53a3cbbbae5c9d3ba718bc3546eaad989) +
                      (Ic7af968d25c444d210ebbc7ae563688f4f8a48f38035ce5bccee100e10555047) +
                      (Icb61d0767612534695d9de0380a1febbda612604f373afa55f0339c7a679e99e) +
                      (I58d2fcb7085fddc9250ca075b010afdc2d019c4091f5d115d9520586224a1ae8) +
                      (I4e5dfe1c7112e24769a5e6aa86584c09ed659fa5d05af38d18183db31189a3a7) +
                      (Iff97998b0778cb649d03228ed3acc81c1b3a97f6bc47041c423120b1311112d0) +
                      (({q0_1[44],q0_0[44]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[44],q0_0[44]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171  <=
                      (I422fb05bbac12ca5df13eb7c0c3fd96a4e819de9669ccd64d40060b5db3f3421) +
                      (I782d29ca9e53ffe86cec8809d7d413c9c5ebd9edb6a0d76db2d0c321312d224a) +
                      (I0705e6f1954b14f35dd7fa8a64370c2f9e6e39b6e265857e72946815d1f994fe) +
                      (I3f9e2f1be98a5d14a8b79b252e9b5a2b3a09304f27a3526a4a66b365b682787c) +
                      (I134dfd9d579ba8b2d72bf1c47119a086fcfb6b7d591cc2c5558e451f57636d0c) +
                      (I5f4870fc880aac0f84130a26e3cd493954ea49eb3804dd17a91b2ba1cea599f3) +
                      (I918037e81d2f9c05c6a8b94c64724b1d0ec8afafe5666df433fee3e296171f54) +
                      (I136f70cfdde5473f8944efa2b1093ed76f82dd06a341413ee2a56054ebef5fd2) +
                      (Ic02dae50f30bea04d63949eadbcf892ce936efc5373a6185668a20311dd59f4f) +
                      (I54296c97ecd9a699f171f4d7271c761aeea50255010a0a90d2dabc16a0cbef79) +
                      (I50a310ea41e0637bf28b5f56cf11560bc936e15c73acee063c60668bfa905fed) +
                      (I25d2b0d3ff7f684e508a62271f3d29c729dc46478248627013dd91075f8d2146) +
                      (I7f9f83601cb61fece60f94c3120b43ca0c737ee36b8c67ccc917d3a428d8750a) +
                      (If4fa37977e1db59d1bd7a30b2b0919c997b6e25e0438e01b62dc273d10497867) +
                      (I66291192ca8d81c8e3f667651d5201cb41b6872f73283d13c6718159b008d8cf) +
                      (I4bfef3f43cb1a77ce8b2bf4b26160a161e7f28308b8d2817e6e2840f09463e37) +
                      (({q0_1[45],q0_0[45]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[45],q0_0[45]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4  <=
                      (I0aafab9f9205eb4a8c16e213e116d949a5c625f7cb2b0f3d124deb80aad2c6c7) +
                      (I9095fb177f965807ae5a73a45c76b1c0b6300c6800b17259e5836adea5a78ec8) +
                      (I3780e5266741d9a9435818f002588f4c44ae518b77a30ede57a3823e1e1e5867) +
                      (I360ab21cba3dfd419f0ca83f85d9633b918c3d24a00214399b0465d7106466ad) +
                      (I2c061ca6ba4299d676b5c6f1e1cc920bc1104e7ac730d207949b952d1a98300f) +
                      (Ief44fc6df0864dd0766877e0d673847250f53ab137cd9029916ab7149446f9c2) +
                      (I353e1673347daf260e61fbba813cd14f83c52ce3f6e5168c0fa6308d41e93590) +
                      (Idf77a6217d51b2439f71afbf5956a52a241f2bf8722f54cb166d83c3b45f6721) +
                      (I8ea9b55580c15fa584fb934e010debd92e2e893630de456e85036d583921011b) +
                      (Ic36cf3da50983e4168cc0a31ec0a86c171714355c0fab18398b8daf57bee1a45) +
                      (I7469c1791d81d0924eb0faa6303565dc78fe9eb371fa13039ff89b92b7f51a6b) +
                      (I9b8a4dcee9668bb71803c25e0ece0eebbf704eb29cfa7b91c47cf48d61076803) +
                      (Icf4d3544466d430d71abf2513cfbc16b575af540d369d405ed831753f304673c) +
                      (I0568efb50e0bb85c39c9ac6d2ab3474ab38799257dac5693085eeb0d74859ade) +
                      (If072f43c0b06c41c30d9bc40dae674ad9052e5533b1308adb97cff2e03821bab) +
                      (I2f05dd0209278c1e661998552da73728c1521c024a7d26f4652d4f151c6e5f80) +
                      (({q0_1[46],q0_0[46]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[46],q0_0[46]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a  <=
                      (I17dbb17fb2770beac552dafeb238c5e8e7a948c35c7c543508e652cbcda01dee) +
                      (I68ed84b705e3c00d0fb66182d6eeb93f43999532d713f81fab39a36259e0e7da) +
                      (I9d1a378e4d5703b65f197cb76a1982cc10e0c17654eabcf10d9df091086d8acd) +
                      (Iba503643311c9dc3366b9bb843dcc1ee2f0243c4cf78004a660fca224b36c5f2) +
                      (I05806fb5d45e4d6f569c12116644b625b7ba071eb052ab97525f06fca03dd88b) +
                      (Ib2630bec8f9f78489ca6cfe0bf25746b720aa422b9d529d67d6dde2d045d9c3c) +
                      (Ic57569daaae5eb0e66117615c8c6043b5f76b114b5c34b0df50445f66a22849e) +
                      (I5cbbcfd1cfc35b3e78d01b29831195106ebd9ba5907f44dee6761c2b047c4a60) +
                      (I6dc5ebe003a649f0e4106dc27f25387651d43259f0ddafad10411795ee48b40c) +
                      (I238a5c9cd1dcce0d745817081a4b240f74de3de6f18a3abcc42cafbb19a0ad69) +
                      (I53c29303c76ac3c1c02fc9a74eaff9595153ba06d67c08e07790c58e53b674f1) +
                      (Ia92993e9a66294adf7a4dbe1ea88a9e8be6367da1c05b8df343b3c7a38bfd8b6) +
                      (I329448311438699d3d590bba6ab4bfc9cead805f96015b77617f42d957bde7d5) +
                      (I717aab2686adb8a0688009c23d92aa4475e240ec0747735e6fee5e196a50c444) +
                      (I13a54b612481fe0fdfe8b52909179bb82298c2bff4f10adc4f41215fa4396311) +
                      (I26a27b64a7aafdbcf4a6d058181fb84e0e16767f4bd7a9c45211c4c1246d3b9e) +
                      (({q0_1[47],q0_0[47]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[47],q0_0[47]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d  <=
                      (Ie46448d24890ed6ffa2736abb97331dc3ed219b9324bc0e8453eed6aa2a4806c) +
                      (I8ab86da421b01a03999daa91e41ae95ff58c6bc38566a3deff72633a5ad1cc18) +
                      (I20ddfee724da47731a2062b2732598b429c42f7d22bcfb300dc084de362a2bdb) +
                      (I8d8dbd62189397b5e9189ead2126a615d5b6cea393901e21cd89c255d6672615) +
                      (Ie79db7f22cab9cd57482ce0141d83d5c1ff720a7c3dca2c3664feb4a1e2f4850) +
                      (Idcdcb2dd5e2f2aff0d7b362ddb4ae1ee4db08edc2c3df3589a7143bafeec0bcf) +
                      (I525b9b85b14df7a6533a7e54bdc9bf40a303c890a4a410251c8d556d38b33125) +
                      (I65afc937c55081dabf16dbfd02eb03c97204efbdcfbb523609571bb32d537d5e) +
                      (I45a11cd2f581121ac03fe112ec78bd07c070673712fe6112a3e4fb4eba298e27) +
                      (({q0_1[48],q0_0[48]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[48],q0_0[48]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c  <=
                      (I9342de9fe82f2273da138f99da619acf144edf1f9c33682fe3b1a09d0121c4d1) +
                      (If6cd81d168d83d5f6a7ca18051bbbcea5c7a9e017cfffcf72f31f73275c3a4d4) +
                      (Ie2c7966ff2c1e84a7ae016f31b0f8b9ca7aa42eec03467c7e3dda37dc34f070c) +
                      (I468b28bee4fe1c0d20fe7abd9338bf844ce0a2e322ed6b6de11e2ac621572c48) +
                      (I08c55e08731cbdc9703e607b481a65177e7e1e242fdab9bfb014964bb0d1d22c) +
                      (I6c252caff8f1ab047efc25a950ce3e3ffb47a5b779e37a667c48bc1487528218) +
                      (I2ade6ee1b52da04fce9491cad314947a07eb9aaa8b0a430db2f96e2d290384dc) +
                      (If6e953221a61b86b1fc339b69af853f6ad538b60770f2f7b880d7aa15bd625b3) +
                      (I6c6885b180013a16955ddefa0dc75c25ac85fb76059df9bf8b63af72c8c1fb4d) +
                      (({q0_1[49],q0_0[49]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[49],q0_0[49]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757  <=
                      (I907aa3f6584035b934017a601019d35f353b3f99c7573bef60fad167f9d9ffe0) +
                      (I7ae7cc2f052d37b650c0abeccd841b1b18abb4049c976fbdbab72ea579a5d206) +
                      (I5c0776e9826af1a98810296a7cb86adde5b1b41c434e6040bc6a5a30172d1bf7) +
                      (Ia244be7d571a1e41348c37534a23f7cc942b689cbcd5dff8c10043325b80e322) +
                      (I14730b2825dc07428388347472491ef3abe06da3bcea9b7dc9c919079c22325c) +
                      (I22670670d7018cb361ca0ffd92516837302d5528c26915b62d22505471ab7384) +
                      (Ibc34c6979b8f5adc5421ca8603b6dca91161055286758ac10d0c612263077758) +
                      (Id39c55c4f0df8a0d8ee4f8b47f3de8cebf5343bf75521edfe38a695565eea926) +
                      (I06a5cdf2e430e40b5c08ab617356f6b4b0389236041b77e2a57d9d314bfe77f3) +
                      (({q0_1[50],q0_0[50]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[50],q0_0[50]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84  <=
                      (I22c3d90c4ad5f41054f9b3dc7ddae143f567182c7fc695c5cd087f126ccdbcf8) +
                      (I533d6897ed500a803f6f6468e36a2a922495b3effbeb405b47ffb7a5f4d82c89) +
                      (Ib8d3655f6360b2b189b79353d38c9c9989af811109144d45af0f8b68a3276149) +
                      (I6b264ac5221269381b155a30c051523f4488ecdc6eb2cf60da80a8b84c49bd96) +
                      (I5c3a945e8bd4c55e9cb38d19100b13668bd652bc1162d16b30f1562a6595a032) +
                      (Ief691d56b56a000651b0a4c6cc9f26bc44da82f4a6382550d96ea4101b81ecb9) +
                      (Icf55933dce8b9f95a57d7d019c9b29f72e08454428013009cf0e4d2c5b6edf0b) +
                      (I5b0da0701e7399ca2e668c1602f494f41127e4c90e6fa91632da0016e7b395e9) +
                      (I6106f96669a63f337b78a6bad5894881230f0ab6467c23ec877cf27a5bc76cb6) +
                      (({q0_1[51],q0_0[51]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[51],q0_0[51]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc  <=
                      (I566a76fd27d46125a614f5e0c72dff06a0c1d836c7fe4a2c4086129386b34dde) +
                      (Ic754ed4f2d29b948b422876f371df4f89b86976e25183ce1b9f664e1a9b19f56) +
                      (Id7310932ca8964fd49adc052220c04855b028e29fb7a48521a36e2dbe1d6d5f4) +
                      (Ibae8222f76059e8f61dff938a64e23080eb668880ac50ecbb50de852472a22ad) +
                      (I09673e64aaf6f35dbf4aae16ffba969d08a800d32ab25413bfcdbd540d7b01f3) +
                      (I3ae1a42457a669272eeff1bc293c80c67239ef6b725a09eacb82b06ec84edd65) +
                      (I5b4c4554a78c551dd34a93ceb225237a2d2540a0e05311c4595bdaa5a4cb14ea) +
                      (If27288056468d3ef3052303952f2e4be67796c40d6224383047d71d996f98cf3) +
                      (I12dfae8d4c1a0612c6d65c6f5493247af5e06ca1d8c72dc28f9ca41b0bbc6ea3) +
                      (I295da244d8dab1563a5947230e49171eb905c3758c289526ff6d3e0c3efcebbb) +
                      (I89cf2ce418b6d96c0e2b9c8e82167a47d40ade45a8f08255a1b849a9df9e6d06) +
                      (I47ba4d6ad7b1889cb52ff7a1d42176e166270e39a1d2875f3a0cd260a1fc92ab) +
                      (({q0_1[52],q0_0[52]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[52],q0_0[52]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54  <=
                      (I08240dfbc0f698324c1ffdb8e769016bb8b947fb0b8dbb72839375cdb4cc47e1) +
                      (Ia9ea47bb0829c979af002fb7aa0e22072671c2876bcdf79365ff2b3691172149) +
                      (I58df4f7ee4282cdb7bb80c9f1d907ff37590b1db22994f3a07b521132ab80087) +
                      (Iadfdcb3c0764107a2b0deaaf039babe6a08f1018f3718f5539718ed6a5aa962d) +
                      (Ia2417744c8f15898d5d951e15cdf8c03d932cdac6acd27e32045e0fbfbfe4f30) +
                      (I6d70d8c6d44eb58daff53226cbb59eb647b6dec6bed37021a64e16ac5318d484) +
                      (Ice3b06f04279add8283c8173340c2bfd4b4801d85610179943f070aef508a893) +
                      (I4fa5ada2d589c7a90e700745aba8e09edcfb0252f532e4c74eb0809c712a36f0) +
                      (I71c6f88cbabd48d41f42f2b16170c8955b79d20b8a8b211e174d1c1473567ad4) +
                      (I1e7e130607ec849c80f9e687f0215ceb767a2650626f20ee44a6fe677fde2299) +
                      (I4c02563233638e273f05bac3e277c702b38c204fda200dc5ac163662c77a429b) +
                      (I85d8f259f770b22a380d6eb5ace0281c57f0952506152be05f38482c47334988) +
                      (({q0_1[53],q0_0[53]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[53],q0_0[53]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99  <=
                      (I989259874d3f12b373358db47fed6245f192edac9e7df00531ea7ba75c360d4c) +
                      (I2ef69d9eec4f925b598115d569d2d85a4545871f2ac62635f9b072ba718b595f) +
                      (If8cefdab8d831c3db83e1ef615ca534f34c58b9903520c7741cafbc84e28d207) +
                      (I00e5abb30adb527f6b32257212dc21f9797e9793ebbcc10feae9e524188539d2) +
                      (I9349cba960e03e6068aa27e997993b0c466e040a1ee9e6053536d3346c84214f) +
                      (I19797110801d39a7970e6d8665215c967071ad9a1bad12c33401b44f595772b7) +
                      (I0d25b3618b50ff21e3f301fe44087368e38fd6b37b6f6fab004824aa9df51f0b) +
                      (Iba62c53d136b455b7d575b868f2ebd2dadc6003981aa2aae72863a0eb812bd1a) +
                      (Ia6f2e4979fa9229a647a81a4fa3f8b2af809199049d2554ea15fa9a6ba2f90a9) +
                      (I83d70d4886f48dce0888e203c2c333c76d35f0c73767dd9443ec8fa4790ecb09) +
                      (I3f92074e96f2c2711248b1d770b4ad718a565a323e6fe4ebb379e6494039af47) +
                      (Ia478acf4034b69d392277c3d5c6683346547ff26d418b3a6c36a3f9a56e3cfe0) +
                      (({q0_1[54],q0_0[54]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[54],q0_0[54]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec  <=
                      (I06186aec49594899011a9d7bce163a3a43ec094d7c92033df033594ed5eb43ac) +
                      (Icd8ef17fc44642a3c86a1cb62727eb607e3a4e6d0b021406b9b710ea5c96c06f) +
                      (I2a3d1a32b282fd624497621815c6ff85c904f5f3fb50f18cf345c5a5d7a557ef) +
                      (Ibb57ab5a5468d08c8b299ee67b535b83995e94d6223d0c6d93dba8580906e319) +
                      (I6fdc128e94d85f0f7f884ee1ff44fdb6de2ad5b93d83c3e36ae235afcd3d23c0) +
                      (I2790277776fa84c3edba2332cf538f8ea3a40c1b06cece7463a3b4757b1fe213) +
                      (I068f00aade8307d2a2e2ddb37d7429a04c2f6786232134a041e62733cadb03ac) +
                      (I07087056bd31363bfb1f76f8fbeb18d1deafd5e4816ca1200d362c0797a77bb4) +
                      (I01c264f9a89aec9dc11fa16206ffee1c8fb03bcb279e9e9f53fea1e94e9d8b23) +
                      (Ie42f89c20abd223240a9f93a89ce650ed2f581e1ceab0587a4fea2ddf9f4f98f) +
                      (I44ba42cf2460fce5fde6d8a9fba799517336268d29b5817597d819a9eb83df0e) +
                      (Ie4fafd34aeca2efbfd3bfd3bf45f73ceea27b613ed242a43666d85f3680ada44) +
                      (({q0_1[55],q0_0[55]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[55],q0_0[55]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7689b1f287170d28fc72712f5ff2fd209108b000a63e268b12da08dfed6d60b0  <=
                      (I65cb4f1288affe61a7cd9981878d8519db25d724cecbb80eb3932ccedafcd5bb) +
                      (({q0_1[56],q0_0[56]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[56],q0_0[56]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic114200c11d550dcee2bd668ffd91dbdd193a00571dda2d6f99b4985ef999f83  <=
                      (I577e642ba232b9a606abfddc4d84ce4354744e2f953da3b285e417dbfc5aef16) +
                      (({q0_1[57],q0_0[57]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[57],q0_0[57]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2090cbe74e266e4385d5075f2913013cc38b26c5332d982cabead5dbe52d7775  <=
                      (Ic68515eee7d422be9cf8950e48b81d743d5491851d5a117d1f9b70d1d9b55060) +
                      (({q0_1[58],q0_0[58]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[58],q0_0[58]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7802f219761d40fb4b24650bdbbc6faea69cf01618fbddae575028e96aa7c627  <=
                      (I0ca47358f982879bb85bd78f6bc19192a5ed8c62214073342b37b040aea331b2) +
                      (({q0_1[59],q0_0[59]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[59],q0_0[59]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I9e11bb32c337ed1d87274c3040deee6d8813fd3f6795de87aeab9f93686ee409  <=
                      (I1606027ef88387f2150285b55cef89212359f49ab1a49fb71e457a3dba0c438a) +
                      (({q0_1[60],q0_0[60]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[60],q0_0[60]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I08382faacfb31fa012c97cbde6527792abbdf2c9124d886540d385dbf39e24a7  <=
                      (Ic09f51154140ef91861243d7b35f05961565b368264d44c8fd5d0f85bd0fa213) +
                      (({q0_1[61],q0_0[61]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[61],q0_0[61]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5c8ffe997fea9d77126fb36c6deb4f9b9c9b38e6aa562b574011ee5915a00857  <=
                      (Ie28425115106f4b2405fad6fb2994a76e64dfa60e7bc165f46ae67411932a1cf) +
                      (({q0_1[62],q0_0[62]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[62],q0_0[62]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6f9b56f1fa7e83cc6acf75b74037938bcd08ba89ac2cb3dbf4df512fc9d521f8  <=
                      (I64862889bfd7d2a15503bc07af594be59cbaa8758863f78311d6f15ecadcc99f) +
                      (({q0_1[63],q0_0[63]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[63],q0_0[63]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3ea241ea179029fe0c486fead3909ff2c05b2d47e4484549d1d521a4f891a9a8  <=
                      (Ied4424f3e85f3fb92f4e40bc63909f4e77698a18a1d0ee651e54e4de06ee330f) +
                      (({q0_1[64],q0_0[64]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[64],q0_0[64]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6f9fd1c4756d8d1250b0ed96355e2739d3bcdaa3603b7e1cb5cb0dd0ad5985e5  <=
                      (I6c850d46af2f31f4e3d31c3fd2b2d9c7471ccf817b452a4fa2602485f5e7f164) +
                      (({q0_1[65],q0_0[65]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[65],q0_0[65]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If084c3e6863c87018f76e95d715c83cc83dd85ddf7664f98c6ff35e8a0ea40d9  <=
                      (I1a1a9f7ee74e17c4a0d7064ca9fae938002b1b685f3cb6309569081b0d971aed) +
                      (({q0_1[66],q0_0[66]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[66],q0_0[66]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7fcd9ade547e48c042200e4bae7d4699b326df8a285204b7e23eee2a019cb01d  <=
                      (Ib5929b32be13a8436b74dadded1f26d3742e1424b6025d1eacda112bf4749a15) +
                      (({q0_1[67],q0_0[67]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[67],q0_0[67]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I9207b21b45d4265cc52ef02ed257ea78cc5a269d98165b2a7714a25b1c477521  <=
                      (Ibcb7809e1db6cb82ba62be017c5b8685cb6f988f85a0d29ce2459f6ac80498dd) +
                      (({q0_1[68],q0_0[68]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[68],q0_0[68]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I4322d4cf469c3caa560e48f6eb1fea264c42dd76b65977c24c676681518691f8  <=
                      (Idb971d0017094cf8b28e639623f85e6e5fc2c03a1da1e19a1ef87b959fe8e1cf) +
                      (({q0_1[69],q0_0[69]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[69],q0_0[69]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I924625bbe810db6c8d5cca4407571d5819d0f7361e2d7f1906bbeb822457aae4  <=
                      (I89373d12365deb440d5337a2586fcdab81347ca28ff6f261a12e35a235bd23c6) +
                      (({q0_1[70],q0_0[70]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[70],q0_0[70]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3a01e4ea96fcd387a6bda68d7d07cd6b4e89ca653c798f08ac8402696b42a371  <=
                      (Ib8f9b76d6cf7a74f0d437f634ce888096a0d6d81d66dc6c60b62a60006b661e9) +
                      (({q0_1[71],q0_0[71]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[71],q0_0[71]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I96114d8145aafde7f8f5666ca2f6dcea9ddfe9796f2e3a54556fb1b23fb1a331  <=
                      (Ie55394a5e3d49de60fbc4f33b3f9813b885da2049376036c935e8cd7c85010d7) +
                      (({q0_1[72],q0_0[72]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[72],q0_0[72]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I006672e4b2c9c693fe5b05655ebb6f31e96ca8e2c92eb488cd28e5a940e49766  <=
                      (Ia6240db37d8e82731a264e5e3eeabb88e632dc6445647a26b4abdb142ff44c03) +
                      (({q0_1[73],q0_0[73]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[73],q0_0[73]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I408f22a4a77906024a2e6ceb970b39ba9ca76300fb2584bff35e37da452c6613  <=
                      (I4dfaddc409bf6d3698f255e55590182c2c8c067e0766311322460720dbd0967d) +
                      (({q0_1[74],q0_0[74]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[74],q0_0[74]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie84e7eb709edc06e55ae27284cb93a0c656ce8559679c49a47c7f03f0d64fce2  <=
                      (I1dd3e1e1e78d9e24a54fc937e7a25fc0e2514eabd1c1cc662d81ba73aa44680b) +
                      (({q0_1[75],q0_0[75]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[75],q0_0[75]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I84fb24aeaf533382e57c00dd73683ce0e4f5f33a0e7a3b36f2ab00732891682f  <=
                      (I80d4a0cc8b63f2ce0dcb344da5a47c95cc28b5f93d5bc6b77e9b875cdd58db99) +
                      (({q0_1[76],q0_0[76]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[76],q0_0[76]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ifc8b49d8467101e2eedcab4b6ad6a73e4f657c0e995ccaee5dee276a5ae916b2  <=
                      (Iec19b0b63d20ea69dbcb23411a298bb6e833ee523fdf082f9343a695891a990f) +
                      (({q0_1[77],q0_0[77]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[77],q0_0[77]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I001fd8ecbe068f57df7498db3f519cbb5a65bc5af187f1d34b5eab3df45447d9  <=
                      (Ib612f39370c6527c5f6eedb0eb5e7676212642673e940402586e823ddcbfb4c6) +
                      (({q0_1[78],q0_0[78]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[78],q0_0[78]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I11745815606a2dcec9059a24625e93a31b0f15d9b81c97403905e00d3fd64f43  <=
                      (Ifa501efa24e47050960fb3c383458a20f54abcbc5ca45bbe2d15a037670cd5cd) +
                      (({q0_1[79],q0_0[79]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[79],q0_0[79]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I37a341bca6a12362e49dae8435798cd8e7550a16cd506a7f852f4223088bdb4d  <=
                      (I8f088dd043a22011add21694f90df62fe1d2f6670cc72cfee805c9fb49756c77) +
                      (({q0_1[80],q0_0[80]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[80],q0_0[80]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I8ab2f0a2c9cf1f1e0401a67f3749b106fac7d45293bb9648325f330e3230517e  <=
                      (Id86d515c6d081de87b9ed3c3521ab079e93ee082d8a0b396d44b3b70cac06b9b) +
                      (({q0_1[81],q0_0[81]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[81],q0_0[81]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic6ce7ef3f9390c17ef23e718bce985f168504ddff0d66e2babddf08b37dd2819  <=
                      (I4f94812066080b656de1a2807f5f669b2a81085bfc0470f9868bf5945856b451) +
                      (({q0_1[82],q0_0[82]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[82],q0_0[82]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I26c16ba52eb0f661ca599263265d1d0d7e1f155b4afec85407f3ece6fff3c391  <=
                      (Ia92baf4463c96e210b460ea02d7775353edc6d475d7a315b594b9798cfd17900) +
                      (({q0_1[83],q0_0[83]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[83],q0_0[83]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I31afedbc324d4ddcd04b3ef766154a6414cc6e31eedb0ff24b40698430e84927  <=
                      (I9d4c230c86454c5c5f9ec98917ffc8d23fd19105ef93ba860ac2650bcf43ba4d) +
                      (({q0_1[84],q0_0[84]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[84],q0_0[84]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I807fdac75cca555b8d81d1b4d7e53ae7cfa0e4b83bcb260cadae218faed4f781  <=
                      (Ia4a28d520896fadbeabee4130dcf862a9542852d87be480b1df2b67817f0ce65) +
                      (({q0_1[85],q0_0[85]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[85],q0_0[85]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I0f8a9c8deb02bf990a6ac2ac0569f9d0ad9f167d7c18dc70ba544912aed4bf78  <=
                      (Ide9498000905141bb106efc7e2184bd460d0e59a2270b10d42f981cf3bd514cb) +
                      (({q0_1[86],q0_0[86]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[86],q0_0[86]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib3e6663aab02fdb649843c552944b6e325240f5010acb414c311ae56e78f8459  <=
                      (Ie9a6b0e499ede3f80403e8f9c795ef4e93108ee8db755e12fb931259f1699712) +
                      (({q0_1[87],q0_0[87]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[87],q0_0[87]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I41339bac55a76a05186d632423b1fef8173940f0cbddfb64c83282af5cd04cf6  <=
                      (I362132341c8e8a464a2bc93e7cc5b1d9d7804dd93965614dc340b48fad5c92da) +
                      (({q0_1[88],q0_0[88]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[88],q0_0[88]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I28fb4df9f762474ad496e8689f21d13bcc5bd4fd79190892b78409a06720e2f3  <=
                      (I4b3c222863418745872c878545e419ee8f9c531f2cba89d28f0787992b0be8ed) +
                      (({q0_1[89],q0_0[89]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[89],q0_0[89]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I84ce9c6711b257cb8cf2f09bcc02e0f03490605e543ba12942207df6fabed5ac  <=
                      (Ie39e570f1b5dd9f1ae893af78d81e458d077fcde2aeaba432209269b79785582) +
                      (({q0_1[90],q0_0[90]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[90],q0_0[90]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I8f3d31b6843ca54e80e8f61be651cb7788b43302b001d791357fad349785eb1d  <=
                      (I50ebc7f8f7cf324814b5885b2b18c90bf5007d8030744263d6e66880d836eea0) +
                      (({q0_1[91],q0_0[91]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[91],q0_0[91]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6fb6112b591f6f1495935e422361833f041f7231996d88a3936b5da186e4c48d  <=
                      (I326b57b49d3fcfe654c4cb9ebcd6edc0ad7969e3b531f498e3c31270a5c4aa70) +
                      (({q0_1[92],q0_0[92]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[92],q0_0[92]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I959de6064e6c31bf0d18c2d6b4c274ebd5e9fadd996fcb32e695047831716951  <=
                      (Id3898be2185f86831f58bd16651edee3d1bb21fa07b33a1928740ab496404178) +
                      (({q0_1[93],q0_0[93]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[93],q0_0[93]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I0f46fb1c05f0f882ae878e86285077da38a459201c305e13fb4925ba34eaef8e  <=
                      (I2aa77512781cba636ab96a5d09527e1ac34623ea2bb6c6a8d742bbcf6eff499a) +
                      (({q0_1[94],q0_0[94]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[94],q0_0[94]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I99e249a8eaee9127d347ab629dc27a21d5b55d2826c354eaffd9e6fec47b1043  <=
                      (I225543794992ac9aa68ac3eeea38d41077ab5512b9f3b95fbd65a839294088e9) +
                      (({q0_1[95],q0_0[95]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[95],q0_0[95]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2f779bcb2996facec77594ce5efd7c78acaa443f2b6ab3a5506ae96dcb986b23  <=
                      (Idd1dac44a6f35d558d400160a087fe7628ef80ad72c3962df2b3a3809b89bcdd) +
                      (({q0_1[96],q0_0[96]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[96],q0_0[96]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ia765277dd8a5fbb2a65aedce2934fd6c4dc9daa4e0b316604f6f137f19fd5d25  <=
                      (Ic039114ea8ac4120b09973c79fdc044251fc66bdeb18a498dd6ed7265cdfba2a) +
                      (({q0_1[97],q0_0[97]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[97],q0_0[97]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I1a47d1294e98ebbb0493fe3cf7743d1932eac70fe9d2754367a51d9a49448d12  <=
                      (I21b3fa431ddc4bc8eacfb17a90fdac2bb32e4d0f4d0118715642c37601a1f883) +
                      (({q0_1[98],q0_0[98]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[98],q0_0[98]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I71c11e07942c42d17f5b85b1da8857e91f789966944c1e0948bf5f0285c91079  <=
                      (I1c6d953c9a0e96d328cc4b515867b2ac21d2947a85e96be19f38e67a8b15001c) +
                      (({q0_1[99],q0_0[99]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[99],q0_0[99]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id810b154e951f2b2d0b8ae826f31effa4f39b3a0396d446ebcceedd7225c5018  <=
                      (Ib823a58e9d4db87e4d73a81a772a02435af32a11d3c2265fb8a16021cfe4503d) +
                      (({q0_1[100],q0_0[100]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[100],q0_0[100]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2a96d9fee197ec3bcdd50abe43ee0d3992f5b03db5cdc958771ed812bf3a0b4e  <=
                      (I3427390162b0952481e5f0728a20075c9cfb814431ecbb1a4014d407ab3b3afd) +
                      (({q0_1[101],q0_0[101]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[101],q0_0[101]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I280a4a7c5231cbfe245c071a856f7d1560c4154e9f9a4c5fb6895baa2f4f5871  <=
                      (I35a9ae1cf23d8697091de65a1d0678632bd6889ae32408d7658e542a756e95ca) +
                      (({q0_1[102],q0_0[102]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[102],q0_0[102]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I01562027a6c7a542ae356bb1d0db0dc55b2094f3470a1894e67a3b7fee9e4361  <=
                      (I37e54e8ae28cf1a36cb9101d5afd4d523ca9a6ae244efe641c547a4114726bea) +
                      (({q0_1[103],q0_0[103]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[103],q0_0[103]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie3eb1aebcdf48fc8f41590f0e9524e989193fd14fae379a200c20d1fd3755db3  <=
                      (I9544a194d3d75c6c414169ea2536e111c09711ee602eb3462c4022350906a21e) +
                      (({q0_1[104],q0_0[104]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[104],q0_0[104]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic585c7a7014e8bff08f28b2d432e9783bea57ff5b456d851503a2c3eee80a768  <=
                      (I1e4bc72a55efb8462410905dcb2c9a8412e2533ded854d23ca648e0e36802960) +
                      (({q0_1[105],q0_0[105]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[105],q0_0[105]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I4f0a460fa116f5a45cd0c435e594ccc7597b449cf5205391a2dc6e977f4bdeb1  <=
                      (If2cec64e868d25d7fbad45ce4889c6a4cac0084aae00d2aa8963678edbb88875) +
                      (({q0_1[106],q0_0[106]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[106],q0_0[106]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib7f3bef766d8e66cc9002dbcf3538dbe974b70de4d7a8a3d9cc3bfbe815841d5  <=
                      (I73ad61911b0822e313aab2c484d1699cf2655a42a2bb0a1c9ab36228e41d0f7f) +
                      (({q0_1[107],q0_0[107]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[107],q0_0[107]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I027d6136f1b64e5e2f94af338f8fbc0ef9fdf8dd0a2d58aa0eb6879557361681  <=
                      (I218255d96e659dc8f60cddd40cac94a56d93556ed609b60157d88b298ec95f0c) +
                      (({q0_1[108],q0_0[108]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[108],q0_0[108]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic62f1d181b6452f30ab2146b4e43113b2ca1bf21962f686be46f59084d39fa0e  <=
                      (I11284a18d6115421b4c76054c1a580c41987dec66caa7d5bd9107bbd4ac8bc2c) +
                      (({q0_1[109],q0_0[109]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[109],q0_0[109]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iecddbb8ccabf830117fa8836a6eafc8dda6fa463d9c907ea25d298249bd066dc  <=
                      (I8516ef195e4ba8f6e29a02ab5ea349a26bb68f6ebb4da847d56c03c942e9c20c) +
                      (({q0_1[110],q0_0[110]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[110],q0_0[110]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5a2b6e5bff0ffadb36a7f02dbb3cf48ffd37e6e29ef09200db12ccf9fa9d8450  <=
                      (I2411dfbbf605c7590bc678373dd20b7241356a433756332f9a3445ba8dad57fb) +
                      (({q0_1[111],q0_0[111]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[111],q0_0[111]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3a9d955359963dadbc16853d82bc2495f84c37d8cabb868a144c5f24d9edb2c9  <=
                      (I69d896cdb2303b99b73c4d6886f2686381230feca86c62fc064a85e4d11266f4) +
                      (({q0_1[112],q0_0[112]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[112],q0_0[112]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Idaf457dba6ceb8f056ac34d3bd84bb9e9554c0d55db8928b9b48692c316e6fc5  <=
                      (If6ca882e537cdf5f458a2e11b7a11f057a3d2a00923825fe236afa0b0e1442c0) +
                      (({q0_1[113],q0_0[113]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[113],q0_0[113]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iec8531839aeb35f1c356e474abfc871d1ce889c4aaee1b37b272dd9650fb6981  <=
                      (Ie35443efbbf821e07284652a4b37347c4cfb959495dafa4fd2f81ffa2edc56db) +
                      (({q0_1[114],q0_0[114]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[114],q0_0[114]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6a320bd601e721d94d7ac0aeb59e2c81a0a9737d2f7b49d668369336dec2ebfe  <=
                      (Id6d0b1fe00e5324e0ed7c37d41ee3e848f9c7dcfb4a85f5da2b82ed4d8942b21) +
                      (({q0_1[115],q0_0[115]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[115],q0_0[115]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Icd9be4d5172c268eba385d2cf858caf3450d81a87bb90fde24fccae0d1637d99  <=
                      (I0a309e8aa7f7e07abd837c99be6d8bb8c29dc1679b449111a02f49442d5cb432) +
                      (({q0_1[116],q0_0[116]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[116],q0_0[116]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I64227cc72d5c6450ebded626fdcdfd149c8e29dcd6839ad76b2b9a932817fdf0  <=
                      (I416c7ff28cd1d182ba2e08c3882c04d5073a014f7b9b41e56a3850cdc289ffb4) +
                      (({q0_1[117],q0_0[117]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[117],q0_0[117]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic754b281b704937ea08e702dcb74b7175f8901b29809052424f867a6685c1d41  <=
                      (Ie44d1a587dcdbb709546c6c567988fb0a19c276a1df7aced4c09a029196dfd4b) +
                      (({q0_1[118],q0_0[118]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[118],q0_0[118]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I861b39dacbc8ae1c9cb21a407a53608f0d5adf148148ddb8c3ab1cbce25e2497  <=
                      (Ic2b8d811fd01f5cd88dd60bb1b89b33163b3cbeae48d04e2316f15500c6a1a40) +
                      (({q0_1[119],q0_0[119]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[119],q0_0[119]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I994137ceebfa9f1bfb6f3342c02ef25b1a5e881f6fcf6c2e7f274663b5b4a3ba  <=
                      (I85ff9ab4f9a4a3301bb8fcdc7107202263af0c37f091445efb5fa163a6b47a51) +
                      (({q0_1[120],q0_0[120]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[120],q0_0[120]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5193db4e129f33dd7cd8691b74f52f030a066b583bbe2d9a4a6e9962f1c43280  <=
                      (I39ab1bf4bdde9805c5bc7695c4700975d5a6094c40e107b82477192005d9ce21) +
                      (({q0_1[121],q0_0[121]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[121],q0_0[121]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iecd0fbf7643812e36e8d17ed6782ecf4b181df9d284988b1f416de07cdfe6095  <=
                      (I602591ae56f1a42c64e50378841e065e79aee138622a0a571effe20cb48645a3) +
                      (({q0_1[122],q0_0[122]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[122],q0_0[122]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I390b2f0e16e0de51443f9cbf8ae301009d17581f5e20ec4956a8e95ede2c0822  <=
                      (If37e9ed3af8a31c989dc6ad554207cd464c591b630ca1e5cf56b2eca57a18d8c) +
                      (({q0_1[123],q0_0[123]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[123],q0_0[123]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ia733b3c17807a98828719894627b0a1fb161ffee86fb28c11d92f5b185a6284e  <=
                      (I80099c7b01770cc5f7edb3a3551d8edfe9dccbcd2a12daf8ebbafdfccd141bd4) +
                      (({q0_1[124],q0_0[124]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[124],q0_0[124]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6b87b44befe3363656697619cf3dd967526646ced0f90813c24c960ad4d57d5f  <=
                      (Ie479ccbabaa8a00009152557e4de08bd240fd28f1b131c674dafbcc2505711f7) +
                      (({q0_1[125],q0_0[125]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[125],q0_0[125]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I29ee4a3cefb214cdfe60e6907e63799323eec92930d4a48797c96a7c1f3e3a15  <=
                      (I6364406b04427fe3a4cecbed48e12a67cb08dc632b2914b0fe52fab0ca541c0d) +
                      (({q0_1[126],q0_0[126]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[126],q0_0[126]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I748cf7beef2ac47341c77503d0042b6e1570248031f1d9880d0bf14969378379  <=
                      (I610dd39f1d44d84764b0acd6b3fb1219fb6b6d6ca92e1b226ca76a389bf6c937) +
                      (({q0_1[127],q0_0[127]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[127],q0_0[127]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I559b90a32f7cfdeb35bcf30683787c6357460614330553ffd4f5732cc03507ed  <=
                      (Ib9f9384ac4ec4bad29fbb4ce683ffda7dcab311135f02b6336e6209f5742fddd) +
                      (({q0_1[128],q0_0[128]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[128],q0_0[128]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie6d770decdaac3d75cd6c9eba7edc89898bd152a7c75f43a464a47c9994c9a87  <=
                      (I60980f76d468775bcc8a7052681fbb6ef4b2243e5e30e5365cda6cf598bd0bde) +
                      (({q0_1[129],q0_0[129]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[129],q0_0[129]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6541e01880f3c658b3404a81e96fd03b861ba4a26ec927e9c2c64aa9973dafc2  <=
                      (I892a754f0322d92126d4731e8066760a24897f93e2afb858ee1393604d2cbb26) +
                      (({q0_1[130],q0_0[130]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[130],q0_0[130]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I184fea1e133f0a5b9b8a88926ebceffbb79cf7816941eaf9a326764d876c924f  <=
                      (Ib0f8816eafd3b950f67cfbdb6a44c59ab7c0918979817a4a998d8305da847e72) +
                      (({q0_1[131],q0_0[131]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[131],q0_0[131]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I78d3ad872172f1089358c601e00c98f526455a961f30bfd6a966e8d8bb6bd098  <=
                      (I04b55f2c45002f1f1f7a6176773a22730dcfea14662f0badb102ddb60b84cf9d) +
                      (({q0_1[132],q0_0[132]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[132],q0_0[132]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ibe18bd1138dcd8295a35b807d811d5b05b07df9efd2326d0cae0cac6589e7bbb  <=
                      (I5edc072d158ac583bd1cdb2449086d4f0b17e36d724f4cfde79820788ce57f31) +
                      (({q0_1[133],q0_0[133]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[133],q0_0[133]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I68fb3ebbcbcaf18cb81eeae19529cbcf7fe4175df44bd847d87ba9675ffa862c  <=
                      (Ieb128919ed64e331affb6adba798c267e8c3ec924a7ef58f50b1bc0b29702c23) +
                      (({q0_1[134],q0_0[134]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[134],q0_0[134]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id2154e04af88ba8cccdbe100e1c4e4bccbffee35bebd3d43f9229d2915bc1deb  <=
                      (I90cc372cc2f3b23eaaf2cb32da95ee715af64ca2eaee77195d9813647d2a0d08) +
                      (({q0_1[135],q0_0[135]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[135],q0_0[135]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic95be152c428a61c5e57fa5a5e776b9341efe9f2d08c73fe0a9d2663b0a974e0  <=
                      (Idaf65411d995039ea730b6ee4b5ae727325da17dc79c8664270d60f063828453) +
                      (({q0_1[136],q0_0[136]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[136],q0_0[136]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6e7d06d6c6a765e6994847af070c889f9c7059754ed634122e0204f750919234  <=
                      (I977557441002c273f9b9b8748ffa9edceadb342e028ceb581c3bbce9af103a74) +
                      (({q0_1[137],q0_0[137]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[137],q0_0[137]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If0343bdeee565245554859329a0188f1267cab02c325fbe93d4df18606760025  <=
                      (Icc10ac19a64065f5923ecef4f1353f13c7796c23f2555f8ae6566eb538d77677) +
                      (({q0_1[138],q0_0[138]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[138],q0_0[138]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie090cc0a910baacb33f7e858eddac0b221b9a5c567ebde9bba44380b06e8dc29  <=
                      (I725c369a5013eeb6b581209bc8a921fccfcf1754137191e26757abdb72ced94b) +
                      (({q0_1[139],q0_0[139]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[139],q0_0[139]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ia0e41f1ae6bbe04c95f97b4d03e31d86b4399463bbd9fb5bd714b9c2b58bb23f  <=
                      (Iaa02b7ddfffcecb763aa916a2bc4c3aea58027c89b515c40b72214d9dd44ba21) +
                      (({q0_1[140],q0_0[140]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[140],q0_0[140]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               If4a86cc5d7bf6b2552861b330822e6bf86fa60debb5d503d86e081b720f3432e  <=
                      (If8737fa82b71d9b0e7223baabca7405e148621600bdaef02e65cd7bd175b2d88) +
                      (({q0_1[141],q0_0[141]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[141],q0_0[141]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I0d2ad8151436f1c3336aae018a92e8bd400452c12972fef401e7ab55030d285b  <=
                      (Id85c2b905d61bcdc87d500d6ede3ca02d52bc3eaf278f087f27fe6f277c91262) +
                      (({q0_1[142],q0_0[142]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[142],q0_0[142]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id2881f7fc5d7a68a4583d24b1a8a9e09928ea1e5e3ec22fff19d4d59e12a201e  <=
                      (I5923f41aa444bebfc18d13202747ff84e20a4753bc9cedf697b9ae8ec3418afa) +
                      (({q0_1[143],q0_0[143]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[143],q0_0[143]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I8733749031c60ed31e2867dedeae4f9ddd4da169ff086c567288ece5da43decd  <=
                      (I4ac498dc826a9dbeaddf2f013ae7116e92dc772ea55987a4661f18e56a4123a8) +
                      (({q0_1[144],q0_0[144]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[144],q0_0[144]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I9180b03e001160fe9a51818e7641c427a35e0b2cbeda9e6bc0e32878bca05815  <=
                      (Iaadbb1b235a85c555a6f37d003e87a987b7d9b07148207555eb717b7332f67ec) +
                      (({q0_1[145],q0_0[145]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[145],q0_0[145]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2f00eb344711414f5f6efe7eee64b5690b4610385673a7186711075eeb319cf9  <=
                      (I6afb533ec993de4f9b04007b355a9cadf08488ee6ca02aec2d7916a4c98a7fad) +
                      (({q0_1[146],q0_0[146]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[146],q0_0[146]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iea8f3fa357088442ab8048febba14f1e6ae367c6b1a854ce0b2c4861c4a2ed27  <=
                      (I01313177417c899543a67763ede925dea3ee58ef4a31714ad15a7a3746bb5be5) +
                      (({q0_1[147],q0_0[147]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[147],q0_0[147]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I0d3923859952e0ab6d926924645383b83904ee287f1783cdaa7f314b171f4171  <=
                      (Ibd0ba147d1a08acea707b8c60da14ebcc4ad62e67ef26634777b5dae38af6d61) +
                      (({q0_1[148],q0_0[148]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[148],q0_0[148]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I45f444d890e00116a19e16e3c50c555419e910e2413c0277f62032d6ff66ca15  <=
                      (I1e92e18a915678cc96aa493a00627dffecbd341dc8e022615610061e52c1ac3f) +
                      (({q0_1[149],q0_0[149]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[149],q0_0[149]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic67dc4f0898ca883d489eab901e11caae2adbe1c1c502ab57f5366cc26d4d335  <=
                      (Ia7b91fa4a1ef16f859ee162b91daedc97927244dc19aaedede898049daf85a19) +
                      (({q0_1[150],q0_0[150]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[150],q0_0[150]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I89150482cc550af995633308cb14fc4aac6984b8c5bb09ed4018e5692f8866e4  <=
                      (I9918d91748722a47f8526008bc3fd4c498bc80205211d5c92acbc511fdb667bf) +
                      (({q0_1[151],q0_0[151]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[151],q0_0[151]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id4c7f10c8e46d38df8e36571905e342a0b283e8badd00d3e4081890010c25f34  <=
                      (I95d109e37a87827de1455b5ec479dda78a0218cb9db245b80710cdb1e8ead67a) +
                      (({q0_1[152],q0_0[152]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[152],q0_0[152]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3c6ebb6c57609827961bfb1e39059b0805cec40a48787adfc9b2b138a5012c9b  <=
                      (Ia0c7162290e415f24699688e45850c243397b5cccf07daf0398dda04810b0690) +
                      (({q0_1[153],q0_0[153]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[153],q0_0[153]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic8177ee86d033bd8ab95b63937a4f80b02ebbb66d4c16d84c8822d133e7cdd0d  <=
                      (Ib9dc17b2b9fc7c228eba40cf625a49a27ec16f8c8a91957de14fb6849ea49212) +
                      (({q0_1[154],q0_0[154]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[154],q0_0[154]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I65cdf21d7c52f9a1fd2d4bb265a678e8b543e0dedd9fdc5cf9e12ecf756e66ae  <=
                      (Ied32ced79448b3f92faf0dca1673559e07372ec338e8c51a750be1c6975a298e) +
                      (({q0_1[155],q0_0[155]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[155],q0_0[155]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib047d12eab2012f21895617ed9bff57a0678c2c85235301fa1276f99ecc8625f  <=
                      (Iaddb000276bde734c13ec1395f06c1b3bf5606ad5cb138579d711cecf26ac88a) +
                      (({q0_1[156],q0_0[156]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[156],q0_0[156]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I4864402239c958072b187da428e64688ab13cd5a3ba940785ac5086f81c50e92  <=
                      (I211ada7f9095ced6b3d20f8f7f67b56cd2e73595481ed5d4c08175ca874d16ae) +
                      (({q0_1[157],q0_0[157]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[157],q0_0[157]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I8d03bb3beaf84d3f94a15648cd5536d5f14020daffea4160bbd12426018140e3  <=
                      (I0d49182fe7486bcf54c8f68904b4b90436de6f3bc42fab67a4e47f61154e22c4) +
                      (({q0_1[158],q0_0[158]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[158],q0_0[158]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id3b64ab87f29683b9210364e13398a54c486d0b8b8a7a5ec6f15c29cf752b5cf  <=
                      (If79b91295d25c503f6bf5ca7c6eebd2ebf6807dd9990ce31e844cee0d8f89dac) +
                      (({q0_1[159],q0_0[159]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[159],q0_0[159]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2f3b819fb1f865426e38d2b39a1a4a8ea0560e0888f19913e2393d416205f3b3  <=
                      (Iec1d04d20ec09595743b7a35860b5cb2ec862c20da87c6f899284069c60bdd71) +
                      (({q0_1[160],q0_0[160]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[160],q0_0[160]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I23e7ddde350dba3f41b08c523c29dae580b57e09b8fd9d35af6ba3bd4b104b6e  <=
                      (I2126b1597a95d7aeb7d20d4e0f4270e1fc5cb0fe6eb5003b05abbb7e5e9a2819) +
                      (({q0_1[161],q0_0[161]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[161],q0_0[161]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ifbd6430f8434621a650f4942f3be3669bfaa802cd912188e4139542d2a64a511  <=
                      (I72a115d9b3659f31366e1d73d6d9a0793e20be233c3ccab2b513fd79786224bb) +
                      (({q0_1[162],q0_0[162]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[162],q0_0[162]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I1cb9b876fadc25322c3f466b101084a68e5a283260303beb238d55ca788523c7  <=
                      (I469b0bcfe9cfc27a8596782bab479f30aedaa132a5cd404feb1fec4b52a17d3a) +
                      (({q0_1[163],q0_0[163]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[163],q0_0[163]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I9bd2fc6de34fc3d410b3d5e30c2e9e811c7063afaa6888afd119cdc02e39afae  <=
                      (Ib4c52550766a2cbe0de236d6783edfb1a6a7cb4c2bb9333a9379e1b75680dad1) +
                      (({q0_1[164],q0_0[164]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[164],q0_0[164]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I9e9c82e0f8d919f8e2e03046a1654698592da05002140ff69fdd551598618d59  <=
                      (Iaa72101e8c3e7fa248ac4d4336b3847c4f602b6db009e9cd74cdd25251d5178e) +
                      (({q0_1[165],q0_0[165]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[165],q0_0[165]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic9fded9a702f4299431ec45bc00c9111907d62279133f1a5f62e5f6527823aaf  <=
                      (Ic1381219782d18c1cb880970c062eb260d9d3be0b597e1465fc604c0c0c32c68) +
                      (({q0_1[166],q0_0[166]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[166],q0_0[166]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib95adef89f659c6d98e43f4a9c43340a0acdf273ea6bfea0b8e99f0751c250e2  <=
                      (Icf0c3c82c9e458a347212415d3029f192c40152e8525a20b5c9bfed88ccdb32e) +
                      (({q0_1[167],q0_0[167]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[167],q0_0[167]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2f3612471464f3108bd427b6427c8fe79dce2b8e23dc4bb74cecb7e89a3b64a1  <=
                      (Ic5a87abf4c6018e9555de321c141d9754a7de91f1743d980e339ff9cebd63b7a) +
                      (({q0_1[168],q0_0[168]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[168],q0_0[168]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iccedefdcae7039447a6901e1cac8bf962a9f520d3b343c2b00e654c7e11a24f2  <=
                      (I3a27e4e3322c28e7fe85d7e76b7d5477f4d4f6acb8cdb876b9a54cba98b189b9) +
                      (({q0_1[169],q0_0[169]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[169],q0_0[169]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I8252bcef404ae08a2a748c98d672c368fbe4187f26e788e54d93af9077f92a20  <=
                      (I11edfeb948852dab396975b53b12d09da7a5fbedc2dae9fe7c687768cfef05b4) +
                      (({q0_1[170],q0_0[170]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[170],q0_0[170]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iaa2493521eb50d228c5b0619dca5c86b89a165f9855552ce98021778cc196f8d  <=
                      (I578437932d2d1156445b41a1238e0fd96ab5702bc3158ea337a9e37d14d6731e) +
                      (({q0_1[171],q0_0[171]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[171],q0_0[171]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I69d7f0497be77c5b1457ccdc35789d454bbe83f7d9eb458527d737a2222c7796  <=
                      (I3c2c5b5cd798851c7fcb0d0e66ddf81a516ef9bdf4aa4ebd4901532bfb2a651b) +
                      (({q0_1[172],q0_0[172]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[172],q0_0[172]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2c40224a96616b7749f39d78a0c07514232a019bf2c9ecd7340560f5aa5ce6bd  <=
                      (I8153d6f17d832da24daaba2909a88f1609e523ad3b6eac7ad42521979aae96da) +
                      (({q0_1[173],q0_0[173]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[173],q0_0[173]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id95e503df18410329be5e7761b6857182c75f7d2b0268d0fc377a415c89cad3f  <=
                      (Ic10ea001dcd0b864b987bc3080e95b338c1e91247bb90e884e161c926183fd2b) +
                      (({q0_1[174],q0_0[174]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[174],q0_0[174]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5cca65d1f11141b49a1136898dac8226cb1ec1654c8b8846471f1e4c36bcf3fc  <=
                      (I61efe7187a1aaa28235dacf68eb1e1dd97e7cb5900862790bb4d5872d7adbd67) +
                      (({q0_1[175],q0_0[175]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[175],q0_0[175]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6abf4748a0be2d4365fd1d9b53a44c3183015e1bdfb9a3f671eb5beed231eda1  <=
                      (I3c710fbd5e4dce0c97eb9da2d8e526f9d44d87fa75088c0421353614e6ef5da9) +
                      (({q0_1[176],q0_0[176]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[176],q0_0[176]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I56bb103437d88864c0ecd5bea1ab5a0313fef2b904c52adb559e19bef8f716bb  <=
                      (Ie02f677979058dda2291ddb93acd64f4461f6d75f3a33c21dac97129344f7055) +
                      (({q0_1[177],q0_0[177]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[177],q0_0[177]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5596d8fa3572e105a1618deba542906f0ba5acef8d7b0a48d0fe2e4eb3cf7481  <=
                      (I2b78100b50f7334d563daa27cab8078fa374dca0c438157d1ad44ed3fd9e3456) +
                      (({q0_1[178],q0_0[178]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[178],q0_0[178]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic00f466513895a54a6974af570c7bd5aba8c0ecab5612798bf512ca88f27081d  <=
                      (Icdfa68bdad11213dbaa576cbf43ca9deeb1f9f24225264eaeeede7d1aba5fd8a) +
                      (({q0_1[179],q0_0[179]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[179],q0_0[179]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I456f1fae558de9875bb1f76cfbb1840945f61ea1bce9c9bbcd0ead15d4b2803e  <=
                      (Idb39db95234cbfdbbc89fdee230784c703e170b9e932643a5e1b811b24ae021a) +
                      (({q0_1[180],q0_0[180]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[180],q0_0[180]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7b2c627cf9d530af8ad8ebc0d3dbc53988ea1819d98b5e36e1517e21cc954782  <=
                      (I7141b42fce475b5502fd33035bf37addde06271b2259e158ba03a66843b66075) +
                      (({q0_1[181],q0_0[181]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[181],q0_0[181]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic61cceb25c811577024c75e771c53089a2adb9f80e6a622eb82f9d8e5bbb6c16  <=
                      (I245e922da0aa5470370db389d5bc9db33327c905528a1740aa015b7ccdfcc29e) +
                      (({q0_1[182],q0_0[182]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[182],q0_0[182]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id8edf0b11a998a6c5737c8877c9b203e44c777ca9ee01cce63f046a6bd375c13  <=
                      (Ia2ff4d61c4f4fdf29be87b50e206c308cf970cbad2638e86ba8c2be8d025b534) +
                      (({q0_1[183],q0_0[183]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[183],q0_0[183]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2813295228131e78d6af31808dc1d9a6f712ddc60b2629d5329dc6ee2d07c9d9  <=
                      (Idd383630385363471e1b17ea946a61194a3cb287d833af386876c3b4ee66e406) +
                      (({q0_1[184],q0_0[184]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[184],q0_0[184]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I6736fca4e33cbc58b4658d91a401b558b1fbf9b3496e1830a8d7b4237d0ef125  <=
                      (I3daa8702e9dbd047a05e5ea044d14b670c2ae3849526cc514be6a511c5c45c35) +
                      (({q0_1[185],q0_0[185]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[185],q0_0[185]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Id66c49fe8c0d931dab1b901945cc3926c6e7e3d220480a28e0099a0656241a03  <=
                      (Ia695c63ae87e9a6742c6fecea648a214f5b24ea2b652bb5d83f35d9a59b94f72) +
                      (({q0_1[186],q0_0[186]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[186],q0_0[186]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I1d8a87a805073dbe04ce0f76953a234bceb3e6027b2a187071b492f644843715  <=
                      (Ifc31b600cbbf26e78cee82cd354c17b872586c1a53ddd132edbd25ce87d8aa9a) +
                      (({q0_1[187],q0_0[187]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[187],q0_0[187]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ieb9ae0dc5ee16583e8d05536052b61089e8004344fa0e3fdbc88c5af5119f293  <=
                      (I261e70e693cdbc572e40e81c594f3dac624febb03465bfd0fb864d337e753499) +
                      (({q0_1[188],q0_0[188]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[188],q0_0[188]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iff41f572ab79a4cc8e83538b32d4861e88ebdd0a9ce51555053943225158c5af  <=
                      (Ia6f7ae0adde8136c7a25f4fed69bbcaa376b5f28cbb4990afabb57a87ec03019) +
                      (({q0_1[189],q0_0[189]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[189],q0_0[189]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7f8fe2415810e04fccd129edfe956981aea020e4b24dd85d59991f4ef0131380  <=
                      (Ic40e94217a2d2c13f4b1ad2766ab1ae4e8ded0b5e0a3522dd51ec806c3e9feef) +
                      (({q0_1[190],q0_0[190]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[190],q0_0[190]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I5eafefae338dc0fdd7610a7cc3093d323fbd397263d3c8b7546bf540e77d60de  <=
                      (I78602c68a4a00f530bda7ba1dfa4820b7faeb0edabc636d6a2d8bf97005755d1) +
                      (({q0_1[191],q0_0[191]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[191],q0_0[191]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ie5d6a774e706204102b6a2d413e41c538f5e61284a19c7a47c42e356ea77d072  <=
                      (Id8e684d92e6d0b6e10b5e7f7ff9656e6fc67c99edaa59b49e453844ae33d23f6) +
                      (({q0_1[192],q0_0[192]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[192],q0_0[192]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Iab62db2e5fab6a7735067ea4afe23d7904f71c5b92219a1ea7848fa358da3cdd  <=
                      (Ic9d9001a209401fca8a3f28e39c4b89adc8f4e9d225aeffbb5d30893bea1a7b2) +
                      (({q0_1[193],q0_0[193]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[193],q0_0[193]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Icdf027acf32cc766a4ab1f19373a58cad87f74c1ca1791f66e958de6f18803ab  <=
                      (I97f666707f6afacfc6156ef498941fe5feeb7424834b4a283139aefb5f50a68f) +
                      (({q0_1[194],q0_0[194]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[194],q0_0[194]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib087093eca2530f923f55a4b4cddc83869730b169ab16bf26f6378b580da58f2  <=
                      (Ibdaeb96b71f9ccccfe79b1b3bab77122aa32217b58037d80a3183bf888b60c72) +
                      (({q0_1[195],q0_0[195]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[195],q0_0[195]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ice19f7340dbb41a6b126bdae27e69b813b5d6f73ba4db6ee79715328be678511  <=
                      (I574e4843ab81be7ad95cb7027fc3284a8780b07fb8a194a9c991997988d7ff8f) +
                      (({q0_1[196],q0_0[196]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[196],q0_0[196]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I575538bdc858fc8c843bc6b68625f1ba5fd33a904937071914caccc65f324a49  <=
                      (Iaa4463f258ed92a2c85fef0790c47e725c555f37c80dbe366d973c9599a5484d) +
                      (({q0_1[197],q0_0[197]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[197],q0_0[197]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Idea12ce0edfa5df65e47f6496f2a457a03907e9d62de2cb3797ec2cc6c5adf07  <=
                      (I7102386e760e34e2d0fc4563b497acec7222bd171333a2169fac800df94ea27c) +
                      (({q0_1[198],q0_0[198]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[198],q0_0[198]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib368839377e69cd28a997a22724c32efdc8820a04f9b5f93d9877bf398ec6e61  <=
                      (Iee34d958bf4feec1e5bde8a866a9919f29edd54f1bc51cc9c8216b71101d640b) +
                      (({q0_1[199],q0_0[199]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[199],q0_0[199]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I67be614a904dd4d47457ba0dc7a19b2e9f8e4231797917ef3610aea55d5ba3a8  <=
                      (I64b0ef6642050de0690c95be2af9606797be36c1656f1306b87ce3e8131c4629) +
                      (({q0_1[200],q0_0[200]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[200],q0_0[200]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I7cd598a52037f986959ad3f02b4b2783a613170f53a7e49573c5da74f1cbf614  <=
                      (I23f31ebee34c7f4f9c46fba41d41df176a7465c074ad8527205a5782edab6524) +
                      (({q0_1[201],q0_0[201]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[201],q0_0[201]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ide70b17967ff52e323b4a51db51e71445ad3c5483c745b2cec2cc338e5f42f6f  <=
                      (I628b9674d7d6caaa70c54539241df2e7a4be0441dde1739b442513c6e4ded8a4) +
                      (({q0_1[202],q0_0[202]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[202],q0_0[202]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ib28a3a83a3be0baf561a184b6de18de0c4847ff892c403bb9da441f017dd5efb  <=
                      (Ib066c9d790586949b27c4cf09dc957e7d28161ab00e8dc6920e4e0cc5ac665d9) +
                      (({q0_1[203],q0_0[203]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[203],q0_0[203]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2416ae27b898336a36264980b371003c06275245f514135d0adac28d88379cf7  <=
                      (I57419941b1979cd06c4fa0e6be943f004dd80da502425ee5b6dabd2239139cd7) +
                      (({q0_1[204],q0_0[204]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[204],q0_0[204]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I2d58b3296656a43e75a58883e59a576c0bf73dcd6bc28a939582be7ce0a0ffbd  <=
                      (Iabb5703a54942b1bdcfe2213d2011c659ec812f751dc75943b2ce511c81ffaf9) +
                      (({q0_1[205],q0_0[205]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[205],q0_0[205]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               I3f548241255df4c4a5a8b71a4352ffad6c3e5278c73de2b1afd1a1f1f1f94684  <=
                      (I798a6a6074b50fc61bd4e1b4696560abd2e515c86d47f85e9a3077cf6672acc8) +
                      (({q0_1[206],q0_0[206]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[206],q0_0[206]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"
               Ic3ef9d69272fb936b5ada08c6eb60ccaa6acf7b139689e5cb44e0ab76c0ee24c  <=
                      (I3f4a8ec7c554b1f0b9d3d2963b0e3dec4654bf07c5b836f8fd07c639cd19d588) +
                      (({q0_1[207],q0_0[207]} ==2'b11) ? ~percent_probability_int + 1 : (( {q0_1[207],q0_0[207]}  == 2'b01) ? percent_probability_int : 32'h0));
                    // 2'b11 === -1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b1
                    // 2'b01 ===  1 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for 1'b0
                    // 2'b00 ===  Ia4888af4e46c129c695ee32775a8c233f113c82e7cd4e6fd3cbb1fda5659f36a I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 -1:1 and 1:0 I51a733b740d2bdbf4b02ea2ec24007ef3cf36ab9b6261a3003ed24730acc888a I77bc06c55d29ee3cfa295b4592e4b2a85a16bb06a8974726b7bfa3d4ca36d5ae Ifa51fd49abf67705d6a35d18218c115ff5633aec1f9ebfdc9d5d4956416f57f6 bit Icd42404d52ad55ccfa9aca4adc828aa5800ad9d385a0671fbcbf724118320619 for "Ib23a6a8439c0dde5515893e7c90c1e3233b8616e634470f20dc4928bcf3609bc"

                 if ({q0_1[0],q0_0[0]} != 1 ) begin
                 end
                 if ({q0_1[1],q0_0[1]} != 1 ) begin
                 end
                 if ({q0_1[2],q0_0[2]} != 0 ) begin
                 end
                 if ({q0_1[3],q0_0[3]} != 1 ) begin
                 end
                 if ({q0_1[4],q0_0[4]} != 0 ) begin
                 end
                 if ({q0_1[5],q0_0[5]} != 0 ) begin
                 end
                 if ({q0_1[6],q0_0[6]} != 0 ) begin
                 end
                 if ({q0_1[7],q0_0[7]} != 0 ) begin
                 end
                 if ({q0_1[8],q0_0[8]} != 0 ) begin
                 end
                 if ({q0_1[9],q0_0[9]} != 1 ) begin
                 end
                 if ({q0_1[10],q0_0[10]} != 1 ) begin
                 end
                 if ({q0_1[11],q0_0[11]} != 1 ) begin
                 end
                 if ({q0_1[12],q0_0[12]} != 1 ) begin
                 end
                 if ({q0_1[13],q0_0[13]} != 1 ) begin
                 end
                 if ({q0_1[14],q0_0[14]} != 0 ) begin
                 end
                 if ({q0_1[15],q0_0[15]} != 1 ) begin
                 end
                 if ({q0_1[16],q0_0[16]} != 0 ) begin
                 end
                 if ({q0_1[17],q0_0[17]} != 0 ) begin
                 end
                 if ({q0_1[18],q0_0[18]} != 1 ) begin
                 end
                 if ({q0_1[19],q0_0[19]} != 0 ) begin
                 end
                 if ({q0_1[20],q0_0[20]} != 1 ) begin
                 end
                 if ({q0_1[21],q0_0[21]} != 1 ) begin
                 end
                 if ({q0_1[22],q0_0[22]} != 0 ) begin
                 end
                 if ({q0_1[23],q0_0[23]} != 0 ) begin
                 end
                 if ({q0_1[24],q0_0[24]} != 0 ) begin
                 end
                 if ({q0_1[25],q0_0[25]} != 1 ) begin
                 end
                 if ({q0_1[26],q0_0[26]} != 1 ) begin
                 end
                 if ({q0_1[27],q0_0[27]} != 0 ) begin
                 end
                 if ({q0_1[28],q0_0[28]} != 0 ) begin
                 end
                 if ({q0_1[29],q0_0[29]} != 1 ) begin
                 end
                 if ({q0_1[30],q0_0[30]} != 1 ) begin
                 end
                 if ({q0_1[31],q0_0[31]} != 1 ) begin
                 end
                 if ({q0_1[32],q0_0[32]} != 0 ) begin
                 end
                 if ({q0_1[33],q0_0[33]} != 0 ) begin
                 end
                 if ({q0_1[34],q0_0[34]} != 1 ) begin
                 end
                 if ({q0_1[35],q0_0[35]} != 0 ) begin
                 end
                 if ({q0_1[36],q0_0[36]} != 0 ) begin
                 end
                 if ({q0_1[37],q0_0[37]} != 0 ) begin
                 end
                 if ({q0_1[38],q0_0[38]} != 0 ) begin
                 end
                 if ({q0_1[39],q0_0[39]} != 0 ) begin
                 end
                 if ({q0_1[40],q0_0[40]} != 1 ) begin
                 end
                 if ({q0_1[41],q0_0[41]} != 0 ) begin
                 end
                 if ({q0_1[42],q0_0[42]} != 0 ) begin
                 end
                 if ({q0_1[43],q0_0[43]} != 1 ) begin
                 end
                 if ({q0_1[44],q0_0[44]} != 1 ) begin
                 end
                 if ({q0_1[45],q0_0[45]} != 1 ) begin
                 end
                 if ({q0_1[46],q0_0[46]} != 1 ) begin
                 end
                 if ({q0_1[47],q0_0[47]} != 0 ) begin
                 end
                 if ({q0_1[48],q0_0[48]} != 0 ) begin
                 end
                 if ({q0_1[49],q0_0[49]} != 1 ) begin
                 end
                 if ({q0_1[50],q0_0[50]} != 1 ) begin
                 end
                 if ({q0_1[51],q0_0[51]} != 0 ) begin
                 end
                 if ({q0_1[52],q0_0[52]} != 1 ) begin
                 end
                 if ({q0_1[53],q0_0[53]} != 1 ) begin
                 end
                 if ({q0_1[54],q0_0[54]} != 0 ) begin
                 end
                 if ({q0_1[55],q0_0[55]} != 1 ) begin
                 end
                 if ({q0_1[56],q0_0[56]} != 1 ) begin
                 end
                 if ({q0_1[57],q0_0[57]} != 0 ) begin
                 end
                 if ({q0_1[58],q0_0[58]} != 0 ) begin
                 end
                 if ({q0_1[59],q0_0[59]} != 1 ) begin
                 end
                 if ({q0_1[60],q0_0[60]} != 0 ) begin
                 end
                 if ({q0_1[61],q0_0[61]} != 0 ) begin
                 end
                 if ({q0_1[62],q0_0[62]} != 0 ) begin
                 end
                 if ({q0_1[63],q0_0[63]} != 1 ) begin
                 end
                 if ({q0_1[64],q0_0[64]} != 0 ) begin
                 end
                 if ({q0_1[65],q0_0[65]} != 1 ) begin
                 end
                 if ({q0_1[66],q0_0[66]} != 1 ) begin
                 end
                 if ({q0_1[67],q0_0[67]} != 1 ) begin
                 end
                 if ({q0_1[68],q0_0[68]} != 1 ) begin
                 end
                 if ({q0_1[69],q0_0[69]} != 1 ) begin
                 end
                 if ({q0_1[70],q0_0[70]} != 1 ) begin
                 end
                 if ({q0_1[71],q0_0[71]} != 1 ) begin
                 end
                 if ({q0_1[72],q0_0[72]} != 0 ) begin
                 end
                 if ({q0_1[73],q0_0[73]} != 0 ) begin
                 end
                 if ({q0_1[74],q0_0[74]} != 1 ) begin
                 end
                 if ({q0_1[75],q0_0[75]} != 0 ) begin
                 end
                 if ({q0_1[76],q0_0[76]} != 0 ) begin
                 end
                 if ({q0_1[77],q0_0[77]} != 0 ) begin
                 end
                 if ({q0_1[78],q0_0[78]} != 0 ) begin
                 end
                 if ({q0_1[79],q0_0[79]} != 0 ) begin
                 end
                 if ({q0_1[80],q0_0[80]} != 0 ) begin
                 end
                 if ({q0_1[81],q0_0[81]} != 1 ) begin
                 end
                 if ({q0_1[82],q0_0[82]} != 1 ) begin
                 end
                 if ({q0_1[83],q0_0[83]} != 0 ) begin
                 end
                 if ({q0_1[84],q0_0[84]} != 0 ) begin
                 end
                 if ({q0_1[85],q0_0[85]} != 0 ) begin
                 end
                 if ({q0_1[86],q0_0[86]} != 0 ) begin
                 end
                 if ({q0_1[87],q0_0[87]} != 0 ) begin
                 end
                 if ({q0_1[88],q0_0[88]} != 0 ) begin
                 end
                 if ({q0_1[89],q0_0[89]} != 1 ) begin
                 end
                 if ({q0_1[90],q0_0[90]} != 0 ) begin
                 end
                 if ({q0_1[91],q0_0[91]} != 1 ) begin
                 end
                 if ({q0_1[92],q0_0[92]} != 0 ) begin
                 end
                 if ({q0_1[93],q0_0[93]} != 0 ) begin
                 end
                 if ({q0_1[94],q0_0[94]} != 0 ) begin
                 end
                 if ({q0_1[95],q0_0[95]} != 0 ) begin
                 end
                 if ({q0_1[96],q0_0[96]} != 0 ) begin
                 end
                 if ({q0_1[97],q0_0[97]} != 0 ) begin
                 end
                 if ({q0_1[98],q0_0[98]} != 0 ) begin
                 end
                 if ({q0_1[99],q0_0[99]} != 0 ) begin
                 end
                 if ({q0_1[100],q0_0[100]} != 1 ) begin
                 end
                 if ({q0_1[101],q0_0[101]} != 1 ) begin
                 end
                 if ({q0_1[102],q0_0[102]} != 1 ) begin
                 end
                 if ({q0_1[103],q0_0[103]} != 1 ) begin
                 end
                 if ({q0_1[104],q0_0[104]} != 0 ) begin
                 end
                 if ({q0_1[105],q0_0[105]} != 1 ) begin
                 end
                 if ({q0_1[106],q0_0[106]} != 1 ) begin
                 end
                 if ({q0_1[107],q0_0[107]} != 1 ) begin
                 end
                 if ({q0_1[108],q0_0[108]} != 0 ) begin
                 end
                 if ({q0_1[109],q0_0[109]} != 0 ) begin
                 end
                 if ({q0_1[110],q0_0[110]} != 0 ) begin
                 end
                 if ({q0_1[111],q0_0[111]} != 1 ) begin
                 end
                 if ({q0_1[112],q0_0[112]} != 1 ) begin
                 end
                 if ({q0_1[113],q0_0[113]} != 0 ) begin
                 end
                 if ({q0_1[114],q0_0[114]} != 0 ) begin
                 end
                 if ({q0_1[115],q0_0[115]} != 1 ) begin
                 end
                 if ({q0_1[116],q0_0[116]} != 1 ) begin
                 end
                 if ({q0_1[117],q0_0[117]} != 1 ) begin
                 end
                 if ({q0_1[118],q0_0[118]} != 1 ) begin
                 end
                 if ({q0_1[119],q0_0[119]} != 0 ) begin
                 end
                 if ({q0_1[120],q0_0[120]} != 1 ) begin
                 end
                 if ({q0_1[121],q0_0[121]} != 0 ) begin
                 end
                 if ({q0_1[122],q0_0[122]} != 0 ) begin
                 end
                 if ({q0_1[123],q0_0[123]} != 1 ) begin
                 end
                 if ({q0_1[124],q0_0[124]} != 0 ) begin
                 end
                 if ({q0_1[125],q0_0[125]} != 0 ) begin
                 end
                 if ({q0_1[126],q0_0[126]} != 1 ) begin
                 end
                 if ({q0_1[127],q0_0[127]} != 1 ) begin
                 end
                 if ({q0_1[128],q0_0[128]} != 1 ) begin
                 end
                 if ({q0_1[129],q0_0[129]} != 0 ) begin
                 end
                 if ({q0_1[130],q0_0[130]} != 1 ) begin
                 end
                 if ({q0_1[131],q0_0[131]} != 0 ) begin
                 end
                 if ({q0_1[132],q0_0[132]} != 0 ) begin
                 end
                 if ({q0_1[133],q0_0[133]} != 0 ) begin
                 end
                 if ({q0_1[134],q0_0[134]} != 1 ) begin
                 end
                 if ({q0_1[135],q0_0[135]} != 1 ) begin
                 end
                 if ({q0_1[136],q0_0[136]} != 1 ) begin
                 end
                 if ({q0_1[137],q0_0[137]} != 0 ) begin
                 end
                 if ({q0_1[138],q0_0[138]} != 1 ) begin
                 end
                 if ({q0_1[139],q0_0[139]} != 1 ) begin
                 end
                 if ({q0_1[140],q0_0[140]} != 1 ) begin
                 end
                 if ({q0_1[141],q0_0[141]} != 0 ) begin
                 end
                 if ({q0_1[142],q0_0[142]} != 0 ) begin
                 end
                 if ({q0_1[143],q0_0[143]} != 1 ) begin
                 end
                 if ({q0_1[144],q0_0[144]} != 0 ) begin
                 end
                 if ({q0_1[145],q0_0[145]} != 1 ) begin
                 end
                 if ({q0_1[146],q0_0[146]} != 0 ) begin
                 end
                 if ({q0_1[147],q0_0[147]} != 1 ) begin
                 end
                 if ({q0_1[148],q0_0[148]} != 1 ) begin
                 end
                 if ({q0_1[149],q0_0[149]} != 1 ) begin
                 end
                 if ({q0_1[150],q0_0[150]} != 1 ) begin
                 end
                 if ({q0_1[151],q0_0[151]} != 0 ) begin
                 end
                 if ({q0_1[152],q0_0[152]} != 1 ) begin
                 end
                 if ({q0_1[153],q0_0[153]} != 0 ) begin
                 end
                 if ({q0_1[154],q0_0[154]} != 0 ) begin
                 end
                 if ({q0_1[155],q0_0[155]} != 0 ) begin
                 end
                 if ({q0_1[156],q0_0[156]} != 0 ) begin
                 end
                 if ({q0_1[157],q0_0[157]} != 1 ) begin
                 end
                 if ({q0_1[158],q0_0[158]} != 0 ) begin
                 end
                 if ({q0_1[159],q0_0[159]} != 1 ) begin
                 end
                 if ({q0_1[160],q0_0[160]} != 1 ) begin
                 end
                 if ({q0_1[161],q0_0[161]} != 0 ) begin
                 end
                 if ({q0_1[162],q0_0[162]} != 0 ) begin
                 end
                 if ({q0_1[163],q0_0[163]} != 1 ) begin
                 end
                 if ({q0_1[164],q0_0[164]} != 0 ) begin
                 end
                 if ({q0_1[165],q0_0[165]} != 0 ) begin
                 end
                 if ({q0_1[166],q0_0[166]} != 1 ) begin
                 end
                 if ({q0_1[167],q0_0[167]} != 1 ) begin
                 end
                 if ({q0_1[168],q0_0[168]} != 0 ) begin
                 end
                 if ({q0_1[169],q0_0[169]} != 0 ) begin
                 end
                 if ({q0_1[170],q0_0[170]} != 1 ) begin
                 end
                 if ({q0_1[171],q0_0[171]} != 0 ) begin
                 end
                 if ({q0_1[172],q0_0[172]} != 1 ) begin
                 end
                 if ({q0_1[173],q0_0[173]} != 1 ) begin
                 end
                 if ({q0_1[174],q0_0[174]} != 0 ) begin
                 end
                 if ({q0_1[175],q0_0[175]} != 0 ) begin
                 end
                 if ({q0_1[176],q0_0[176]} != 1 ) begin
                 end
                 if ({q0_1[177],q0_0[177]} != 0 ) begin
                 end
                 if ({q0_1[178],q0_0[178]} != 1 ) begin
                 end
                 if ({q0_1[179],q0_0[179]} != 1 ) begin
                 end
                 if ({q0_1[180],q0_0[180]} != 1 ) begin
                 end
                 if ({q0_1[181],q0_0[181]} != 0 ) begin
                 end
                 if ({q0_1[182],q0_0[182]} != 1 ) begin
                 end
                 if ({q0_1[183],q0_0[183]} != 1 ) begin
                 end
                 if ({q0_1[184],q0_0[184]} != 1 ) begin
                 end
                 if ({q0_1[185],q0_0[185]} != 1 ) begin
                 end
                 if ({q0_1[186],q0_0[186]} != 0 ) begin
                 end
                 if ({q0_1[187],q0_0[187]} != 1 ) begin
                 end
                 if ({q0_1[188],q0_0[188]} != 0 ) begin
                 end
                 if ({q0_1[189],q0_0[189]} != 0 ) begin
                 end
                 if ({q0_1[190],q0_0[190]} != 0 ) begin
                 end
                 if ({q0_1[191],q0_0[191]} != 0 ) begin
                 end
                 if ({q0_1[192],q0_0[192]} != 1 ) begin
                 end
                 if ({q0_1[193],q0_0[193]} != 0 ) begin
                 end
                 if ({q0_1[194],q0_0[194]} != 0 ) begin
                 end
                 if ({q0_1[195],q0_0[195]} != 0 ) begin
                 end
                 if ({q0_1[196],q0_0[196]} != 0 ) begin
                 end
                 if ({q0_1[197],q0_0[197]} != 0 ) begin
                 end
                 if ({q0_1[198],q0_0[198]} != 0 ) begin
                 end
                 if ({q0_1[199],q0_0[199]} != 0 ) begin
                 end
                 if ({q0_1[200],q0_0[200]} != 0 ) begin
                 end
                 if ({q0_1[201],q0_0[201]} != 0 ) begin
                 end
                 if ({q0_1[202],q0_0[202]} != 1 ) begin
                 end
                 if ({q0_1[203],q0_0[203]} != 0 ) begin
                 end
                 if ({q0_1[204],q0_0[204]} != 0 ) begin
                 end
                 if ({q0_1[205],q0_0[205]} != 0 ) begin
                 end
                 if ({q0_1[206],q0_0[206]} != 1 ) begin
                 end
                 if ({q0_1[207],q0_0[207]} != 0 ) begin
                 end


           end

           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[0]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[0] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[0] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[0]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[1]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[1] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[1] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[1]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[2]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[2] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[2] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[2]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[3]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[3] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[3] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[3]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[4]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[4] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[4] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[4]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[5]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[5] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[5] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[5]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[6]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[6] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[6] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[6]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[7]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[7] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[7] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[7]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[8]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[8] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[8] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[8]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[9]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[9] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[9] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[9]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[10]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[10] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[10] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[10]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[11]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[11] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[11] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[11]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[12]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[12] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[12] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[12]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[13]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[13] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[13] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[13]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[14]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[14] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[14] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[14]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[15]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[15] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[15] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[15]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[16]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[16] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[16] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[16]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[17]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[17] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[17] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[17]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[18]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[18] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[18] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[18]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[19]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[19] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[19] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[19]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[20]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[20] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[20] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[20]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[21]        <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[21] + 1 :
                                             I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[21] ;
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[21]  <=  I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[0]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[0] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[0] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[0]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[1]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[1] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[1] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[1]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[2]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[2] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[2] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[2]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[3]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[3] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[3] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[3]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[4]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[4] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[4] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[4]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[5]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[5] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[5] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[5]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[6]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[6] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[6] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[6]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[7]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[7] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[7] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[7]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[8]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[8] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[8] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[8]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[9]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[9] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[9] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[9]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[10]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[10] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[10] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[10]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[11]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[11] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[11] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[11]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[12]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[12] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[12] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[12]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[13]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[13] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[13] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[13]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[14]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[14] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[14] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[14]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[15]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[15] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[15] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[15]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[16]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[16] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[16] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[16]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[17]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[17] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[17] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[17]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[18]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[18] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[18] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[18]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[19]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[19] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[19] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[19]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[20]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[20] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[20] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[20]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[21]        <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[21] + 1 :
                                             I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[21] ;
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[21]  <=  I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[0]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[0] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[0] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[0]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[1]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[1] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[1] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[1]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[2]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[2] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[2] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[2]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[3]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[3] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[3] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[3]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[4]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[4] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[4] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[4]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[5]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[5] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[5] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[5]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[6]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[6] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[6] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[6]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[7]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[7] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[7] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[7]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[8]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[8] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[8] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[8]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[9]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[9] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[9] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[9]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[10]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[10] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[10] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[10]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[11]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[11] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[11] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[11]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[12]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[12] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[12] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[12]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[13]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[13] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[13] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[13]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[14]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[14] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[14] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[14]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[15]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[15] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[15] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[15]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[16]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[16] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[16] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[16]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[17]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[17] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[17] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[17]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[18]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[18] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[18] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[18]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[19]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[19] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[19] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[19]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[20]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[20] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[20] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[20]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[21]        <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[21] + 1 :
                                             I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[21] ;
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[21]  <=  I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[0]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[0] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[0] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[0]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[1]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[1] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[1] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[1]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[2]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[2] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[2] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[2]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[3]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[3] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[3] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[3]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[4]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[4] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[4] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[4]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[5]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[5] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[5] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[5]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[6]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[6] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[6] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[6]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[7]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[7] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[7] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[7]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[8]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[8] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[8] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[8]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[9]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[9] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[9] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[9]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[10]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[10] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[10] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[10]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[11]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[11] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[11] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[11]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[12]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[12] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[12] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[12]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[13]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[13] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[13] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[13]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[14]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[14] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[14] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[14]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[15]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[15] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[15] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[15]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[16]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[16] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[16] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[16]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[17]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[17] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[17] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[17]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[18]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[18] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[18] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[18]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[19]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[19] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[19] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[19]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[20]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[20] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[20] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[20]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[21]        <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[21] + 1 :
                                             Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[21] ;
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[21]  <=  Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[0]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[0] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[0] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[0]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[1]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[1] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[1] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[1]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[2]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[2] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[2] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[2]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[3]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[3] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[3] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[3]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[4]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[4] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[4] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[4]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[5]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[5] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[5] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[5]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[6]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[6] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[6] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[6]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[7]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[7] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[7] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[7]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[8]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[8] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[8] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[8]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[9]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[9] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[9] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[9]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[10]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[10] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[10] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[10]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[11]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[11] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[11] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[11]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[12]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[12] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[12] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[12]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[13]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[13] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[13] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[13]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[14]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[14] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[14] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[14]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[15]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[15] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[15] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[15]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[16]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[16] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[16] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[16]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[17]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[17] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[17] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[17]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[18]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[18] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[18] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[18]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[19]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[19] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[19] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[19]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[20]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[20] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[20] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[20]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[21]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[21] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[21] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[21]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[22]        <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[22][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[22] + 1 :
                                             Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[22] ;
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[22]  <=  Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[22][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[0]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[0] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[0] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[0]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[1]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[1] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[1] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[1]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[2]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[2] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[2] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[2]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[3]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[3] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[3] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[3]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[4]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[4] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[4] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[4]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[5]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[5] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[5] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[5]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[6]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[6] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[6] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[6]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[7]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[7] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[7] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[7]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[8]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[8] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[8] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[8]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[9]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[9] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[9] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[9]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[10]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[10] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[10] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[10]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[11]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[11] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[11] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[11]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[12]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[12] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[12] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[12]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[13]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[13] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[13] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[13]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[14]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[14] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[14] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[14]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[15]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[15] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[15] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[15]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[16]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[16] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[16] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[16]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[17]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[17] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[17] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[17]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[18]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[18] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[18] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[18]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[19]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[19] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[19] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[19]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[20]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[20] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[20] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[20]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[21]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[21] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[21] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[21]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[22]        <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[22][MAX_SUM_WDTH_LONG-1] ?
                                             ~I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[22] + 1 :
                                             I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[22] ;
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[22]  <=  I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[22][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[0]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[0] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[0] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[0]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[1]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[1] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[1] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[1]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[2]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[2] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[2] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[2]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[3]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[3] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[3] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[3]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[4]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[4] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[4] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[4]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[5]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[5] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[5] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[5]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[6]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[6] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[6] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[6]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[7]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[7] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[7] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[7]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[8]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[8] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[8] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[8]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[9]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[9] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[9] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[9]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[10]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[10] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[10] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[10]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[11]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[11] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[11] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[11]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[12]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[12] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[12] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[12]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[13]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[13] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[13] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[13]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[14]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[14] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[14] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[14]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[15]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[15] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[15] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[15]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[16]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[16] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[16] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[16]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[17]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[17] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[17] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[17]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[18]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[18] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[18] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[18]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[19]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[19] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[19] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[19]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[20]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[20] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[20] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[20]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[21]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[21] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[21] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[21]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[22]        <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[22][MAX_SUM_WDTH_LONG-1] ?
                                             ~I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[22] + 1 :
                                             I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[22] ;
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[22]  <=  I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[22][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[0]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[0] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[0] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[0]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[1]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[1] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[1] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[1]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[2]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[2] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[2] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[2]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[3]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[3] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[3] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[3]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[4]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[4] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[4] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[4]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[5]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[5] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[5] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[5]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[6]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[6] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[6] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[6]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[7]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[7] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[7] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[7]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[8]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[8] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[8] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[8]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[9]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[9] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[9] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[9]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[10]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[10] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[10] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[10]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[11]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[11] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[11] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[11]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[12]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[12] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[12] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[12]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[13]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[13] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[13] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[13]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[14]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[14] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[14] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[14]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[15]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[15] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[15] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[15]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[16]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[16][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[16] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[16] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[16]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[16][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[17]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[17][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[17] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[17] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[17]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[17][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[18]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[18][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[18] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[18] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[18]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[18][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[19]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[19][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[19] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[19] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[19]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[19][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[20]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[20][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[20] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[20] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[20]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[20][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[21]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[21][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[21] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[21] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[21]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[21][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[22]        <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[22][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[22] + 1 :
                                             I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[22] ;
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[22]  <=  I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[22][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[0]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[0] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[0] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[0]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[1]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[1] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[1] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[1]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[2]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[2] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[2] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[2]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[3]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[3] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[3] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[3]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[4]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[4] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[4] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[4]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[5]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[5] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[5] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[5]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[6]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[6] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[6] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[6]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[7]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[7] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[7] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[7]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[8]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[8] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[8] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[8]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[9]        <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[9] + 1 :
                                             Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[9] ;
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[9]  <=  Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[0]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[0] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[0] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[0]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[1]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[1] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[1] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[1]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[2]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[2] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[2] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[2]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[3]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[3] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[3] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[3]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[4]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[4] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[4] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[4]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[5]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[5] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[5] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[5]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[6]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[6] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[6] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[6]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[7]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[7] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[7] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[7]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[8]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[8] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[8] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[8]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[9]        <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[9] + 1 :
                                             I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[9] ;
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[9]  <=  I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[0]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[0] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[0] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[0]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[1]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[1] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[1] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[1]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[2]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[2] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[2] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[2]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[3]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[3] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[3] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[3]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[4]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[4] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[4] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[4]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[5]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[5] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[5] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[5]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[6]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[6] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[6] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[6]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[7]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[7] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[7] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[7]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[8]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[8] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[8] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[8]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[9]        <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[9] + 1 :
                                             Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[9] ;
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[9]  <=  Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[0]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[0] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[0] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[0]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[1]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[1] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[1] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[1]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[2]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[2] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[2] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[2]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[3]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[3] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[3] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[3]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[4]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[4] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[4] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[4]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[5]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[5] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[5] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[5]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[6]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[6] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[6] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[6]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[7]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[7] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[7] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[7]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[8]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[8] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[8] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[8]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[9]        <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[9] + 1 :
                                             Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[9] ;
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[9]  <=  Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[0]        <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[0] + 1 :
                                             Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[0] ;
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[0]  <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[1]        <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[1] + 1 :
                                             Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[1] ;
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[1]  <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[2]        <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[2] + 1 :
                                             Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[2] ;
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[2]  <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[3]        <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[3] + 1 :
                                             Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[3] ;
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[3]  <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[4]        <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[4] + 1 :
                                             Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[4] ;
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[4]  <=  Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[0]        <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[0] + 1 :
                                             Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[0] ;
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[0]  <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[1]        <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[1] + 1 :
                                             Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[1] ;
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[1]  <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[2]        <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[2] + 1 :
                                             Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[2] ;
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[2]  <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[3]        <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[3] + 1 :
                                             Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[3] ;
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[3]  <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[4]        <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[4] + 1 :
                                             Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[4] ;
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[4]  <=  Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[0]        <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[0] + 1 :
                                             Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[0] ;
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[0]  <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[1]        <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[1] + 1 :
                                             Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[1] ;
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[1]  <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[2]        <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[2] + 1 :
                                             Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[2] ;
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[2]  <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[3]        <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[3] + 1 :
                                             Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[3] ;
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[3]  <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[4]        <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[4] + 1 :
                                             Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[4] ;
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[4]  <=  Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[0]        <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[0] + 1 :
                                             I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[0] ;
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[0]  <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[1]        <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[1] + 1 :
                                             I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[1] ;
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[1]  <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[2]        <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[2] + 1 :
                                             I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[2] ;
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[2]  <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[3]        <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[3] + 1 :
                                             I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[3] ;
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[3]  <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[4]        <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[4] + 1 :
                                             I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[4] ;
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[4]  <=  I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[0]        <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[0] + 1 :
                                             I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[0] ;
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[0]  <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[1]        <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[1] + 1 :
                                             I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[1] ;
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[1]  <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[2]        <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[2] + 1 :
                                             I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[2] ;
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[2]  <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[3]        <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[3] + 1 :
                                             I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[3] ;
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[3]  <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[4]        <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[4] + 1 :
                                             I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[4] ;
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[4]  <=  I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[0]        <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[0] + 1 :
                                             I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[0] ;
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[0]  <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[1]        <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[1] + 1 :
                                             I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[1] ;
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[1]  <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[2]        <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[2] + 1 :
                                             I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[2] ;
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[2]  <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[3]        <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[3] + 1 :
                                             I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[3] ;
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[3]  <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[4]        <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[4] + 1 :
                                             I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[4] ;
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[4]  <=  I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[0]        <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[0] + 1 :
                                             I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[0] ;
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[0]  <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[1]        <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[1] + 1 :
                                             I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[1] ;
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[1]  <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[2]        <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[2] + 1 :
                                             I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[2] ;
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[2]  <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[3]        <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[3] + 1 :
                                             I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[3] ;
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[3]  <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[4]        <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[4] + 1 :
                                             I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[4] ;
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[4]  <=  I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[0]        <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[0] + 1 :
                                             Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[0] ;
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[0]  <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[1]        <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[1] + 1 :
                                             Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[1] ;
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[1]  <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[2]        <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[2] + 1 :
                                             Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[2] ;
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[2]  <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[3]        <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[3] + 1 :
                                             Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[3] ;
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[3]  <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[4]        <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[4] + 1 :
                                             Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[4] ;
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[4]  <=  Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[0]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[0] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[0] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[0]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[1]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[1] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[1] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[1]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[2]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[2] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[2] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[2]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[3]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[3] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[3] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[3]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[4]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[4] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[4] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[4]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[5]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[5] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[5] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[5]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[6]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[6] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[6] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[6]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[7]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[7] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[7] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[7]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[8]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[8] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[8] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[8]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[9]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[9] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[9] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[9]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[10]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[10] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[10] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[10]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[11]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[11] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[11] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[11]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[12]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[12] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[12] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[12]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[13]        <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[13] + 1 :
                                             I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[13] ;
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[13]  <=  I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[0]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[0] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[0] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[0]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[1]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[1] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[1] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[1]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[2]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[2] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[2] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[2]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[3]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[3] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[3] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[3]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[4]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[4] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[4] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[4]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[5]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[5] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[5] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[5]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[6]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[6] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[6] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[6]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[7]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[7] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[7] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[7]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[8]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[8] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[8] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[8]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[9]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[9] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[9] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[9]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[10]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[10] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[10] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[10]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[11]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[11] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[11] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[11]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[12]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[12] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[12] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[12]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[13]        <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[13] + 1 :
                                             Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[13] ;
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[13]  <=  Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[0]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[0] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[0] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[0]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[1]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[1] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[1] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[1]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[2]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[2] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[2] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[2]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[3]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[3] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[3] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[3]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[4]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[4] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[4] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[4]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[5]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[5] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[5] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[5]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[6]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[6] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[6] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[6]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[7]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[7] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[7] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[7]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[8]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[8] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[8] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[8]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[9]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[9] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[9] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[9]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[10]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[10] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[10] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[10]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[11]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[11] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[11] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[11]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[12]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[12] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[12] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[12]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[13]        <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[13] + 1 :
                                             I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[13] ;
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[13]  <=  I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[0]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[0] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[0] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[0]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[1]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[1] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[1] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[1]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[2]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[2] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[2] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[2]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[3]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[3] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[3] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[3]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[4]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[4] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[4] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[4]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[5]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[5] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[5] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[5]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[6]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[6] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[6] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[6]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[7]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[7] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[7] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[7]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[8]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[8] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[8] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[8]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[9]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[9] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[9] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[9]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[10]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[10] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[10] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[10]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[11]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[11] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[11] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[11]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[12]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[12] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[12] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[12]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[13]        <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[13] + 1 :
                                             I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[13] ;
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[13]  <=  I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[0]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[0] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[0] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[0]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[1]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[1] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[1] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[1]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[2]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[2] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[2] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[2]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[3]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[3] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[3] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[3]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[4]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[4] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[4] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[4]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[5]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[5] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[5] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[5]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[6]        <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[6] + 1 :
                                             I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[6] ;
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[6]  <=  I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[0]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[0] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[0] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[0]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[1]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[1] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[1] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[1]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[2]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[2] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[2] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[2]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[3]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[3] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[3] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[3]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[4]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[4] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[4] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[4]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[5]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[5] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[5] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[5]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[6]        <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[6] + 1 :
                                             I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[6] ;
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[6]  <=  I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[0]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[0] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[0] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[0]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[1]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[1] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[1] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[1]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[2]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[2] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[2] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[2]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[3]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[3] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[3] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[3]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[4]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[4] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[4] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[4]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[5]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[5] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[5] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[5]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[6]        <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[6] + 1 :
                                             Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[6] ;
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[6]  <=  Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[0]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[0] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[0] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[0]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[1]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[1] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[1] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[1]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[2]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[2] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[2] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[2]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[3]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[3] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[3] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[3]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[4]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[4] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[4] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[4]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[5]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[5] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[5] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[5]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[6]        <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[6] + 1 :
                                             Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[6] ;
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[6]  <=  Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[0]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[0] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[0] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[0]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[1]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[1] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[1] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[1]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[2]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[2] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[2] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[2]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[3]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[3] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[3] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[3]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[4]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[4] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[4] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[4]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[5]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[5] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[5] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[5]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[6]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[6] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[6] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[6]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[7]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[7] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[7] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[7]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[8]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[8] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[8] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[8]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[9]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[9] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[9] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[9]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[10]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[10] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[10] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[10]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[11]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[11] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[11] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[11]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[12]        <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[12] + 1 :
                                             Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[12] ;
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[12]  <=  Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[0]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[0] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[0] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[0]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[1]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[1] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[1] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[1]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[2]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[2] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[2] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[2]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[3]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[3] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[3] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[3]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[4]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[4] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[4] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[4]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[5]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[5] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[5] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[5]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[6]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[6] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[6] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[6]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[7]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[7] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[7] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[7]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[8]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[8] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[8] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[8]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[9]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[9] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[9] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[9]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[10]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[10] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[10] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[10]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[11]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[11] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[11] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[11]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[12]        <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[12] + 1 :
                                             Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[12] ;
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[12]  <=  Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[0]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[0] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[0] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[0]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[1]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[1] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[1] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[1]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[2]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[2] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[2] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[2]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[3]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[3] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[3] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[3]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[4]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[4] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[4] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[4]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[5]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[5] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[5] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[5]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[6]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[6] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[6] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[6]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[7]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[7] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[7] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[7]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[8]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[8] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[8] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[8]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[9]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[9] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[9] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[9]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[10]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[10] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[10] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[10]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[11]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[11] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[11] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[11]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[12]        <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[12] + 1 :
                                             Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[12] ;
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[12]  <=  Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[0]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[0] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[0] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[0]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[1]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[1] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[1] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[1]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[2]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[2] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[2] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[2]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[3]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[3] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[3] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[3]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[4]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[4] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[4] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[4]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[5]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[5] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[5] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[5]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[6]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[6] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[6] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[6]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[7]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[7] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[7] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[7]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[8]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[8] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[8] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[8]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[9]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[9] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[9] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[9]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[10]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[10] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[10] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[10]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[11]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[11] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[11] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[11]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[12]        <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[12] + 1 :
                                             I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[12] ;
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[12]  <=  I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[0]        <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[0] + 1 :
                                             Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[0] ;
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[0]  <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[1]        <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[1] + 1 :
                                             Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[1] ;
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[1]  <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[2]        <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[2] + 1 :
                                             Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[2] ;
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[2]  <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[3]        <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[3] + 1 :
                                             Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[3] ;
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[3]  <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[4]        <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[4] + 1 :
                                             Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[4] ;
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[4]  <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[5]        <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[5] + 1 :
                                             Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[5] ;
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[5]  <=  Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[0]        <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[0] + 1 :
                                             I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[0] ;
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[0]  <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[1]        <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[1] + 1 :
                                             I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[1] ;
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[1]  <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[2]        <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[2] + 1 :
                                             I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[2] ;
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[2]  <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[3]        <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[3] + 1 :
                                             I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[3] ;
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[3]  <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[4]        <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[4] + 1 :
                                             I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[4] ;
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[4]  <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[5]        <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[5] + 1 :
                                             I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[5] ;
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[5]  <=  I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[0]        <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[0] + 1 :
                                             Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[0] ;
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[0]  <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[1]        <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[1] + 1 :
                                             Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[1] ;
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[1]  <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[2]        <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[2] + 1 :
                                             Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[2] ;
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[2]  <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[3]        <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[3] + 1 :
                                             Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[3] ;
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[3]  <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[4]        <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[4] + 1 :
                                             Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[4] ;
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[4]  <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[5]        <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[5] + 1 :
                                             Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[5] ;
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[5]  <=  Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[0]        <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[0] + 1 :
                                             I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[0] ;
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[0]  <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[1]        <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[1] + 1 :
                                             I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[1] ;
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[1]  <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[2]        <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[2] + 1 :
                                             I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[2] ;
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[2]  <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[3]        <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[3] + 1 :
                                             I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[3] ;
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[3]  <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[4]        <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[4] + 1 :
                                             I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[4] ;
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[4]  <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[5]        <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[5] + 1 :
                                             I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[5] ;
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[5]  <=  I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[0]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[0] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[0] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[0]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[1]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[1] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[1] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[1]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[2]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[2] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[2] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[2]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[3]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[3] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[3] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[3]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[4]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[4] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[4] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[4]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[5]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[5] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[5] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[5]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[6]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[6] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[6] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[6]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[7]        <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[7] + 1 :
                                             I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[7] ;
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[7]  <=  I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[0]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[0] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[0] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[0]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[1]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[1] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[1] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[1]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[2]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[2] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[2] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[2]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[3]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[3] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[3] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[3]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[4]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[4] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[4] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[4]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[5]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[5] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[5] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[5]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[6]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[6] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[6] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[6]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[7]        <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[7] + 1 :
                                             If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[7] ;
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[7]  <=  If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[0]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[0] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[0] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[0]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[1]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[1] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[1] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[1]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[2]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[2] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[2] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[2]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[3]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[3] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[3] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[3]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[4]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[4] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[4] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[4]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[5]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[5] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[5] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[5]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[6]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[6] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[6] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[6]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[7]        <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[7] + 1 :
                                             I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[7] ;
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[7]  <=  I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[0]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[0] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[0] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[0]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[1]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[1] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[1] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[1]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[2]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[2] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[2] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[2]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[3]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[3] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[3] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[3]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[4]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[4] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[4] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[4]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[5]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[5] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[5] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[5]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[6]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[6] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[6] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[6]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[7]        <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[7] + 1 :
                                             I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[7] ;
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[7]  <=  I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[0]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[0] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[0] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[0]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[1]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[1] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[1] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[1]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[2]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[2] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[2] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[2]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[3]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[3] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[3] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[3]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[4]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[4] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[4] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[4]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[5]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[5] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[5] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[5]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[6]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[6] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[6] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[6]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[7]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[7] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[7] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[7]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[8]        <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[8] + 1 :
                                             I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[8] ;
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[8]  <=  I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[0]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[0] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[0] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[0]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[1]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[1] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[1] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[1]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[2]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[2] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[2] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[2]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[3]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[3] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[3] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[3]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[4]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[4] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[4] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[4]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[5]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[5] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[5] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[5]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[6]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[6] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[6] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[6]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[7]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[7] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[7] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[7]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[8]        <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[8] + 1 :
                                             Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[8] ;
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[8]  <=  Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[0]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[0] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[0] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[0]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[1]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[1] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[1] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[1]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[2]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[2] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[2] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[2]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[3]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[3] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[3] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[3]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[4]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[4] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[4] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[4]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[5]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[5] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[5] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[5]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[6]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[6] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[6] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[6]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[7]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[7] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[7] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[7]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[8]        <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[8] + 1 :
                                             I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[8] ;
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[8]  <=  I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[0]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[0] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[0] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[0]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[1]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[1] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[1] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[1]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[2]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[2] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[2] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[2]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[3]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[3] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[3] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[3]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[4]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[4] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[4] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[4]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[5]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[5] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[5] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[5]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[6]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[6] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[6] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[6]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[7]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[7] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[7] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[7]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[8]        <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[8] + 1 :
                                             I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[8] ;
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[8]  <=  I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[0]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[0] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[0] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[0]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[1]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[1] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[1] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[1]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[2]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[2] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[2] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[2]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[3]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[3] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[3] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[3]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[4]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[4] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[4] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[4]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[5]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[5] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[5] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[5]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[6]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[6] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[6] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[6]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[7]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[7] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[7] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[7]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[8]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[8] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[8] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[8]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[9]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[9] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[9] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[9]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[10]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[10] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[10] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[10]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[11]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[11] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[11] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[11]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[12]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[12] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[12] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[12]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[13]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[13] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[13] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[13]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[14]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[14] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[14] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[14]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[15]        <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[15] + 1 :
                                             I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[15] ;
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[15]  <=  I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[0]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[0] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[0] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[0]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[1]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[1] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[1] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[1]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[2]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[2] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[2] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[2]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[3]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[3] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[3] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[3]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[4]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[4] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[4] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[4]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[5]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[5] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[5] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[5]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[6]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[6] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[6] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[6]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[7]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[7] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[7] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[7]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[8]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[8] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[8] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[8]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[9]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[9] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[9] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[9]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[10]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[10] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[10] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[10]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[11]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[11] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[11] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[11]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[12]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[12] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[12] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[12]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[13]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[13] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[13] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[13]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[14]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[14] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[14] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[14]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[15]        <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[15] + 1 :
                                             I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[15] ;
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[15]  <=  I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[0]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[0] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[0] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[0]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[1]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[1] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[1] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[1]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[2]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[2] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[2] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[2]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[3]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[3] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[3] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[3]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[4]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[4] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[4] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[4]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[5]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[5] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[5] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[5]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[6]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[6] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[6] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[6]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[7]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[7] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[7] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[7]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[8]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[8] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[8] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[8]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[9]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[9] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[9] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[9]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[10]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[10] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[10] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[10]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[11]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[11] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[11] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[11]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[12]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[12] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[12] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[12]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[13]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[13] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[13] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[13]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[14]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[14] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[14] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[14]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[15]        <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[15] + 1 :
                                             Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[15] ;
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[15]  <=  Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[0]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[0] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[0] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[0]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[1]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[1] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[1] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[1]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[2]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[2] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[2] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[2]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[3]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[3] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[3] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[3]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[4]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[4] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[4] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[4]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[5]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[5] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[5] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[5]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[6]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[6] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[6] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[6]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[7]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[7] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[7] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[7]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[8]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[8] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[8] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[8]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[9]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[9] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[9] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[9]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[10]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[10] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[10] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[10]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[11]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[11] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[11] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[11]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[12]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[12][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[12] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[12] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[12]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[12][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[13]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[13][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[13] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[13] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[13]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[13][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[14]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[14][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[14] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[14] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[14]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[14][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[15]        <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[15][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[15] + 1 :
                                             Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[15] ;
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[15]  <=  Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[15][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[0]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[0] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[0] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[0]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[1]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[1] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[1] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[1]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[2]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[2] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[2] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[2]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[3]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[3] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[3] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[3]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[4]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[4] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[4] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[4]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[5]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[5] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[5] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[5]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[6]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[6] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[6] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[6]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[7]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[7] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[7] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[7]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[8]        <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[8] + 1 :
                                             I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[8] ;
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[8]  <=  I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[0]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[0] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[0] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[0]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[1]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[1] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[1] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[1]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[2]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[2] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[2] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[2]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[3]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[3] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[3] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[3]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[4]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[4] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[4] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[4]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[5]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[5] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[5] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[5]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[6]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[6] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[6] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[6]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[7]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[7] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[7] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[7]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[8]        <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[8] + 1 :
                                             Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[8] ;
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[8]  <=  Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[0]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[0] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[0] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[0]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[1]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[1] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[1] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[1]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[2]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[2] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[2] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[2]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[3]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[3] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[3] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[3]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[4]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[4] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[4] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[4]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[5]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[5] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[5] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[5]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[6]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[6] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[6] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[6]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[7]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[7] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[7] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[7]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[8]        <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[8] + 1 :
                                             I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[8] ;
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[8]  <=  I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[0]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[0] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[0] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[0]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[1]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[1] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[1] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[1]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[2]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[2] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[2] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[2]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[3]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[3] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[3] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[3]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[4]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[4] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[4] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[4]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[5]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[5] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[5] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[5]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[6]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[6] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[6] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[6]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[7]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[7] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[7] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[7]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[8]        <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[8] + 1 :
                                             Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[8] ;
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[8]  <=  Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[0]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[0] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[0] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[0]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[1]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[1] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[1] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[1]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[2]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[2] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[2] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[2]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[3]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[3] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[3] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[3]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[4]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[4] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[4] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[4]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[5]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[5] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[5] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[5]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[6]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[6] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[6] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[6]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[7]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[7] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[7] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[7]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[8]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[8] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[8] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[8]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[9]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[9] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[9] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[9]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[10]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[10] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[10] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[10]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[11]        <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[11] + 1 :
                                             I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[11] ;
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[11]  <=  I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[0]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[0] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[0] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[0]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[1]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[1] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[1] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[1]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[2]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[2] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[2] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[2]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[3]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[3] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[3] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[3]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[4]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[4] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[4] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[4]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[5]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[5] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[5] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[5]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[6]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[6] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[6] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[6]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[7]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[7] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[7] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[7]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[8]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[8] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[8] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[8]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[9]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[9] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[9] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[9]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[10]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[10] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[10] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[10]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[11]        <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[11] + 1 :
                                             Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[11] ;
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[11]  <=  Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[0]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[0] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[0] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[0]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[1]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[1] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[1] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[1]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[2]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[2] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[2] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[2]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[3]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[3] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[3] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[3]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[4]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[4] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[4] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[4]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[5]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[5] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[5] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[5]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[6]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[6] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[6] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[6]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[7]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[7] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[7] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[7]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[8]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[8] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[8] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[8]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[9]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[9] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[9] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[9]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[10]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[10] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[10] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[10]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[11]        <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[11] + 1 :
                                             Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[11] ;
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[11]  <=  Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[0]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[0] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[0] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[0]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[1]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[1][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[1] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[1] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[1]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[1][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[2]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[2][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[2] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[2] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[2]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[2][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[3]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[3][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[3] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[3] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[3]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[3][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[4]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[4][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[4] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[4] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[4]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[4][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[5]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[5][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[5] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[5] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[5]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[5][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[6]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[6][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[6] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[6] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[6]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[6][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[7]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[7][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[7] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[7] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[7]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[7][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[8]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[8][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[8] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[8] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[8]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[8][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[9]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[9][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[9] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[9] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[9]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[9][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[10]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[10][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[10] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[10] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[10]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[10][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[11]        <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[11][MAX_SUM_WDTH_LONG-1] ?
                                             ~I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[11] + 1 :
                                             I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[11] ;
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[11]  <=  I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[11][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9aea0703810e5cd52352d3b0ede17aa0ccb943f1e0507585e4cccd0d0c427e98[0]        <=  Ida88a2dbb8109dff5f061f3ecaf9586a219f6355e92312ffd580a09126c72376[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ida88a2dbb8109dff5f061f3ecaf9586a219f6355e92312ffd580a09126c72376[0] + 1 :
                                             Ida88a2dbb8109dff5f061f3ecaf9586a219f6355e92312ffd580a09126c72376[0] ;
            Iea53e5522afe762dd4185f0262512abbb94b905893974c13e954df5553942b1d[0]  <=  Ida88a2dbb8109dff5f061f3ecaf9586a219f6355e92312ffd580a09126c72376[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I42c6c1d7cfb81335f01807b1d1c6b77c109482d338e81eda1ed174f739a6bf1b[0]        <=  I73f2fe34b7ee9a375ae43b6d3cbd515175de303a77f64ad277094e9bb8e45177[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I73f2fe34b7ee9a375ae43b6d3cbd515175de303a77f64ad277094e9bb8e45177[0] + 1 :
                                             I73f2fe34b7ee9a375ae43b6d3cbd515175de303a77f64ad277094e9bb8e45177[0] ;
            If481e9fd41cf8181d432f397381b8376d9da7ddfba17b52e65e301e74c3b9b0d[0]  <=  I73f2fe34b7ee9a375ae43b6d3cbd515175de303a77f64ad277094e9bb8e45177[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I839de42c6f3369ef5c6200c12baee8c9e698b3108fd6dcd58a71351d9bedae54[0]        <=  I9f9254e3af43fc1c116a2d33bee39fb18594b7696e59d5aa4c3884363616a5d6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9f9254e3af43fc1c116a2d33bee39fb18594b7696e59d5aa4c3884363616a5d6[0] + 1 :
                                             I9f9254e3af43fc1c116a2d33bee39fb18594b7696e59d5aa4c3884363616a5d6[0] ;
            If2e4ac195be838db9dd7b062319aba299887896862f1a340013226fa025b18fc[0]  <=  I9f9254e3af43fc1c116a2d33bee39fb18594b7696e59d5aa4c3884363616a5d6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0a1e88a592eeec68c060dd84ca2d75809b8fd80dd97a01a8d12cd9869bf94532[0]        <=  Idbd45e6a4aa2cf66d740fb7d3c41c5d4af78bdfe13d321e6ee7eceb153e03de4[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idbd45e6a4aa2cf66d740fb7d3c41c5d4af78bdfe13d321e6ee7eceb153e03de4[0] + 1 :
                                             Idbd45e6a4aa2cf66d740fb7d3c41c5d4af78bdfe13d321e6ee7eceb153e03de4[0] ;
            I40914301545dfe0b6673f76e0dc0d1ab3968ca3b18fe8f4ff63d5623c31bafa7[0]  <=  Idbd45e6a4aa2cf66d740fb7d3c41c5d4af78bdfe13d321e6ee7eceb153e03de4[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9114e17d37b4346674c23a6ef3a2aee35426292fbf73d7f30c895090bb749034[0]        <=  Ie3a6f677abff075b84cd72fb72f4b4ad16dc2a915b2d3e06d8136c5073549499[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie3a6f677abff075b84cd72fb72f4b4ad16dc2a915b2d3e06d8136c5073549499[0] + 1 :
                                             Ie3a6f677abff075b84cd72fb72f4b4ad16dc2a915b2d3e06d8136c5073549499[0] ;
            Idf30e1a70a723113d32f621f0375dd85270da2f7386cff5ef4ff88cfca78b848[0]  <=  Ie3a6f677abff075b84cd72fb72f4b4ad16dc2a915b2d3e06d8136c5073549499[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ife5225eb20e50e3cc959d9080f6faa318b4977bc9d04a67414a6cdf16c98e295[0]        <=  I6444b0cde8c0fcb1cc0b51c11d3937bd156b26f21a0eca3cabe0c6b0e696f7c0[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6444b0cde8c0fcb1cc0b51c11d3937bd156b26f21a0eca3cabe0c6b0e696f7c0[0] + 1 :
                                             I6444b0cde8c0fcb1cc0b51c11d3937bd156b26f21a0eca3cabe0c6b0e696f7c0[0] ;
            Ic246bc24fb918b7c4a32727a332df57bfb205adc05150ae8d944a77cbdc62822[0]  <=  I6444b0cde8c0fcb1cc0b51c11d3937bd156b26f21a0eca3cabe0c6b0e696f7c0[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I28dfde2c443cd84194231fc87b8a1c6382ff3c2ff9b6d43e31e3a7116be41169[0]        <=  I1d41ad001c01e3dc84cd02ab5ba24e8239e273f81dad37de1fdf873305e073c3[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I1d41ad001c01e3dc84cd02ab5ba24e8239e273f81dad37de1fdf873305e073c3[0] + 1 :
                                             I1d41ad001c01e3dc84cd02ab5ba24e8239e273f81dad37de1fdf873305e073c3[0] ;
            I6cac9957a16e7cfa8a125b40d8ce42cb7f502078a791b177d9bbe9589b612426[0]  <=  I1d41ad001c01e3dc84cd02ab5ba24e8239e273f81dad37de1fdf873305e073c3[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I55da00c15261d3abb33c69ecc3f2090fb2bb3c29a3653fd999f6232982cf31ac[0]        <=  I75cef0e0547fa056ba6e20b68cadef6bea875e9b12fe99c286e8d79a40c9043f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I75cef0e0547fa056ba6e20b68cadef6bea875e9b12fe99c286e8d79a40c9043f[0] + 1 :
                                             I75cef0e0547fa056ba6e20b68cadef6bea875e9b12fe99c286e8d79a40c9043f[0] ;
            Iee4ad1e7709a56d53cd8b97f587f1f791fb88bf278fcfef32a29fa05247ca13d[0]  <=  I75cef0e0547fa056ba6e20b68cadef6bea875e9b12fe99c286e8d79a40c9043f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I05ca033870ef7adc8ce911a962bbd120591a1fe3b3044782b7e569e2b94ac629[0]        <=  Ie4bd6fa32fac971db980d5dae63887ea1f4b75f375f1953975e4ead5b727d37a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie4bd6fa32fac971db980d5dae63887ea1f4b75f375f1953975e4ead5b727d37a[0] + 1 :
                                             Ie4bd6fa32fac971db980d5dae63887ea1f4b75f375f1953975e4ead5b727d37a[0] ;
            I16a4499c48e5c24fd8a6d49ec3bf63c20c85f440c0c897cdb840e9f28fa2e68a[0]  <=  Ie4bd6fa32fac971db980d5dae63887ea1f4b75f375f1953975e4ead5b727d37a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4ef4ed6e15f48f289815b7e00b2454a26e076b8dc9b8903e118507c9688e905d[0]        <=  I40f5e53051d38a2da1e0c992989c7740e6a7be23273e1412d01e853851b97a0b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I40f5e53051d38a2da1e0c992989c7740e6a7be23273e1412d01e853851b97a0b[0] + 1 :
                                             I40f5e53051d38a2da1e0c992989c7740e6a7be23273e1412d01e853851b97a0b[0] ;
            Ibed209db0bc502e3fceb4ab86ac20a2ebf87c43391a546d592e5aa32709aa8bd[0]  <=  I40f5e53051d38a2da1e0c992989c7740e6a7be23273e1412d01e853851b97a0b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I25e57b538f9a08a355a5ff8d26d94f81bbf2ebd0039881e74aec76ffb1dd48aa[0]        <=  I0e9c027df8259f9e499658f9ee700b50ea04b829312da04e92f13edd2af302ad[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I0e9c027df8259f9e499658f9ee700b50ea04b829312da04e92f13edd2af302ad[0] + 1 :
                                             I0e9c027df8259f9e499658f9ee700b50ea04b829312da04e92f13edd2af302ad[0] ;
            I05dc9e8db597a2123632b2934d864ae64cab5192401d8f66ebebd95618590ba2[0]  <=  I0e9c027df8259f9e499658f9ee700b50ea04b829312da04e92f13edd2af302ad[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I070ee6bd21603d58d3243ac556db2ca3c0476c64fde6d32aff54e0577b0472f0[0]        <=  If5d8bf4cfab249bae208cb278b5fc90873cebd7a677b1d1e22df49b576863146[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If5d8bf4cfab249bae208cb278b5fc90873cebd7a677b1d1e22df49b576863146[0] + 1 :
                                             If5d8bf4cfab249bae208cb278b5fc90873cebd7a677b1d1e22df49b576863146[0] ;
            Ib309786164a7d646c17533008b3aaf0fd86eda3c5ee167efc2080ef5b26a9ddf[0]  <=  If5d8bf4cfab249bae208cb278b5fc90873cebd7a677b1d1e22df49b576863146[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id2ede5f3d3ce0652bc9ceeadf1de91fb99234718893eea8cc1779cf900284e88[0]        <=  I03501709a4343537388784e4e39cb9c1b52beb3749d09e2daaf1910dc5b1e2b2[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I03501709a4343537388784e4e39cb9c1b52beb3749d09e2daaf1910dc5b1e2b2[0] + 1 :
                                             I03501709a4343537388784e4e39cb9c1b52beb3749d09e2daaf1910dc5b1e2b2[0] ;
            Id9bbd0f5c16ba0ffae6a0e5304e1726b97df06f06feaccbb1bbcaf0e01be3823[0]  <=  I03501709a4343537388784e4e39cb9c1b52beb3749d09e2daaf1910dc5b1e2b2[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie251294e2cb883a913e91485cecfa90bbd107955ceb6d60d4a9b1808aaadb2d4[0]        <=  I46aa1767826fecc6fede490a807238d69235f3cdf96dc753215e008a12454119[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I46aa1767826fecc6fede490a807238d69235f3cdf96dc753215e008a12454119[0] + 1 :
                                             I46aa1767826fecc6fede490a807238d69235f3cdf96dc753215e008a12454119[0] ;
            I4294b001f220e009c2a65fbf8b36ce1d8961c317ae8ded31cbe5aa288191e009[0]  <=  I46aa1767826fecc6fede490a807238d69235f3cdf96dc753215e008a12454119[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I983e8c64c323025590663edf53b0666d93d838f15879b5e3df245a8e9ac6fb80[0]        <=  Id749da645d127d8ff383558a6e7ab4a5c2a59f513cb7808fa4dc4e9f6f14f2b9[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id749da645d127d8ff383558a6e7ab4a5c2a59f513cb7808fa4dc4e9f6f14f2b9[0] + 1 :
                                             Id749da645d127d8ff383558a6e7ab4a5c2a59f513cb7808fa4dc4e9f6f14f2b9[0] ;
            Id1fe66d1340965020f513e73a4f77d18f4703c194c3954d40a7f1bc37fc1342b[0]  <=  Id749da645d127d8ff383558a6e7ab4a5c2a59f513cb7808fa4dc4e9f6f14f2b9[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46e5ca785f6f4304dbc4fbbf3816d83106047f0eceea77717a1ad5c41a9ca441[0]        <=  Ib15e62b641f64f20a1d3baff39f2dc6a403616e09955f5d7f47ba4fc093badc9[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib15e62b641f64f20a1d3baff39f2dc6a403616e09955f5d7f47ba4fc093badc9[0] + 1 :
                                             Ib15e62b641f64f20a1d3baff39f2dc6a403616e09955f5d7f47ba4fc093badc9[0] ;
            Ie95c9af987f352eca30c8546d306af7cdada8d2a8037200d303e6afbd5a4f448[0]  <=  Ib15e62b641f64f20a1d3baff39f2dc6a403616e09955f5d7f47ba4fc093badc9[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ibefeb67be2754ad6b9a6cda09c66529a7ca51536f5c6ca6b05e6ac1de34ae514[0]        <=  I603d7bbab10dd31f19047e4a73046c804506ba70d1504351984be41bae1d180e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I603d7bbab10dd31f19047e4a73046c804506ba70d1504351984be41bae1d180e[0] + 1 :
                                             I603d7bbab10dd31f19047e4a73046c804506ba70d1504351984be41bae1d180e[0] ;
            Id34d005cdd89bf304f95101c6fbfdd40d6c0b1742b5f3bee3bf043bf88c3d063[0]  <=  I603d7bbab10dd31f19047e4a73046c804506ba70d1504351984be41bae1d180e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0dd45b65c82498edff9ac44b5b07ed30818dc1ea2af48e5c1394466865f36adf[0]        <=  Ia7b80ae8cf2697315846253262614611c079c53ada59bf7d982596ff8df770b6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia7b80ae8cf2697315846253262614611c079c53ada59bf7d982596ff8df770b6[0] + 1 :
                                             Ia7b80ae8cf2697315846253262614611c079c53ada59bf7d982596ff8df770b6[0] ;
            I79d61ad4114817a49b1dc8e9314d9e3be9758d861974ead362ff0ac862d1d77f[0]  <=  Ia7b80ae8cf2697315846253262614611c079c53ada59bf7d982596ff8df770b6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ica92be8c7303e09b9f549ec558e655816c1d23a39b8d5324060f64a391984c1b[0]        <=  I58250efea716c203d1475c4046ca67a47a156f9e4709d26d4b05a29ed1578337[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I58250efea716c203d1475c4046ca67a47a156f9e4709d26d4b05a29ed1578337[0] + 1 :
                                             I58250efea716c203d1475c4046ca67a47a156f9e4709d26d4b05a29ed1578337[0] ;
            Icfe1fffea36cf64044389903be9550fe283d4dbb7f1b47aff2005e70765a6045[0]  <=  I58250efea716c203d1475c4046ca67a47a156f9e4709d26d4b05a29ed1578337[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I726b6a7ed2ab76b049762263a08d5121a597f30ce25a6880b51d6b01aff801d7[0]        <=  I50cccb280c7d65372645e94b4a4d472860f246a8a6d89c02e4feee7dac903e8e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I50cccb280c7d65372645e94b4a4d472860f246a8a6d89c02e4feee7dac903e8e[0] + 1 :
                                             I50cccb280c7d65372645e94b4a4d472860f246a8a6d89c02e4feee7dac903e8e[0] ;
            Ib08cf17b2065d04f587d1a8231ec1e4bbb6b2b15819de8a7efe18b477515ccf8[0]  <=  I50cccb280c7d65372645e94b4a4d472860f246a8a6d89c02e4feee7dac903e8e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I89362accf0644c192f06b113020d2071f1389e8ddd8d4fee492205db15b25b66[0]        <=  I01d4a1a1123a68c80a967604072ca420c79d4e205c354221591cdbcaa24c4050[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I01d4a1a1123a68c80a967604072ca420c79d4e205c354221591cdbcaa24c4050[0] + 1 :
                                             I01d4a1a1123a68c80a967604072ca420c79d4e205c354221591cdbcaa24c4050[0] ;
            I21832b7270210e1bb6a23930ad9ced36d3da201d80310263e26eb96bebd23612[0]  <=  I01d4a1a1123a68c80a967604072ca420c79d4e205c354221591cdbcaa24c4050[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4473c0cfd2d569bc671ba814a524058946271eb49a04fc384e9373185e1f4a6b[0]        <=  I702778e2f8308e720ae6aebd003938631b4a76341308834c90d10eeb3611ce3f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I702778e2f8308e720ae6aebd003938631b4a76341308834c90d10eeb3611ce3f[0] + 1 :
                                             I702778e2f8308e720ae6aebd003938631b4a76341308834c90d10eeb3611ce3f[0] ;
            I5dcc76c47f3c9129431152fa6f7047be203fc556198b45db15a9991647bb8c85[0]  <=  I702778e2f8308e720ae6aebd003938631b4a76341308834c90d10eeb3611ce3f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2ba73f603d9cb767572f2b2f2a9732e2ebc066392aa85888df87da4dd8b84113[0]        <=  Id2ba36bb60a1673c62e790e5ad15a4fdd49bc397b3cba8e6251a88e63c249091[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id2ba36bb60a1673c62e790e5ad15a4fdd49bc397b3cba8e6251a88e63c249091[0] + 1 :
                                             Id2ba36bb60a1673c62e790e5ad15a4fdd49bc397b3cba8e6251a88e63c249091[0] ;
            I450f5b0f5d2b96636ae010048040ebd744fc4ca164cd764bb33615741ecaa62f[0]  <=  Id2ba36bb60a1673c62e790e5ad15a4fdd49bc397b3cba8e6251a88e63c249091[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I82f10eef14d4ad82b1f7f8c5d056c398386a6cf790095113a615a8bb6cfba233[0]        <=  Ifb22aa4df653a2afecbf1dc570c526ccf003e19a0f5972b9bc5ba9458e316ba6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifb22aa4df653a2afecbf1dc570c526ccf003e19a0f5972b9bc5ba9458e316ba6[0] + 1 :
                                             Ifb22aa4df653a2afecbf1dc570c526ccf003e19a0f5972b9bc5ba9458e316ba6[0] ;
            I35d64df6881fde0d4836aa408258db7cc1bfb2f066abf8c9345670b78c466b9e[0]  <=  Ifb22aa4df653a2afecbf1dc570c526ccf003e19a0f5972b9bc5ba9458e316ba6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2fd5dd69a5f551c26d9970d09ab0e26ac5183a0022af58e2bec1dd1efefb139c[0]        <=  I43fb6b8f15f49b741ef111f2b4a57e5da84af4d6f3ce9b92e0a2bedb18eef4bf[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I43fb6b8f15f49b741ef111f2b4a57e5da84af4d6f3ce9b92e0a2bedb18eef4bf[0] + 1 :
                                             I43fb6b8f15f49b741ef111f2b4a57e5da84af4d6f3ce9b92e0a2bedb18eef4bf[0] ;
            I11944fb91fa1b1d5f076cc36db77f0f8434f0edbb1236c7a9bcb45f79432ea9f[0]  <=  I43fb6b8f15f49b741ef111f2b4a57e5da84af4d6f3ce9b92e0a2bedb18eef4bf[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2fd258374a5bda5c58c1fdc6e305789a598fbe70657d6dc18e8878b6c2b0441a[0]        <=  Ibc1b6326c8e2b05aef237f6ded855eb730c445a3cb6c7d49293ef68b6ec623ea[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibc1b6326c8e2b05aef237f6ded855eb730c445a3cb6c7d49293ef68b6ec623ea[0] + 1 :
                                             Ibc1b6326c8e2b05aef237f6ded855eb730c445a3cb6c7d49293ef68b6ec623ea[0] ;
            I49642204473312df5a3bcab2692aa7558f44f21416226675a4ec10b0543cc5e9[0]  <=  Ibc1b6326c8e2b05aef237f6ded855eb730c445a3cb6c7d49293ef68b6ec623ea[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I76942d3b012aef2097112a1c1adfa2bf986414df19a633b87d2f3c2a61d27351[0]        <=  I3a8bec62f5e0501c90baaa2f6f7288929d91d107a2197e1c574428638cd020d7[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I3a8bec62f5e0501c90baaa2f6f7288929d91d107a2197e1c574428638cd020d7[0] + 1 :
                                             I3a8bec62f5e0501c90baaa2f6f7288929d91d107a2197e1c574428638cd020d7[0] ;
            I24e0d361a2679430549932a968d7cc25f980275fea5554e3453ed0a652d31caa[0]  <=  I3a8bec62f5e0501c90baaa2f6f7288929d91d107a2197e1c574428638cd020d7[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ida428d199205588ecd8cc963ceb39e24bf6f2d004b675f3cb883960e0f089842[0]        <=  Ie8930f54b7806297e3bb1082b70d74d5eaeaf269112a0d5f82caf5c941ff7a2b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie8930f54b7806297e3bb1082b70d74d5eaeaf269112a0d5f82caf5c941ff7a2b[0] + 1 :
                                             Ie8930f54b7806297e3bb1082b70d74d5eaeaf269112a0d5f82caf5c941ff7a2b[0] ;
            I386015f8daacd2ac9cfed376d3418b56ac13f075a43dde939e4056c29565a926[0]  <=  Ie8930f54b7806297e3bb1082b70d74d5eaeaf269112a0d5f82caf5c941ff7a2b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I91f0247d07693c53d716345c810ffa0ee8d3f4b793ca8831763f5465db649c89[0]        <=  I948dbc4fe20518395aaa5356bb504e41a80332a8adbba9ae4c6d8a4ca0704b7b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I948dbc4fe20518395aaa5356bb504e41a80332a8adbba9ae4c6d8a4ca0704b7b[0] + 1 :
                                             I948dbc4fe20518395aaa5356bb504e41a80332a8adbba9ae4c6d8a4ca0704b7b[0] ;
            I32832b039ae7e6f4b1e38cfdf680e5044e383b921a76189054511ebe5b8c0d7c[0]  <=  I948dbc4fe20518395aaa5356bb504e41a80332a8adbba9ae4c6d8a4ca0704b7b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I754c4c2dda64bb938ac60db8cd469c6f3ee0831a3a6b6b98e902c1b72663ff28[0]        <=  I5140e483e7397c66b8d4835ac2e465f125e62c4feb9835d7a5f5ea7849def4dc[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5140e483e7397c66b8d4835ac2e465f125e62c4feb9835d7a5f5ea7849def4dc[0] + 1 :
                                             I5140e483e7397c66b8d4835ac2e465f125e62c4feb9835d7a5f5ea7849def4dc[0] ;
            I09fff9b84a38f3d19685f9627d01a7183cf65d72110802f11e8da0e01194bf88[0]  <=  I5140e483e7397c66b8d4835ac2e465f125e62c4feb9835d7a5f5ea7849def4dc[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I567c2801d5598a057d5773ea5045f594de038bab88d554ad2c713cf56ef632b4[0]        <=  If049a08cd46a811753b3637ee0a96207144b0a5eade57068ba5712c3ba23c8ae[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If049a08cd46a811753b3637ee0a96207144b0a5eade57068ba5712c3ba23c8ae[0] + 1 :
                                             If049a08cd46a811753b3637ee0a96207144b0a5eade57068ba5712c3ba23c8ae[0] ;
            Ib82c65f09934744abbba984b6e375bd69ce7231a5085bb00ba4e673cfd3aba38[0]  <=  If049a08cd46a811753b3637ee0a96207144b0a5eade57068ba5712c3ba23c8ae[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic9f57a4a1184139b219a3a5e3c554705469b79d3ab175ddc74512ccbfd5898b0[0]        <=  I6b404c4caf16f09360a848f09b33c16a69029ab05067f1bca94eba5e69701d37[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6b404c4caf16f09360a848f09b33c16a69029ab05067f1bca94eba5e69701d37[0] + 1 :
                                             I6b404c4caf16f09360a848f09b33c16a69029ab05067f1bca94eba5e69701d37[0] ;
            I8ec5727130bf67c04580aa1b5b46cdf964db65750f2fc9ce55025b1c117b2bef[0]  <=  I6b404c4caf16f09360a848f09b33c16a69029ab05067f1bca94eba5e69701d37[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2dc38e534505cf47f391eb9f4b090e16136d12619b4fe91cc8029bb5a050689d[0]        <=  I1efde896c2d2e97d2b635b34d6ad30d31a8c855ea5975dfadcf5ea136fa3d063[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I1efde896c2d2e97d2b635b34d6ad30d31a8c855ea5975dfadcf5ea136fa3d063[0] + 1 :
                                             I1efde896c2d2e97d2b635b34d6ad30d31a8c855ea5975dfadcf5ea136fa3d063[0] ;
            I862dddc300df692e8bbf4ca45a24d840e51ac1e975631cf4ebb8337ceefc2eb1[0]  <=  I1efde896c2d2e97d2b635b34d6ad30d31a8c855ea5975dfadcf5ea136fa3d063[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib83aabc196c7633dfb4a9bcb4b8d06959130620de297f9dff77b1454a8f2f96d[0]        <=  I860fff7ccba78c970b447509ccd6de21b521bd8458673134640ce16c6f1ead4e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I860fff7ccba78c970b447509ccd6de21b521bd8458673134640ce16c6f1ead4e[0] + 1 :
                                             I860fff7ccba78c970b447509ccd6de21b521bd8458673134640ce16c6f1ead4e[0] ;
            Id08a37df0c5095196e2d760938c4d0b7e8716c25b55d9a9656d86c2c473f9c2f[0]  <=  I860fff7ccba78c970b447509ccd6de21b521bd8458673134640ce16c6f1ead4e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia23743e423f143b75923bc7b1a4363323d46ace080c8ee9d15ff687afd4bef65[0]        <=  I9786358e2588e06550a490e47029ce233b6d39273ad261316c5f730a7ee4bf17[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9786358e2588e06550a490e47029ce233b6d39273ad261316c5f730a7ee4bf17[0] + 1 :
                                             I9786358e2588e06550a490e47029ce233b6d39273ad261316c5f730a7ee4bf17[0] ;
            I40204cd18eb803f82fc3ef933553c6ec41331f6d4a15538c287b8f57adebb89e[0]  <=  I9786358e2588e06550a490e47029ce233b6d39273ad261316c5f730a7ee4bf17[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id49eabe82a09acf1b3a3aa3be9bfbc0ff958b96b44ada842e892c587fbddb8fc[0]        <=  Ia01e9ec22c644f28b2be05c8002d4f576e816688e30965ae9f3ef78ca1272b9b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia01e9ec22c644f28b2be05c8002d4f576e816688e30965ae9f3ef78ca1272b9b[0] + 1 :
                                             Ia01e9ec22c644f28b2be05c8002d4f576e816688e30965ae9f3ef78ca1272b9b[0] ;
            I677f733f4e801d99dc2fd1987683a7ac6c8609d84da6c95b8a7056ce07845665[0]  <=  Ia01e9ec22c644f28b2be05c8002d4f576e816688e30965ae9f3ef78ca1272b9b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I93584fe5ab7128b24b2372bfeea00f7a2bf09d50b1fb535d01cc141c6d6fc377[0]        <=  I0797e7fab1998d109cd09e4aa801cd2dfe57364a83e9c84bef81be8f59ca729e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I0797e7fab1998d109cd09e4aa801cd2dfe57364a83e9c84bef81be8f59ca729e[0] + 1 :
                                             I0797e7fab1998d109cd09e4aa801cd2dfe57364a83e9c84bef81be8f59ca729e[0] ;
            Ifeb10787a88bae5943b616e3bf751faff5e7eea80e45e24d60a760f4d6b0154c[0]  <=  I0797e7fab1998d109cd09e4aa801cd2dfe57364a83e9c84bef81be8f59ca729e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I44142c70d3ba4660f5b85d895710afc623ed3470ba85eab3dee5e49a59e1b124[0]        <=  I035ba5b524312fb6136ca853695154f9334f6336e5acf5884beebeff72197c7d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I035ba5b524312fb6136ca853695154f9334f6336e5acf5884beebeff72197c7d[0] + 1 :
                                             I035ba5b524312fb6136ca853695154f9334f6336e5acf5884beebeff72197c7d[0] ;
            Iecc97eedc286cd1c3d301e35036e81a10d164d59da9252a92ca5f355a828367b[0]  <=  I035ba5b524312fb6136ca853695154f9334f6336e5acf5884beebeff72197c7d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id8b538e6a6c4a147c7000388923f1d89a193f8ec53ef214556e005218d2c240e[0]        <=  If058a896104351e61394ece6dde5212381937b7d36a4b63f5e99a268d5c7722b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If058a896104351e61394ece6dde5212381937b7d36a4b63f5e99a268d5c7722b[0] + 1 :
                                             If058a896104351e61394ece6dde5212381937b7d36a4b63f5e99a268d5c7722b[0] ;
            Ia9a21e6f22a6cc828e041980ab142b418938a92bf8e868216402a46b8c614a19[0]  <=  If058a896104351e61394ece6dde5212381937b7d36a4b63f5e99a268d5c7722b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I658f9399a929745b4ba467a1e019fdbe214acd543dd4f5f51a95292420281401[0]        <=  I29e36792da89f6ea79232a191af837f9da3739332265e00d97d40b09ef384a58[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I29e36792da89f6ea79232a191af837f9da3739332265e00d97d40b09ef384a58[0] + 1 :
                                             I29e36792da89f6ea79232a191af837f9da3739332265e00d97d40b09ef384a58[0] ;
            I355f4f82732333ae56692d1c7ee89b368d938d9ce1d5f806be7e46482c10e19c[0]  <=  I29e36792da89f6ea79232a191af837f9da3739332265e00d97d40b09ef384a58[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id1ba70174cf019078c719d1d50a82a61fbfdeea2a13e21a1247e567b9266365f[0]        <=  I5e9d25157a8f35aed3b702ea5120ad81de73bafda0cb5811bae0fd0eaf2d11e1[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5e9d25157a8f35aed3b702ea5120ad81de73bafda0cb5811bae0fd0eaf2d11e1[0] + 1 :
                                             I5e9d25157a8f35aed3b702ea5120ad81de73bafda0cb5811bae0fd0eaf2d11e1[0] ;
            I9b2ce64b97ca55921bacb9b6aa4cdc8da5c1e33db4215a2470b7cfab3693576c[0]  <=  I5e9d25157a8f35aed3b702ea5120ad81de73bafda0cb5811bae0fd0eaf2d11e1[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I797dfd66b521bd680024b6e46455d624aa58b4271f5e6ca19fc7abf520f26222[0]        <=  I57f4038fbe1f52bf47fe1cdbb52088b800609231fa2007cb1ff941817005a0ce[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I57f4038fbe1f52bf47fe1cdbb52088b800609231fa2007cb1ff941817005a0ce[0] + 1 :
                                             I57f4038fbe1f52bf47fe1cdbb52088b800609231fa2007cb1ff941817005a0ce[0] ;
            I2d78ac4a4125ec25a02df6484c0ae640a37f915383b72f33b91e87cdf376fdf7[0]  <=  I57f4038fbe1f52bf47fe1cdbb52088b800609231fa2007cb1ff941817005a0ce[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I74f49d84817f2467b8ccdf03acbd7372c58f1a4fddcce45cb882431b2be20b39[0]        <=  I592de5159deb6cf98840aff691c78457fefe7ee33d85506cd1dd400679207812[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I592de5159deb6cf98840aff691c78457fefe7ee33d85506cd1dd400679207812[0] + 1 :
                                             I592de5159deb6cf98840aff691c78457fefe7ee33d85506cd1dd400679207812[0] ;
            Id727bdc545af53e8f89be0ac5627d0c0c0f0bd7d75030bcb41f198a4fe9c7d64[0]  <=  I592de5159deb6cf98840aff691c78457fefe7ee33d85506cd1dd400679207812[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib756dd9d8d9a5233fcd368ffa91f5d7d9c8825b01bc26140e5a717d3ce263e64[0]        <=  I262ef0e0ef60c8effdcfb37ad79058672a12fe1aa6b0099d00f1067fb709c255[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I262ef0e0ef60c8effdcfb37ad79058672a12fe1aa6b0099d00f1067fb709c255[0] + 1 :
                                             I262ef0e0ef60c8effdcfb37ad79058672a12fe1aa6b0099d00f1067fb709c255[0] ;
            I7661c17a1c73dbca82a6d3bfba2ab85ebb0131c1e513f093e1b0aec54907595d[0]  <=  I262ef0e0ef60c8effdcfb37ad79058672a12fe1aa6b0099d00f1067fb709c255[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I1bb2be29dd44258b24a36ad9b1625ead1cf965856f1d9695c62ae80de142169d[0]        <=  Ic69f5c16ae27a74a97e7bc6fce24e0c868c1e1e5b6a348410853d40bb11f5d91[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic69f5c16ae27a74a97e7bc6fce24e0c868c1e1e5b6a348410853d40bb11f5d91[0] + 1 :
                                             Ic69f5c16ae27a74a97e7bc6fce24e0c868c1e1e5b6a348410853d40bb11f5d91[0] ;
            I553a83634252c50164bdde3576d7e1552a147490d02eac6dfd1140a46b813d08[0]  <=  Ic69f5c16ae27a74a97e7bc6fce24e0c868c1e1e5b6a348410853d40bb11f5d91[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icbff209e6c8353c58f46c0688f06da0cdf71a95defd8937f2d52d63d387d74b5[0]        <=  I0bba5d4133f73c77eb3812cb20554c368cfe3a6ddc34cc7405b33921fbbd9a2a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I0bba5d4133f73c77eb3812cb20554c368cfe3a6ddc34cc7405b33921fbbd9a2a[0] + 1 :
                                             I0bba5d4133f73c77eb3812cb20554c368cfe3a6ddc34cc7405b33921fbbd9a2a[0] ;
            Ib450c1ee41d04516060a410bbdfb605f0ce13cd8781596ce5218928ed207de8a[0]  <=  I0bba5d4133f73c77eb3812cb20554c368cfe3a6ddc34cc7405b33921fbbd9a2a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia628bc749f04b3d12509effbd4e0bc5ac0fadf48a2cd5663e4c2094593870a42[0]        <=  I98234b1225d9d3d636129139d51ebd098c46162cd51cf3530b9c8f8c0f12684c[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I98234b1225d9d3d636129139d51ebd098c46162cd51cf3530b9c8f8c0f12684c[0] + 1 :
                                             I98234b1225d9d3d636129139d51ebd098c46162cd51cf3530b9c8f8c0f12684c[0] ;
            Ica745abd4de790f1cd3e2a5a32a9d0b5edf1b64e85759c49f3b4e51779443709[0]  <=  I98234b1225d9d3d636129139d51ebd098c46162cd51cf3530b9c8f8c0f12684c[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5ac2c7b61022af9bd2550f824b8e129ca1c336b1ff900b0af785d86e33cf3358[0]        <=  I31906081d1cabbb8c066a2d5377802f2366fe4f3993b4f749f59d89ed1fe0388[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I31906081d1cabbb8c066a2d5377802f2366fe4f3993b4f749f59d89ed1fe0388[0] + 1 :
                                             I31906081d1cabbb8c066a2d5377802f2366fe4f3993b4f749f59d89ed1fe0388[0] ;
            I6399b29558311ea40cda1388848ce13bb7593bfed01ca2a10fa5d8ed6700df56[0]  <=  I31906081d1cabbb8c066a2d5377802f2366fe4f3993b4f749f59d89ed1fe0388[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie511320217185f90f1e4a23ab51ae9686801b09657c714a5bdd9c4e26f070bff[0]        <=  I735b667ac51f343a3a50cbaf5478e1095cf20f38a650d24285dbb38ba66abbbd[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I735b667ac51f343a3a50cbaf5478e1095cf20f38a650d24285dbb38ba66abbbd[0] + 1 :
                                             I735b667ac51f343a3a50cbaf5478e1095cf20f38a650d24285dbb38ba66abbbd[0] ;
            I6f529a4dd77f75d9af4350baf53ba61c1e9c5ea6227c26690987d244dfe71528[0]  <=  I735b667ac51f343a3a50cbaf5478e1095cf20f38a650d24285dbb38ba66abbbd[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I032b833c683eaf0c1c4c60ad831278ab0ed11ed856361be3be59dae656141fb0[0]        <=  I4156cb61e9e7e8947b6750f177dac22866e9f9ad06d7e45bdad1304988857d6f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I4156cb61e9e7e8947b6750f177dac22866e9f9ad06d7e45bdad1304988857d6f[0] + 1 :
                                             I4156cb61e9e7e8947b6750f177dac22866e9f9ad06d7e45bdad1304988857d6f[0] ;
            I7a94e46f1351801c2edf76bf3b70e3b5100b8e6108d60d9341591aa59f4e95d1[0]  <=  I4156cb61e9e7e8947b6750f177dac22866e9f9ad06d7e45bdad1304988857d6f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib41d86b318a3004b648c9a1b0ad00bbb144511fd63b1c7648cf3ccfb996686d3[0]        <=  I45ae7cee40ada2a73a62a90f141788d37c2a24f503646ce743ae4ac3e43b5bda[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I45ae7cee40ada2a73a62a90f141788d37c2a24f503646ce743ae4ac3e43b5bda[0] + 1 :
                                             I45ae7cee40ada2a73a62a90f141788d37c2a24f503646ce743ae4ac3e43b5bda[0] ;
            I0b761d71a88d70e6228dcf7325206f840d9da85892ba151c317e06079291fc2e[0]  <=  I45ae7cee40ada2a73a62a90f141788d37c2a24f503646ce743ae4ac3e43b5bda[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icc4bebb1db4145f9cce0fd4c250f7501f300b6cde1f31327d80b844adeeca1c7[0]        <=  I5ae0ab8d5ea922fff8bcc268c8f3bea87f11b7d6b824787e972c00a9db0be916[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5ae0ab8d5ea922fff8bcc268c8f3bea87f11b7d6b824787e972c00a9db0be916[0] + 1 :
                                             I5ae0ab8d5ea922fff8bcc268c8f3bea87f11b7d6b824787e972c00a9db0be916[0] ;
            Ic2ae521a3a6fef956f28a89da365b0838d535c9f7801a405cf60cc776ba0af2a[0]  <=  I5ae0ab8d5ea922fff8bcc268c8f3bea87f11b7d6b824787e972c00a9db0be916[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idead9dbad4283dce602c05f81e98610ab7f65f9911342174ceff7c95dfa9ddb0[0]        <=  Id33bc2a3f235239565a24ba23a93a90e564b2ddcc7559044ccd4f2e6aa6fdb6b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id33bc2a3f235239565a24ba23a93a90e564b2ddcc7559044ccd4f2e6aa6fdb6b[0] + 1 :
                                             Id33bc2a3f235239565a24ba23a93a90e564b2ddcc7559044ccd4f2e6aa6fdb6b[0] ;
            I01d9f8a8900be1981c601c0ccb45c1f39a0fdc16179245d80fbb2ad6d7060899[0]  <=  Id33bc2a3f235239565a24ba23a93a90e564b2ddcc7559044ccd4f2e6aa6fdb6b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If7060467d2fac9aee8d69c5ebdc24d515a657bedea3da55d13ed6ed4e3c8e79b[0]        <=  I86a468c8931c4e794856a1c434471a885c62c94dbbc95059bb67ec45a9a722b7[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I86a468c8931c4e794856a1c434471a885c62c94dbbc95059bb67ec45a9a722b7[0] + 1 :
                                             I86a468c8931c4e794856a1c434471a885c62c94dbbc95059bb67ec45a9a722b7[0] ;
            Icdfc2f0ce24f01af7df8a99b58de3a74e1dda0eea5b41ff2c342106cb226abdc[0]  <=  I86a468c8931c4e794856a1c434471a885c62c94dbbc95059bb67ec45a9a722b7[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6aefe769159bdc69fee8e09e46357993c13dd8ec9f059cd51d43944ecd7ce3ff[0]        <=  Ibc857d78e207a3c56616aab90400d7f0b57c62f4a5e421ee4b5b7ac7bfa1c31b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ibc857d78e207a3c56616aab90400d7f0b57c62f4a5e421ee4b5b7ac7bfa1c31b[0] + 1 :
                                             Ibc857d78e207a3c56616aab90400d7f0b57c62f4a5e421ee4b5b7ac7bfa1c31b[0] ;
            I929ef5474f10c76c4686fb044b2833b6ba1571f2e1c82b6d92cfaadfa44946e6[0]  <=  Ibc857d78e207a3c56616aab90400d7f0b57c62f4a5e421ee4b5b7ac7bfa1c31b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icac3a5cc88034cf8211c158a1bee2a04c228afd4eace1b50c7460ad5331ae02d[0]        <=  I275f7df80a91271f558b5ab22bb6a5b46f01973b93cccebe198f0f3c6e2f2cbe[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I275f7df80a91271f558b5ab22bb6a5b46f01973b93cccebe198f0f3c6e2f2cbe[0] + 1 :
                                             I275f7df80a91271f558b5ab22bb6a5b46f01973b93cccebe198f0f3c6e2f2cbe[0] ;
            I55312932ff9d69c8ffa1e42efdb5e775ccb21a8f9e8791b080b67654462e537a[0]  <=  I275f7df80a91271f558b5ab22bb6a5b46f01973b93cccebe198f0f3c6e2f2cbe[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ifa5d23491b028cbdcfd79fdea2e0784f068c1fd381dda7ebfb5d457800e510cd[0]        <=  I8cc2be0175b91e2589ee8980b860af09aaa4a81cedf23de18f9ae69d0514c369[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8cc2be0175b91e2589ee8980b860af09aaa4a81cedf23de18f9ae69d0514c369[0] + 1 :
                                             I8cc2be0175b91e2589ee8980b860af09aaa4a81cedf23de18f9ae69d0514c369[0] ;
            Icbdbaf4eb2f30bb78db34a582e06dc91689b9eab2f8fdfe4fbfb41a8cce93ca5[0]  <=  I8cc2be0175b91e2589ee8980b860af09aaa4a81cedf23de18f9ae69d0514c369[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic27b23bf87ceb2ec2d6460321286d798980f966c89d0f8ea42a79a0549b2128e[0]        <=  Ia6661480da7ffc0644e0a42782e89f84535952e5f17f2ecf3f1e4cfc56c532d5[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia6661480da7ffc0644e0a42782e89f84535952e5f17f2ecf3f1e4cfc56c532d5[0] + 1 :
                                             Ia6661480da7ffc0644e0a42782e89f84535952e5f17f2ecf3f1e4cfc56c532d5[0] ;
            Ifa4cbbd5c3ab5e47a7d5135e4dbaf365e79c4c6a806bfae88c9c0e1c9ffe2fa5[0]  <=  Ia6661480da7ffc0644e0a42782e89f84535952e5f17f2ecf3f1e4cfc56c532d5[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I01500dbf2528609729acf26a24c11bab0adf8cdbc0633527f21644816cfa0dc0[0]        <=  If4a3892f82907488395a090155f489b67d9808fab6c5f4cfccde65fc41d3b92f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If4a3892f82907488395a090155f489b67d9808fab6c5f4cfccde65fc41d3b92f[0] + 1 :
                                             If4a3892f82907488395a090155f489b67d9808fab6c5f4cfccde65fc41d3b92f[0] ;
            I2341907334935e19ef0e392216e39bb35c215730c464a85c0e1b804b364b492c[0]  <=  If4a3892f82907488395a090155f489b67d9808fab6c5f4cfccde65fc41d3b92f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6db96717b6fe00f1f87347adf69ce2d4b4464faa472ca989bb272b36454e868b[0]        <=  I7b2b5024c5f6f54ab62c8e703f603950e46ebd179fc35e2db34ace053564af4a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7b2b5024c5f6f54ab62c8e703f603950e46ebd179fc35e2db34ace053564af4a[0] + 1 :
                                             I7b2b5024c5f6f54ab62c8e703f603950e46ebd179fc35e2db34ace053564af4a[0] ;
            Ic0bbaf8314688690b5a15a5613ab149f604a8bfb92a2b9ed014e7ce2757d0743[0]  <=  I7b2b5024c5f6f54ab62c8e703f603950e46ebd179fc35e2db34ace053564af4a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia8cd57b3b123e08e2bc00f82da941eb4431cc816928254135dd13ef52eb9c03a[0]        <=  I709336ccea8dfb4b988c870e3d5c854d77a7acc5ff842b9c2c7490be8e10b3c3[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I709336ccea8dfb4b988c870e3d5c854d77a7acc5ff842b9c2c7490be8e10b3c3[0] + 1 :
                                             I709336ccea8dfb4b988c870e3d5c854d77a7acc5ff842b9c2c7490be8e10b3c3[0] ;
            I19ff0bebf62a994a2b5814ea41289f72cd62a38d2f37dc0027beb0f488926d4f[0]  <=  I709336ccea8dfb4b988c870e3d5c854d77a7acc5ff842b9c2c7490be8e10b3c3[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4fa8db615d84b02196afb2ad926769bcbfffb7c81170387b4d460c7403f0dfab[0]        <=  I6ad8cd22867ad477cef7562ef157f85bcd0aeb6ff72ceccd15ecf5c00faf12d6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6ad8cd22867ad477cef7562ef157f85bcd0aeb6ff72ceccd15ecf5c00faf12d6[0] + 1 :
                                             I6ad8cd22867ad477cef7562ef157f85bcd0aeb6ff72ceccd15ecf5c00faf12d6[0] ;
            I4f9435bbcce379d6d591547481382ab188003b97877c0f32462ef9e33aa8bc1a[0]  <=  I6ad8cd22867ad477cef7562ef157f85bcd0aeb6ff72ceccd15ecf5c00faf12d6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie81813a1836449254acfcf7674552545d2cbc852ee2bd2f37378345ccdfc61b4[0]        <=  If4a806d211914f82ca329f57517b2d1b1a60a8381bddbd3153e78418258d819e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If4a806d211914f82ca329f57517b2d1b1a60a8381bddbd3153e78418258d819e[0] + 1 :
                                             If4a806d211914f82ca329f57517b2d1b1a60a8381bddbd3153e78418258d819e[0] ;
            I9e497e3ee797c274b82ecca58218c47f9b663bcac21b1431b45c17d5e54e5a4a[0]  <=  If4a806d211914f82ca329f57517b2d1b1a60a8381bddbd3153e78418258d819e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id9fde3ad430d66c92a5aa6797b76ce147e39e4245ea761e36d81214e7a02b4d8[0]        <=  I282657b255db6edb8d72272a04f6c69d5b8f32795992f902cbedae3bffba4a4f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I282657b255db6edb8d72272a04f6c69d5b8f32795992f902cbedae3bffba4a4f[0] + 1 :
                                             I282657b255db6edb8d72272a04f6c69d5b8f32795992f902cbedae3bffba4a4f[0] ;
            Ib929181cef39d751d2726a054cd0478d309e58350ecd11d3363ecba8bd4cb7fa[0]  <=  I282657b255db6edb8d72272a04f6c69d5b8f32795992f902cbedae3bffba4a4f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8f2cae5483691fdf6ea64a4ccb2372967aa676835ffd4f562269bac888840d17[0]        <=  Ia3f8a8cdad50f5772d19748e82e1e9e0558a1d7973bc2cda424ba8d383c15d62[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia3f8a8cdad50f5772d19748e82e1e9e0558a1d7973bc2cda424ba8d383c15d62[0] + 1 :
                                             Ia3f8a8cdad50f5772d19748e82e1e9e0558a1d7973bc2cda424ba8d383c15d62[0] ;
            I64fa7f4fa09b7909840d8edb83f29f6a2379419e65b80f592b37d8ea00e59475[0]  <=  Ia3f8a8cdad50f5772d19748e82e1e9e0558a1d7973bc2cda424ba8d383c15d62[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icd8572ba29de1a399bc077f53730492f4e89deb95b9136608da0d029ba60ddd1[0]        <=  I9ec9a8bbe81467bd2ec058114005f308873b8eb8a8c939f4002003402bc6c486[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9ec9a8bbe81467bd2ec058114005f308873b8eb8a8c939f4002003402bc6c486[0] + 1 :
                                             I9ec9a8bbe81467bd2ec058114005f308873b8eb8a8c939f4002003402bc6c486[0] ;
            I35beac843abd6268c39acb691d3105a5c386f05461bca8c63b951ce1c2ed07bc[0]  <=  I9ec9a8bbe81467bd2ec058114005f308873b8eb8a8c939f4002003402bc6c486[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6eab6bb656dc82d656eea6da9dea574b230f56c6ab898a7f80973183896d8347[0]        <=  I2a951c202348bf2bb4da1f79c63a8515c95484c9a16ac1fe9b857fee59361511[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2a951c202348bf2bb4da1f79c63a8515c95484c9a16ac1fe9b857fee59361511[0] + 1 :
                                             I2a951c202348bf2bb4da1f79c63a8515c95484c9a16ac1fe9b857fee59361511[0] ;
            I9d8fbde44d35c50f5f24ceae6f2e16ca2f280573caeb8a3021b6f69dec3d04b4[0]  <=  I2a951c202348bf2bb4da1f79c63a8515c95484c9a16ac1fe9b857fee59361511[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Id802e388c3b33f7d0a0960e0e51da02e7128da423d518a916f761a16b73c17d7[0]        <=  I009b4951ca9d1200c6e7787f401228a9af483223fbb4150aca223cfbb80c8b7c[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I009b4951ca9d1200c6e7787f401228a9af483223fbb4150aca223cfbb80c8b7c[0] + 1 :
                                             I009b4951ca9d1200c6e7787f401228a9af483223fbb4150aca223cfbb80c8b7c[0] ;
            I507d851a78a765c18af6d529292384fb4cbb06cfec0e22d516adc79b8ea13c7f[0]  <=  I009b4951ca9d1200c6e7787f401228a9af483223fbb4150aca223cfbb80c8b7c[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I47507e717446a9ca85cec7e5fa382cfe435affddcbf5b25d4e74f23a143b02b0[0]        <=  I3af56e36e8422acbbdb52c77327e09618a7b89e21e35787ba522cb8a322ed0bd[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I3af56e36e8422acbbdb52c77327e09618a7b89e21e35787ba522cb8a322ed0bd[0] + 1 :
                                             I3af56e36e8422acbbdb52c77327e09618a7b89e21e35787ba522cb8a322ed0bd[0] ;
            I80fb8d450dd144ffade989cc2cec363cf6bbcdc267f5372163fde38313387499[0]  <=  I3af56e36e8422acbbdb52c77327e09618a7b89e21e35787ba522cb8a322ed0bd[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0d76ba051f3db8c1efd9a8f0bd0ca77cb28c7dfd68cf4c290ab00edfedb15237[0]        <=  Iea773cc6750944ca9d0aaaf2dbd818c485ce25a1e333978a68333b521404516d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iea773cc6750944ca9d0aaaf2dbd818c485ce25a1e333978a68333b521404516d[0] + 1 :
                                             Iea773cc6750944ca9d0aaaf2dbd818c485ce25a1e333978a68333b521404516d[0] ;
            I7844074cddcce1b95a010729a9e4ce2bfc4f7e1962b84af0e0a3cbb2c2c08206[0]  <=  Iea773cc6750944ca9d0aaaf2dbd818c485ce25a1e333978a68333b521404516d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I39dc59000bb2e3fcdebec08ddd22a460fad0c09e8b68adc7e72a6e4c3025da49[0]        <=  I5e0342048fa50ff3b98e175c5c8aabadb97e925dfbc34fb7f68376b8eaa3cb1f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5e0342048fa50ff3b98e175c5c8aabadb97e925dfbc34fb7f68376b8eaa3cb1f[0] + 1 :
                                             I5e0342048fa50ff3b98e175c5c8aabadb97e925dfbc34fb7f68376b8eaa3cb1f[0] ;
            I88be0c0499713ce396832a79853e9918ecdfed2519fba6fd7c0bae51450478e7[0]  <=  I5e0342048fa50ff3b98e175c5c8aabadb97e925dfbc34fb7f68376b8eaa3cb1f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6db1df05e1ea3d8011bbd6e08c9d50d91e672a20aa2448167343b839e8f6f888[0]        <=  Ie03375db3932197354d4fdbdc800b2b7134470f1622806909963ea424d5fe6af[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie03375db3932197354d4fdbdc800b2b7134470f1622806909963ea424d5fe6af[0] + 1 :
                                             Ie03375db3932197354d4fdbdc800b2b7134470f1622806909963ea424d5fe6af[0] ;
            Ib585733bf4c3eb59a772866965420fc7397b01272410cdb701f289daf9549fc9[0]  <=  Ie03375db3932197354d4fdbdc800b2b7134470f1622806909963ea424d5fe6af[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I0d11d2b76d26d33ebe0c7577f5d7bc68ab8f4840deb765b17f4f7fde0a4b2fae[0]        <=  I529cffab52c15bb4db9614fb7a0f353e2867564b31984bd2c5551f5a5d407fbb[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I529cffab52c15bb4db9614fb7a0f353e2867564b31984bd2c5551f5a5d407fbb[0] + 1 :
                                             I529cffab52c15bb4db9614fb7a0f353e2867564b31984bd2c5551f5a5d407fbb[0] ;
            Ida673298c761bab46fb26d4e73caa99f5b3ade7f924d99fcedae4e47c70b5b67[0]  <=  I529cffab52c15bb4db9614fb7a0f353e2867564b31984bd2c5551f5a5d407fbb[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ifbbf33f600185eab85dd2c0dc5ab2f5e0e2cce52373cc2acf5e466a2e27ded58[0]        <=  I3bd4e85424803f9f3607ec830b6c73bf1d273e7de387d11359eae7f842fb1551[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I3bd4e85424803f9f3607ec830b6c73bf1d273e7de387d11359eae7f842fb1551[0] + 1 :
                                             I3bd4e85424803f9f3607ec830b6c73bf1d273e7de387d11359eae7f842fb1551[0] ;
            I60bb81cc7cd9a6212f7b4261a21655accd6cd09e7aaf5f78f7f1f4dec0e8489b[0]  <=  I3bd4e85424803f9f3607ec830b6c73bf1d273e7de387d11359eae7f842fb1551[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia38b628fe0740039fd44aa0a75c751e1a9e176bfc305a978377c1fc9525c00e4[0]        <=  Ie54a4e9ee8bf7646b7e69193c8121ff42b4ab2f266c49916322dec059c92684d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie54a4e9ee8bf7646b7e69193c8121ff42b4ab2f266c49916322dec059c92684d[0] + 1 :
                                             Ie54a4e9ee8bf7646b7e69193c8121ff42b4ab2f266c49916322dec059c92684d[0] ;
            I85d3c885ce504524ab43daed7bbcb599cd7e5d6d3635cf46e278345134e97e22[0]  <=  Ie54a4e9ee8bf7646b7e69193c8121ff42b4ab2f266c49916322dec059c92684d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Iaeb5b860946e41cde629a762ab6e6ea4a0f177083c9ac84d90ca99fcb90e7c9a[0]        <=  Ic07553da54e29d977820e271e50502264b236c156bdf4e3a654cd948a6d4f726[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic07553da54e29d977820e271e50502264b236c156bdf4e3a654cd948a6d4f726[0] + 1 :
                                             Ic07553da54e29d977820e271e50502264b236c156bdf4e3a654cd948a6d4f726[0] ;
            Iaa08a49e0ca4f92f38c7f4d115ae1b275e45c42dfa6fd4b6a2ff40536b7f5f15[0]  <=  Ic07553da54e29d977820e271e50502264b236c156bdf4e3a654cd948a6d4f726[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ibc0b2c21012904530a727f0c5643b5187d7bb8706a308bdd0de67a80147db974[0]        <=  I8ba1954b4d7af696e80f659a70d18bea70c37a8f494827a2778c421ca1dd8ac9[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8ba1954b4d7af696e80f659a70d18bea70c37a8f494827a2778c421ca1dd8ac9[0] + 1 :
                                             I8ba1954b4d7af696e80f659a70d18bea70c37a8f494827a2778c421ca1dd8ac9[0] ;
            I197b3231cb1da107c5001075809e9fa75e4089871d473490981a8b44d3ff5e4c[0]  <=  I8ba1954b4d7af696e80f659a70d18bea70c37a8f494827a2778c421ca1dd8ac9[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I008d6180d4774d2472158544239ee654e73570389873b54b695946cb78ddb7e8[0]        <=  I2d1936d0e3bc9f6320f1311cbde5d8e855ebeb68cea0b8c3dcf77f3dd63ceb84[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I2d1936d0e3bc9f6320f1311cbde5d8e855ebeb68cea0b8c3dcf77f3dd63ceb84[0] + 1 :
                                             I2d1936d0e3bc9f6320f1311cbde5d8e855ebeb68cea0b8c3dcf77f3dd63ceb84[0] ;
            I384c04b75344f97c691f70965d7e08266ab9cd8862e04ba73b502a0f36ac5ea7[0]  <=  I2d1936d0e3bc9f6320f1311cbde5d8e855ebeb68cea0b8c3dcf77f3dd63ceb84[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idaea720265ed96d87e8852c36eebd63e2be5b9768c7803f13fe85e7532b75ea2[0]        <=  Ic0b3a57afcb2e31014f5c80d84c8eaf5f7f20d57abd8e863e6ffe0b8146108fd[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic0b3a57afcb2e31014f5c80d84c8eaf5f7f20d57abd8e863e6ffe0b8146108fd[0] + 1 :
                                             Ic0b3a57afcb2e31014f5c80d84c8eaf5f7f20d57abd8e863e6ffe0b8146108fd[0] ;
            Ibf95afb3941a2272d76cd7256d0789f11fb35a3020c3ccca5b099d335d4a2330[0]  <=  Ic0b3a57afcb2e31014f5c80d84c8eaf5f7f20d57abd8e863e6ffe0b8146108fd[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia7bf8296bff6d2322977b0a31ba519bca04a1d6c6f6c0cb5a47e3408bdfac573[0]        <=  Ia7f87cbac38cab3ef1ce6466b6b419127464ad3172cb03af43e0f75b9575ff2e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia7f87cbac38cab3ef1ce6466b6b419127464ad3172cb03af43e0f75b9575ff2e[0] + 1 :
                                             Ia7f87cbac38cab3ef1ce6466b6b419127464ad3172cb03af43e0f75b9575ff2e[0] ;
            I885622bb1c7371f4afa3e9966f870d2bf7750c2d2280a2a993a5bd9854187994[0]  <=  Ia7f87cbac38cab3ef1ce6466b6b419127464ad3172cb03af43e0f75b9575ff2e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2a69131c92e4454ec846c7528679731db69a2aa63420f0f22289d5c0be743be9[0]        <=  I27a670adbcc49dd11d8a6647a3220c4ac80946eae616e3da78e7a35f5f522502[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I27a670adbcc49dd11d8a6647a3220c4ac80946eae616e3da78e7a35f5f522502[0] + 1 :
                                             I27a670adbcc49dd11d8a6647a3220c4ac80946eae616e3da78e7a35f5f522502[0] ;
            I719a3e78d6a298f7db920bf7e355f6fca2c46135abb8ccd1cc3ea470912d05c1[0]  <=  I27a670adbcc49dd11d8a6647a3220c4ac80946eae616e3da78e7a35f5f522502[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia5fc094477d9d66d7fab491b73a00f50abec21827f63372fc1b7e0bd31ccf375[0]        <=  Ib913fea37f6ef92b53b6ec87dde4020983e78b263662b92008f7241cc029189a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib913fea37f6ef92b53b6ec87dde4020983e78b263662b92008f7241cc029189a[0] + 1 :
                                             Ib913fea37f6ef92b53b6ec87dde4020983e78b263662b92008f7241cc029189a[0] ;
            I1729b841d155c32b617727459f01aa9a9a6af56de5f464e20e900e3a4da30dba[0]  <=  Ib913fea37f6ef92b53b6ec87dde4020983e78b263662b92008f7241cc029189a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I41d88c1cdef0448f878686d88600bd254e722761979a244cb1d00724fc1d35d8[0]        <=  I1b653b0e5ffe67c25c7a73b1e2fc591f5e57174285113fe2c43ab123799c556a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I1b653b0e5ffe67c25c7a73b1e2fc591f5e57174285113fe2c43ab123799c556a[0] + 1 :
                                             I1b653b0e5ffe67c25c7a73b1e2fc591f5e57174285113fe2c43ab123799c556a[0] ;
            I96affe6d042e09b07278ae45744977fd3719a31fa5d578adaa2b3a66b2c3ebd0[0]  <=  I1b653b0e5ffe67c25c7a73b1e2fc591f5e57174285113fe2c43ab123799c556a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I85e825a905ae7dd292f400406048736ce90fa7d47b6dc5507254283662fc7564[0]        <=  I068d321d442274e43788076aecb6c24130003e03ced4df86bf13a33d2ca5e1f0[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I068d321d442274e43788076aecb6c24130003e03ced4df86bf13a33d2ca5e1f0[0] + 1 :
                                             I068d321d442274e43788076aecb6c24130003e03ced4df86bf13a33d2ca5e1f0[0] ;
            I12e1e01b28d2d443785fac1d0314b477b221b17b715f1153c5379a85b4b5e3aa[0]  <=  I068d321d442274e43788076aecb6c24130003e03ced4df86bf13a33d2ca5e1f0[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I80cf17357df8073b050d80de366bbb919c5f6c8983ca87f6606a84df1b92c549[0]        <=  I975a1d7b1fe781bb19e80aba369e5146327185746eb5088542eba76fbd88ddbe[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I975a1d7b1fe781bb19e80aba369e5146327185746eb5088542eba76fbd88ddbe[0] + 1 :
                                             I975a1d7b1fe781bb19e80aba369e5146327185746eb5088542eba76fbd88ddbe[0] ;
            Ie244ea5cb57e0b4c14c0c8c22592347d1389a6b0f53b821335b821ca5130ad6e[0]  <=  I975a1d7b1fe781bb19e80aba369e5146327185746eb5088542eba76fbd88ddbe[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I68a074e808119d0f33d54d3863c907dd5d761b3f6b144b9283e67f956d5932ef[0]        <=  I6668b8618eebf7c40e35e5a06aa3b131a6ea1b668bc36d9731036b61087013c3[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6668b8618eebf7c40e35e5a06aa3b131a6ea1b668bc36d9731036b61087013c3[0] + 1 :
                                             I6668b8618eebf7c40e35e5a06aa3b131a6ea1b668bc36d9731036b61087013c3[0] ;
            I5a07f349b1fd7d668d35583c50dfa3ceda070e5dc241bff1ecdddace6624bd57[0]  <=  I6668b8618eebf7c40e35e5a06aa3b131a6ea1b668bc36d9731036b61087013c3[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4aab61ec97ec8dfc8da6d2ab5898bcdfdaebb0f024fea498a6ecbf0bd15fd1c5[0]        <=  I1b4f3dc17b05ab02ad55643162e80975cc4802ba8cbc4323fb017859b3617abb[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I1b4f3dc17b05ab02ad55643162e80975cc4802ba8cbc4323fb017859b3617abb[0] + 1 :
                                             I1b4f3dc17b05ab02ad55643162e80975cc4802ba8cbc4323fb017859b3617abb[0] ;
            I6e5f194e3acb27a7fdd060e05aff00bb9fcd0904b3f920d7db0fee84c1534558[0]  <=  I1b4f3dc17b05ab02ad55643162e80975cc4802ba8cbc4323fb017859b3617abb[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I26395ccf79a44d582b559acac5845eae4a01464019f7739b7d52d8c8a4c11154[0]        <=  Ic69eaf55d245ae896d42f0f702ef6cd804be0d02cfad9f883b3dac30786352d9[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic69eaf55d245ae896d42f0f702ef6cd804be0d02cfad9f883b3dac30786352d9[0] + 1 :
                                             Ic69eaf55d245ae896d42f0f702ef6cd804be0d02cfad9f883b3dac30786352d9[0] ;
            I09780397509ca78f4b4aed5b08cf22d8eae797d1d1864cdba4a951ac8d583c91[0]  <=  Ic69eaf55d245ae896d42f0f702ef6cd804be0d02cfad9f883b3dac30786352d9[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie9c493e499f4b2aa598c54d5a5afdf39447612225daf7f9f5b3c2a23b5ee0ff0[0]        <=  I8c815413903d61f8d5f9a8abbb8b5e6cb133bcf0e084f4a46ceb98fc67f67515[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8c815413903d61f8d5f9a8abbb8b5e6cb133bcf0e084f4a46ceb98fc67f67515[0] + 1 :
                                             I8c815413903d61f8d5f9a8abbb8b5e6cb133bcf0e084f4a46ceb98fc67f67515[0] ;
            Iefcb9b5b2f238005d0f37bc519349bbbc130e3e072814ec48b4edf9c853a6913[0]  <=  I8c815413903d61f8d5f9a8abbb8b5e6cb133bcf0e084f4a46ceb98fc67f67515[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4368873c6f3e3d6ba5e7e83747fb90120e80de634655a9d2a97bbee88a9d8501[0]        <=  I6abdbd209c6b52b3d4c69e83d51d89be9b3b8e719e4f4e15f50afdccb21ea02b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6abdbd209c6b52b3d4c69e83d51d89be9b3b8e719e4f4e15f50afdccb21ea02b[0] + 1 :
                                             I6abdbd209c6b52b3d4c69e83d51d89be9b3b8e719e4f4e15f50afdccb21ea02b[0] ;
            I9835f6f38580d8765566723f5a9adbfb4935af8bf719b3e4918e1b746cf12241[0]  <=  I6abdbd209c6b52b3d4c69e83d51d89be9b3b8e719e4f4e15f50afdccb21ea02b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I082b315a51a6a180909ea4f576a9a3c8b0550e64aa222610c2e6906ca78aebad[0]        <=  I6f2bfa7344a4516d6e0b959405ab2c16aabea8d70a454d4eab330ffb6bf9ce2d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6f2bfa7344a4516d6e0b959405ab2c16aabea8d70a454d4eab330ffb6bf9ce2d[0] + 1 :
                                             I6f2bfa7344a4516d6e0b959405ab2c16aabea8d70a454d4eab330ffb6bf9ce2d[0] ;
            I2266ca44e019a30bb553f955a158a5b075035c4b20a0b3fca6a3675ec79b9997[0]  <=  I6f2bfa7344a4516d6e0b959405ab2c16aabea8d70a454d4eab330ffb6bf9ce2d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I23872b1af6db7e455f25a7ddcc050167bb10de0afd16973c0a90804349210372[0]        <=  Ie7eedf6171b2af8aa5e550f07c6913fc6e02bde23689f5ff9f035b89ea7f4cfb[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie7eedf6171b2af8aa5e550f07c6913fc6e02bde23689f5ff9f035b89ea7f4cfb[0] + 1 :
                                             Ie7eedf6171b2af8aa5e550f07c6913fc6e02bde23689f5ff9f035b89ea7f4cfb[0] ;
            I684ec077e37638f022f10b5eb31403e6f9117a83a606f2a5013c2c33b8d1a8ab[0]  <=  Ie7eedf6171b2af8aa5e550f07c6913fc6e02bde23689f5ff9f035b89ea7f4cfb[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9796589e7a8535d47d56f792d80838aa402e3c235035b517765096d2a6843215[0]        <=  Ia298bc83a87ee16d194185dec24955ca32e85a919f168cbfc79e0724038e43d4[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia298bc83a87ee16d194185dec24955ca32e85a919f168cbfc79e0724038e43d4[0] + 1 :
                                             Ia298bc83a87ee16d194185dec24955ca32e85a919f168cbfc79e0724038e43d4[0] ;
            I9331428911b817ea45d1b5ae75eb3ee6e05c189785c995e5d2625f12ce4e0846[0]  <=  Ia298bc83a87ee16d194185dec24955ca32e85a919f168cbfc79e0724038e43d4[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46d39260d96216c08b7940ea3bfe542bdbd0966f5e798321bc90a2a00f64360f[0]        <=  I78dfe767d8265759b3b1488f6788812b210a952cba86301b7afe8acd0b194947[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I78dfe767d8265759b3b1488f6788812b210a952cba86301b7afe8acd0b194947[0] + 1 :
                                             I78dfe767d8265759b3b1488f6788812b210a952cba86301b7afe8acd0b194947[0] ;
            I7769e8ceb72790c37b351c32983860280aef172974d19a2e99348607863a97d4[0]  <=  I78dfe767d8265759b3b1488f6788812b210a952cba86301b7afe8acd0b194947[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I1033817563ce88e3b26188a88303cc6703f47afdaae4d5457fab8b73bade5274[0]        <=  I12a747458626b92b4c562f72f3e5fb63a575053284698acfde64b482d44a98b7[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I12a747458626b92b4c562f72f3e5fb63a575053284698acfde64b482d44a98b7[0] + 1 :
                                             I12a747458626b92b4c562f72f3e5fb63a575053284698acfde64b482d44a98b7[0] ;
            If09c36408407b246848b29df63e789fd1041815243beb4f27db0e774e853f1cd[0]  <=  I12a747458626b92b4c562f72f3e5fb63a575053284698acfde64b482d44a98b7[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I343bc73eaaf00a82b2674c8cdfbbc5c6ea52d10fbb9e9453cf4fcf2421b97e47[0]        <=  Id27fc6b236852c780351e17ad6e85bf55621c84757b3014ead5a2b9ef31d2ce8[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id27fc6b236852c780351e17ad6e85bf55621c84757b3014ead5a2b9ef31d2ce8[0] + 1 :
                                             Id27fc6b236852c780351e17ad6e85bf55621c84757b3014ead5a2b9ef31d2ce8[0] ;
            I533b63eedc528cb36abc0a469b66b144a6ae5122c038eef85d8d0557c3dff3ea[0]  <=  Id27fc6b236852c780351e17ad6e85bf55621c84757b3014ead5a2b9ef31d2ce8[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I1af6f4d00567aa1e302e7d8830d761e7a9a616f5e4e958b264701c476216de4f[0]        <=  Ic117e33adf22ba594c3e3c03966b6bb0c6827c2c980f6ba1ee5f6ba40da372dc[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ic117e33adf22ba594c3e3c03966b6bb0c6827c2c980f6ba1ee5f6ba40da372dc[0] + 1 :
                                             Ic117e33adf22ba594c3e3c03966b6bb0c6827c2c980f6ba1ee5f6ba40da372dc[0] ;
            I051e3b709db2e7861d31165ec1e5ee679f1e6dffa5a951072831ce479c16f27f[0]  <=  Ic117e33adf22ba594c3e3c03966b6bb0c6827c2c980f6ba1ee5f6ba40da372dc[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I1682f44d820722e2566b0d6c02fbf3dc72547221d519ed071e7c7d77728ba21e[0]        <=  I223d1009ee5643d0804f1d58bbeee2c3f61d8b120ceadf46556e379e45ccc061[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I223d1009ee5643d0804f1d58bbeee2c3f61d8b120ceadf46556e379e45ccc061[0] + 1 :
                                             I223d1009ee5643d0804f1d58bbeee2c3f61d8b120ceadf46556e379e45ccc061[0] ;
            I2fa018ce903921d0a174a63dbbb29eea8d5700b376335b2ba9bd448e8782018a[0]  <=  I223d1009ee5643d0804f1d58bbeee2c3f61d8b120ceadf46556e379e45ccc061[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If0095cd5e911c91331d2ef6ab3866101080b3cabe8d1ba9104b6b5ae5d18c713[0]        <=  I60bf67e044d9694caec17617c4d9ff59b9be7698c17aa034515ab1cc94d6a5ed[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I60bf67e044d9694caec17617c4d9ff59b9be7698c17aa034515ab1cc94d6a5ed[0] + 1 :
                                             I60bf67e044d9694caec17617c4d9ff59b9be7698c17aa034515ab1cc94d6a5ed[0] ;
            I36e06c1d77080ff75778f3dfa4ed60e66f9a3bedc39b214e3fdb5b6c21f1cd3e[0]  <=  I60bf67e044d9694caec17617c4d9ff59b9be7698c17aa034515ab1cc94d6a5ed[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If7f60dea1e83c3f86ff8ce3adda8214324b2064d06d69ca68477288522ad9de0[0]        <=  I7da66be74fda28e419201be145b24b82c9b29d1155ed00f78e8907d584e214c1[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7da66be74fda28e419201be145b24b82c9b29d1155ed00f78e8907d584e214c1[0] + 1 :
                                             I7da66be74fda28e419201be145b24b82c9b29d1155ed00f78e8907d584e214c1[0] ;
            Id647e3bd88fdc7a3642092d071f66f74657c8364937caf63c723f1e027c157bc[0]  <=  I7da66be74fda28e419201be145b24b82c9b29d1155ed00f78e8907d584e214c1[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I3b1abc53d350b3b39e60c3a5725e5a21632e7f0275988b98c1fdaeed5342f9c0[0]        <=  Idfaa10639faa52207bae09b46b05e70da4e285f83560fc415e3915d0a0e8fa4b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idfaa10639faa52207bae09b46b05e70da4e285f83560fc415e3915d0a0e8fa4b[0] + 1 :
                                             Idfaa10639faa52207bae09b46b05e70da4e285f83560fc415e3915d0a0e8fa4b[0] ;
            I015b73e7e4bc4c2a3073a304e58d24f5c8c32e90299f004bc0f75eb9e18e6d41[0]  <=  Idfaa10639faa52207bae09b46b05e70da4e285f83560fc415e3915d0a0e8fa4b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7943272afdae80761f8b673788c92e4461bf3de3229f7addec1e54743b11beca[0]        <=  Ifc9a7a5a4da00db6f00362e2b2b91e1ca59a65e8e35d66791a13468302dd081f[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ifc9a7a5a4da00db6f00362e2b2b91e1ca59a65e8e35d66791a13468302dd081f[0] + 1 :
                                             Ifc9a7a5a4da00db6f00362e2b2b91e1ca59a65e8e35d66791a13468302dd081f[0] ;
            I7c211cef6a581c5a6871d4c9a2b7ba29a9d05d36b0a758106e006caebfc592e5[0]  <=  Ifc9a7a5a4da00db6f00362e2b2b91e1ca59a65e8e35d66791a13468302dd081f[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I8417f8f367de885ebb86571786bd964d4a81d6712a88c3a8071c08d13cc7cf58[0]        <=  If453fce64c627db639d688b2260fa70ef90f802d31cac666fd4cd757cd574682[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If453fce64c627db639d688b2260fa70ef90f802d31cac666fd4cd757cd574682[0] + 1 :
                                             If453fce64c627db639d688b2260fa70ef90f802d31cac666fd4cd757cd574682[0] ;
            I3f2014435aac47a3c807e9ad3f0829179f9285582b7ff2e3bae250a25e800aee[0]  <=  If453fce64c627db639d688b2260fa70ef90f802d31cac666fd4cd757cd574682[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I653822ee3643c81b817be0d9c3f682d0c806ae17dedb0cae5b1aa0ca914e6857[0]        <=  I1eca2d1c9da79ade1c32a3685553f133098e1e40edd1e8d9c299a961627aefbb[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I1eca2d1c9da79ade1c32a3685553f133098e1e40edd1e8d9c299a961627aefbb[0] + 1 :
                                             I1eca2d1c9da79ade1c32a3685553f133098e1e40edd1e8d9c299a961627aefbb[0] ;
            Ib27fb4891a6edd486a99f23a750057de12a5a3e3fc6a5fad7976aa7e961e0c54[0]  <=  I1eca2d1c9da79ade1c32a3685553f133098e1e40edd1e8d9c299a961627aefbb[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ieb917f5db48f3d352eb252f6ce309bd972cab47f09ba1c140f66192b260f3925[0]        <=  Id3b8c5a0992cfb8a82d0e9857a0a77472fe0435d93e37978bc77770999bc4b4d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id3b8c5a0992cfb8a82d0e9857a0a77472fe0435d93e37978bc77770999bc4b4d[0] + 1 :
                                             Id3b8c5a0992cfb8a82d0e9857a0a77472fe0435d93e37978bc77770999bc4b4d[0] ;
            Ib58cd067e009a5f4b72af8cfb1e5c49c18f51a2ad8880f65aee683bf8ecd40ad[0]  <=  Id3b8c5a0992cfb8a82d0e9857a0a77472fe0435d93e37978bc77770999bc4b4d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I313a01d9fe403e838310c49dc37a50b738025400e99faefbd9b8cbd426edcfaa[0]        <=  Ia5acd518b995f7c0cb3e2f5303601027e6195fb82489331aa60c3fc8dfb21184[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ia5acd518b995f7c0cb3e2f5303601027e6195fb82489331aa60c3fc8dfb21184[0] + 1 :
                                             Ia5acd518b995f7c0cb3e2f5303601027e6195fb82489331aa60c3fc8dfb21184[0] ;
            I7e40bd6625b1d7deff82f67d46817c7af70f1da57561ab528b553b3d244b3f1d[0]  <=  Ia5acd518b995f7c0cb3e2f5303601027e6195fb82489331aa60c3fc8dfb21184[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I1b81a8a827bd2222ea6820d80d13e537868e0157970625d628f0c062733ec3d4[0]        <=  I588a95ce70c7581d9afef4d4a297b619958d34acc8bb75e4d61729b440945a89[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I588a95ce70c7581d9afef4d4a297b619958d34acc8bb75e4d61729b440945a89[0] + 1 :
                                             I588a95ce70c7581d9afef4d4a297b619958d34acc8bb75e4d61729b440945a89[0] ;
            I01949f24f74578cb63dd095e8ce639ce0d273c14da81e75d00097535e391aa4c[0]  <=  I588a95ce70c7581d9afef4d4a297b619958d34acc8bb75e4d61729b440945a89[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5615438871373f7ad838fb5e8c24b9517fb94ecf6627c803e66a78f778fe9c42[0]        <=  Idaeda6020813227d8f52db3ade5daa8152deb71aad3e8cd03094b66b7af5696c[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Idaeda6020813227d8f52db3ade5daa8152deb71aad3e8cd03094b66b7af5696c[0] + 1 :
                                             Idaeda6020813227d8f52db3ade5daa8152deb71aad3e8cd03094b66b7af5696c[0] ;
            Id8f2a0d3524b27621ca5a576bf16e15789e6257060225da04da2a5fcc8cf751e[0]  <=  Idaeda6020813227d8f52db3ade5daa8152deb71aad3e8cd03094b66b7af5696c[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I07f9ecb15d2696b2cacc35c935b497b2f8cedc55e2a661fa57f2d0783e6a1001[0]        <=  I48f239b0c336ab3fdd25e5b7758a5e6c3c0e698832c1f4518d3d1bc6845acd41[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I48f239b0c336ab3fdd25e5b7758a5e6c3c0e698832c1f4518d3d1bc6845acd41[0] + 1 :
                                             I48f239b0c336ab3fdd25e5b7758a5e6c3c0e698832c1f4518d3d1bc6845acd41[0] ;
            I6020dcffd9e047c03740cffcdfe790eaf614ea1036a50fefcec9e13e5b5ac4bc[0]  <=  I48f239b0c336ab3fdd25e5b7758a5e6c3c0e698832c1f4518d3d1bc6845acd41[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7fbeac90b85dfc78e20281021fc1d7cc90f9deacb2091ab55ed07f51fbdbcc11[0]        <=  I7226b2d9a70f4f716635a08aacafd4ef7a6f5fd31edaee6654bac5577e6398c4[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I7226b2d9a70f4f716635a08aacafd4ef7a6f5fd31edaee6654bac5577e6398c4[0] + 1 :
                                             I7226b2d9a70f4f716635a08aacafd4ef7a6f5fd31edaee6654bac5577e6398c4[0] ;
            I815f772d86db329f78fa75c3326c129ccf0f6c5f383b42ef18033e48d11525d2[0]  <=  I7226b2d9a70f4f716635a08aacafd4ef7a6f5fd31edaee6654bac5577e6398c4[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I46dfb75396740f84b7758552420a7ba8693bb1ca5259a67530c588585de1c337[0]        <=  I14a8ff2f5afad37ef2f9494e67d6fc7df5e0960766ad9f9c46964287587df5ed[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I14a8ff2f5afad37ef2f9494e67d6fc7df5e0960766ad9f9c46964287587df5ed[0] + 1 :
                                             I14a8ff2f5afad37ef2f9494e67d6fc7df5e0960766ad9f9c46964287587df5ed[0] ;
            I2c8a33831a21c4c21dd58a300467abcc82d52e7636a73a12a003a4144d43e0dc[0]  <=  I14a8ff2f5afad37ef2f9494e67d6fc7df5e0960766ad9f9c46964287587df5ed[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I60e36bd866a477c35110e2688e7fbb13b0303d210e014c9e151b313d130101a8[0]        <=  I0b4e726e030569d30af5272062eab7426f9a6c50a8e71353fc19fa3b0d576de6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I0b4e726e030569d30af5272062eab7426f9a6c50a8e71353fc19fa3b0d576de6[0] + 1 :
                                             I0b4e726e030569d30af5272062eab7426f9a6c50a8e71353fc19fa3b0d576de6[0] ;
            I8c7b9ead4ab28ae2c2aa5185a0746c9cfe9fd90bdd68f2ba05291045a296d566[0]  <=  I0b4e726e030569d30af5272062eab7426f9a6c50a8e71353fc19fa3b0d576de6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ibb36dcaba8439f48b18ad2dc8399df26b940f7cd815996635da092d41ee5b106[0]        <=  Ib6234dcd7696dadb4fa7903f2da1ddf0a7f469668b59cde104d9fd751ebea2cb[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib6234dcd7696dadb4fa7903f2da1ddf0a7f469668b59cde104d9fd751ebea2cb[0] + 1 :
                                             Ib6234dcd7696dadb4fa7903f2da1ddf0a7f469668b59cde104d9fd751ebea2cb[0] ;
            I32ed4ecd4363760151c1accda085c9afa3efe63daf7a312feefc00b804401c27[0]  <=  Ib6234dcd7696dadb4fa7903f2da1ddf0a7f469668b59cde104d9fd751ebea2cb[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I387a4fa48a52a029d2bb0c8e5163f15c4cd55d570db8d89e5f73d7bd6e21ae5b[0]        <=  I07dcbe17d78ed40700955c3277dc667bccfdb936125e6bf04e0e0ed08eafedea[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I07dcbe17d78ed40700955c3277dc667bccfdb936125e6bf04e0e0ed08eafedea[0] + 1 :
                                             I07dcbe17d78ed40700955c3277dc667bccfdb936125e6bf04e0e0ed08eafedea[0] ;
            I6aa6d6c6213348ea0cc3e8b207bca2c1db81499441e4ed721ca0ee01ae831291[0]  <=  I07dcbe17d78ed40700955c3277dc667bccfdb936125e6bf04e0e0ed08eafedea[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie2ad7096c10eafa6e451ff7793b2dda562b6623b1eaeed56bbad4019662851ac[0]        <=  Ie14f4f4bb4b43f4c07d648f32e6470bc1626117d46a927a286a64d093110e0f9[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie14f4f4bb4b43f4c07d648f32e6470bc1626117d46a927a286a64d093110e0f9[0] + 1 :
                                             Ie14f4f4bb4b43f4c07d648f32e6470bc1626117d46a927a286a64d093110e0f9[0] ;
            Ib4f23d2e5f8c73110ae24212c4ec0e7ef29c09c8178ec3850f061a5b0386feca[0]  <=  Ie14f4f4bb4b43f4c07d648f32e6470bc1626117d46a927a286a64d093110e0f9[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9de97cb2569312c40a541c0038e02c03024581050590e5677dcde888f4c6c3ac[0]        <=  I099c775595305f8021cc03ef225be27441e325455935c0545cdc553d0fea3d44[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I099c775595305f8021cc03ef225be27441e325455935c0545cdc553d0fea3d44[0] + 1 :
                                             I099c775595305f8021cc03ef225be27441e325455935c0545cdc553d0fea3d44[0] ;
            If2be986b27ce8aa2117f87e9a144015a10acf0a07847f83acec2804b9e987e8b[0]  <=  I099c775595305f8021cc03ef225be27441e325455935c0545cdc553d0fea3d44[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7a55e4af3d00a3684ba08ac52c3dc7dd0188efbb684b859ecf017f783fce247a[0]        <=  I9bfa196a8246cf5ae88343b221c084738279254b84fc66495e4669083ac05ad1[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9bfa196a8246cf5ae88343b221c084738279254b84fc66495e4669083ac05ad1[0] + 1 :
                                             I9bfa196a8246cf5ae88343b221c084738279254b84fc66495e4669083ac05ad1[0] ;
            I9f17331c6a9858b60705d889b5b77078042cffe9e956de20eb067ad7e70626b7[0]  <=  I9bfa196a8246cf5ae88343b221c084738279254b84fc66495e4669083ac05ad1[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib1644713e1c2c63d093c8af3a2be146dabd70cfe25a1a6ac062174576477b113[0]        <=  I9fb047739860e32f32c612e35c96205de22487ff301c0fc990f576bf205b98fd[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9fb047739860e32f32c612e35c96205de22487ff301c0fc990f576bf205b98fd[0] + 1 :
                                             I9fb047739860e32f32c612e35c96205de22487ff301c0fc990f576bf205b98fd[0] ;
            I2b70416e96231188e62b7bcf0300c4a5b2d2139449150d31414b92ae075aa0e7[0]  <=  I9fb047739860e32f32c612e35c96205de22487ff301c0fc990f576bf205b98fd[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie907506d9949011db3e41c72b9581fb832dfb29f82249768fd9893a3de358b35[0]        <=  Ib5aae92803bb8df9f7ffc9fe70a6f447be999b64f9d698828709487924cdd4db[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ib5aae92803bb8df9f7ffc9fe70a6f447be999b64f9d698828709487924cdd4db[0] + 1 :
                                             Ib5aae92803bb8df9f7ffc9fe70a6f447be999b64f9d698828709487924cdd4db[0] ;
            I29599a1dac362c87f4780a94478787a718f63401d2051ccbfe543b44e49b35bb[0]  <=  Ib5aae92803bb8df9f7ffc9fe70a6f447be999b64f9d698828709487924cdd4db[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I678204e14a0213dfa7135814f07e5f6c4d12452a503ed555ca2c20c10f047d5d[0]        <=  Id89ea99f9b791029af271f9916f63681c6881dec4351cd30a7fc9e3ff1b81400[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id89ea99f9b791029af271f9916f63681c6881dec4351cd30a7fc9e3ff1b81400[0] + 1 :
                                             Id89ea99f9b791029af271f9916f63681c6881dec4351cd30a7fc9e3ff1b81400[0] ;
            I5ff7defb023005e77164f9f3b852fa60ce897922c6b814015d3436fe1d1b4a44[0]  <=  Id89ea99f9b791029af271f9916f63681c6881dec4351cd30a7fc9e3ff1b81400[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ice68b876a3b3943637914d8d12aec7fd37cb867f7a7c20be11a66dd85803827d[0]        <=  I8f70e2b5b2ffcd04b7a84ba28ab51f0a9dafd95e4628df8b36dba0ccf87c666d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8f70e2b5b2ffcd04b7a84ba28ab51f0a9dafd95e4628df8b36dba0ccf87c666d[0] + 1 :
                                             I8f70e2b5b2ffcd04b7a84ba28ab51f0a9dafd95e4628df8b36dba0ccf87c666d[0] ;
            Ie132a24e667376de85b8fff9a639698df164043422122a8058c968bb7996d3a7[0]  <=  I8f70e2b5b2ffcd04b7a84ba28ab51f0a9dafd95e4628df8b36dba0ccf87c666d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I35e112474e97e65f8e8aa9a4dcce274c7ffda9cdef901ba31801b4daa68888fe[0]        <=  I21a71d60d8728a63954973b41b85f8ec46e1fedcb5208ea2397adfa9e58be880[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I21a71d60d8728a63954973b41b85f8ec46e1fedcb5208ea2397adfa9e58be880[0] + 1 :
                                             I21a71d60d8728a63954973b41b85f8ec46e1fedcb5208ea2397adfa9e58be880[0] ;
            Ie8d5dfc9a77dc01055a551c5f37416d0b13ef83428bf751fb9f95c7d10442697[0]  <=  I21a71d60d8728a63954973b41b85f8ec46e1fedcb5208ea2397adfa9e58be880[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I84992c3714fef30f928dc3330821045f20e176826278d42a9606f2dfadfcb9c8[0]        <=  Icc2b71964c3f1484faf865db6f25dadf0a84b62f85a86cae24a8c01baa1ce8ec[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icc2b71964c3f1484faf865db6f25dadf0a84b62f85a86cae24a8c01baa1ce8ec[0] + 1 :
                                             Icc2b71964c3f1484faf865db6f25dadf0a84b62f85a86cae24a8c01baa1ce8ec[0] ;
            Ic94f2b10208cb23bb5f5b1a46c11c3bbae038308b385373cfaad9a18e09ccb90[0]  <=  Icc2b71964c3f1484faf865db6f25dadf0a84b62f85a86cae24a8c01baa1ce8ec[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I011fbcda61a4f528c38920d0077565c4592c5f6d1a2f5a1a7dcb6a4a734e0c83[0]        <=  Ief6bd3a84efa60cd8d09e7f71dc4b3b882f2eeef86edace8634b6355a0ce5db2[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ief6bd3a84efa60cd8d09e7f71dc4b3b882f2eeef86edace8634b6355a0ce5db2[0] + 1 :
                                             Ief6bd3a84efa60cd8d09e7f71dc4b3b882f2eeef86edace8634b6355a0ce5db2[0] ;
            I3b79a6c69be124aeea9d1444f9f985201b55ad0d7a4767a01f612eee12a6ad73[0]  <=  Ief6bd3a84efa60cd8d09e7f71dc4b3b882f2eeef86edace8634b6355a0ce5db2[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6d2154a30adb0faf296cf58ca9229eb1a298767fccc4a1214092a2b977f7442f[0]        <=  I21ed781b8a01923a17f646d965cd22caccb44b555b8f392387269b9a2ec9b647[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I21ed781b8a01923a17f646d965cd22caccb44b555b8f392387269b9a2ec9b647[0] + 1 :
                                             I21ed781b8a01923a17f646d965cd22caccb44b555b8f392387269b9a2ec9b647[0] ;
            Id3ac4bf805d3981ac1eb1b396b3da5c0dbc68754d89668f0a4cf7c6f2a44ddfa[0]  <=  I21ed781b8a01923a17f646d965cd22caccb44b555b8f392387269b9a2ec9b647[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie500f9b1405b49a263908c145ee4a337f2ba4cd2d4d784a2acb77068d09d1662[0]        <=  If070967e597fbcb6a0ce8a28166d084e71daea6fec72b92cad9a59d03c2dc531[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If070967e597fbcb6a0ce8a28166d084e71daea6fec72b92cad9a59d03c2dc531[0] + 1 :
                                             If070967e597fbcb6a0ce8a28166d084e71daea6fec72b92cad9a59d03c2dc531[0] ;
            Id77fd99c6146776bfc20804c67ae41b88cb0441eecba4f40b87828956b7158b6[0]  <=  If070967e597fbcb6a0ce8a28166d084e71daea6fec72b92cad9a59d03c2dc531[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I26997f7f737ba99dcbde55d67661cf9e4efecf397b1ab3ec59e0cc5d8654a75c[0]        <=  Ie0c16d4ccdd2d7d6d9e45d2eea233e13674b7d5a1f8f41877267074f40f6a2bf[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Ie0c16d4ccdd2d7d6d9e45d2eea233e13674b7d5a1f8f41877267074f40f6a2bf[0] + 1 :
                                             Ie0c16d4ccdd2d7d6d9e45d2eea233e13674b7d5a1f8f41877267074f40f6a2bf[0] ;
            I650a7220fd4eb743f652c6c1f9431191621f9fb1a5b5d64bb9649b43bad5b8bf[0]  <=  Ie0c16d4ccdd2d7d6d9e45d2eea233e13674b7d5a1f8f41877267074f40f6a2bf[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            If6181a32c0ba3cb93e47ed1f1279bd4e739882c2905d6d64d0149f26d052f0d0[0]        <=  I731f6a3be9c5a884fe93ef383fd933c14af1cfb64cd73fc4381d91d4faa2757d[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I731f6a3be9c5a884fe93ef383fd933c14af1cfb64cd73fc4381d91d4faa2757d[0] + 1 :
                                             I731f6a3be9c5a884fe93ef383fd933c14af1cfb64cd73fc4381d91d4faa2757d[0] ;
            Ib7417e90e9dc35367f110c364878657dbbf66b1a714d5807e6347095b833c62d[0]  <=  I731f6a3be9c5a884fe93ef383fd933c14af1cfb64cd73fc4381d91d4faa2757d[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Idb4bd19284288df2a5b701cedcd57347e4f7c37947ec1588daedf3c9ede0a12e[0]        <=  I77f33c069479b582cee609a1e4f6255628bb7f6f667e6536333c8e99dac1e08e[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I77f33c069479b582cee609a1e4f6255628bb7f6f667e6536333c8e99dac1e08e[0] + 1 :
                                             I77f33c069479b582cee609a1e4f6255628bb7f6f667e6536333c8e99dac1e08e[0] ;
            Ie59a4afbd0d65de2149e8c60229bce12b77f8f1b2b232a11fb9714371eced2b9[0]  <=  I77f33c069479b582cee609a1e4f6255628bb7f6f667e6536333c8e99dac1e08e[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I4be880e4f25fc41932b9ab9295794ffa2f334ee5338ef0d59894d18918d3e0be[0]        <=  I9288b2d29db5e8dbeef47da923a8ea2055a38ca1f37d4d8ed5d458408b154924[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9288b2d29db5e8dbeef47da923a8ea2055a38ca1f37d4d8ed5d458408b154924[0] + 1 :
                                             I9288b2d29db5e8dbeef47da923a8ea2055a38ca1f37d4d8ed5d458408b154924[0] ;
            Iad3f7ae48f752d3ee71320875a2d1d170e879dd5ff51cdfd662241e6a30fca6d[0]  <=  I9288b2d29db5e8dbeef47da923a8ea2055a38ca1f37d4d8ed5d458408b154924[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2dacf26260c042fa148fa6c4e97bf878ad2e89e221acc0616141e1841b0c320f[0]        <=  I8e09e68977d9f7456b662b0d7fe4575c48ddf88f897bbda3545f7b1b63d89ccc[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8e09e68977d9f7456b662b0d7fe4575c48ddf88f897bbda3545f7b1b63d89ccc[0] + 1 :
                                             I8e09e68977d9f7456b662b0d7fe4575c48ddf88f897bbda3545f7b1b63d89ccc[0] ;
            I4e9c85ad6975994daf65df213a2d2fa5a6a2abd91e66d9c9a6f540caf4c2afe2[0]  <=  I8e09e68977d9f7456b662b0d7fe4575c48ddf88f897bbda3545f7b1b63d89ccc[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6cc3662b07a43d62f870bc24d55a9e5675a0e50d923f3b293d7004c2c62ad31b[0]        <=  I53ec51c004b0546b3dd0563e2c294a6c4b95b21301321aaf80c838931473cece[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I53ec51c004b0546b3dd0563e2c294a6c4b95b21301321aaf80c838931473cece[0] + 1 :
                                             I53ec51c004b0546b3dd0563e2c294a6c4b95b21301321aaf80c838931473cece[0] ;
            Ic8f9966a2711f4810086d09b86e16ccf0d31339d146ad5c38d34c973c757947d[0]  <=  I53ec51c004b0546b3dd0563e2c294a6c4b95b21301321aaf80c838931473cece[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I670beb5586ec69af20e65eeaa49be81826908f01db21d27643e2561621962b87[0]        <=  I3c0c87041c080ddc72a51a1b6a4fe12cbd62dd40515520e3924dd8cb63728a83[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I3c0c87041c080ddc72a51a1b6a4fe12cbd62dd40515520e3924dd8cb63728a83[0] + 1 :
                                             I3c0c87041c080ddc72a51a1b6a4fe12cbd62dd40515520e3924dd8cb63728a83[0] ;
            Ic1385b7aee4e3b643e13733b56157e3e92e638da28cd1234e275fc9263709f04[0]  <=  I3c0c87041c080ddc72a51a1b6a4fe12cbd62dd40515520e3924dd8cb63728a83[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I88ba583883fb596ad6cc6716008143d6b643816e8e694ea5f32ba95f3cfffe48[0]        <=  Id9bb31b77b580b8375e799bc74c4829818ee16c05c6dad069736736dafa7a8f7[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id9bb31b77b580b8375e799bc74c4829818ee16c05c6dad069736736dafa7a8f7[0] + 1 :
                                             Id9bb31b77b580b8375e799bc74c4829818ee16c05c6dad069736736dafa7a8f7[0] ;
            I3a173e6b224a6415ad442ae28a0af62756975427859bbcfc0af6c8e5effd62a6[0]  <=  Id9bb31b77b580b8375e799bc74c4829818ee16c05c6dad069736736dafa7a8f7[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia8545410ad46518007f6812cf6132f4f4482933818a0fe103dae14b1530518d7[0]        <=  I5800b2a82f1442915cabe6307e4eee8c6b4071bf852ca93d4a7420bd0e6b1e24[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I5800b2a82f1442915cabe6307e4eee8c6b4071bf852ca93d4a7420bd0e6b1e24[0] + 1 :
                                             I5800b2a82f1442915cabe6307e4eee8c6b4071bf852ca93d4a7420bd0e6b1e24[0] ;
            Ia5580120af4590da8aed890f81ca17929e4c998617df957686c095e891649c83[0]  <=  I5800b2a82f1442915cabe6307e4eee8c6b4071bf852ca93d4a7420bd0e6b1e24[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7018895fda9af57bf39b18e9edc144f8854067ef25800ef8eabe76015fc207b5[0]        <=  I40886d5f08de09dc76db805b27c8ca792ccded54cd12ba2e6b70c30121ad9f79[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I40886d5f08de09dc76db805b27c8ca792ccded54cd12ba2e6b70c30121ad9f79[0] + 1 :
                                             I40886d5f08de09dc76db805b27c8ca792ccded54cd12ba2e6b70c30121ad9f79[0] ;
            I58a3910d475757bccbde2da0e6b5dd5723cbe44e1f4d3e71ac2973fd2a03b3a8[0]  <=  I40886d5f08de09dc76db805b27c8ca792ccded54cd12ba2e6b70c30121ad9f79[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ib57f995d569a522f5562976385f777cd6cc39ed15491d0ad8f88cc0e908c326a[0]        <=  I0cd63486c66b03be7f8f629aa2577ef8849fa2408aa41a58514c75db95432892[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I0cd63486c66b03be7f8f629aa2577ef8849fa2408aa41a58514c75db95432892[0] + 1 :
                                             I0cd63486c66b03be7f8f629aa2577ef8849fa2408aa41a58514c75db95432892[0] ;
            I1b76b0f61e714e21a844e429806d641f6a24f0eb19c23a3c2fcfb76baaf3e72a[0]  <=  I0cd63486c66b03be7f8f629aa2577ef8849fa2408aa41a58514c75db95432892[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I35636bd5c56cd95d41880b5c936108a3ab7c1517a8e09f76731b2154d39c87f8[0]        <=  I8dc1d4da11f5cf2226f4d8211654acb056d8fa751da8aab85dc14664d72b21a5[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I8dc1d4da11f5cf2226f4d8211654acb056d8fa751da8aab85dc14664d72b21a5[0] + 1 :
                                             I8dc1d4da11f5cf2226f4d8211654acb056d8fa751da8aab85dc14664d72b21a5[0] ;
            If0211848e6cda136970069df5b6156d4ac213717491c68ed49ab39d2cffe9999[0]  <=  I8dc1d4da11f5cf2226f4d8211654acb056d8fa751da8aab85dc14664d72b21a5[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I84280195e0f72492aadcce8eda907d5de2e05dc16b9c5ba1fc2f345192ade355[0]        <=  Iaa67bf8b75feef8789908b65a38dd8124db04184092d5a584054726339440c63[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Iaa67bf8b75feef8789908b65a38dd8124db04184092d5a584054726339440c63[0] + 1 :
                                             Iaa67bf8b75feef8789908b65a38dd8124db04184092d5a584054726339440c63[0] ;
            Id23ae21f713f4f452abcb1c1839b5524c452bb8bb0b6c35683f9bde212bc5f96[0]  <=  Iaa67bf8b75feef8789908b65a38dd8124db04184092d5a584054726339440c63[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6532aae67414dd9e03b874fd4b6a321437892a7d89bab17ec2d5a684aa9ad55d[0]        <=  I845063b254fc4b71844ce1e01433e1d8ad7e176fc80530a73ecb26c31bcf8bf7[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I845063b254fc4b71844ce1e01433e1d8ad7e176fc80530a73ecb26c31bcf8bf7[0] + 1 :
                                             I845063b254fc4b71844ce1e01433e1d8ad7e176fc80530a73ecb26c31bcf8bf7[0] ;
            Id5bdb0f5a920710b1af7cc3abade245196df9d1ab4b7f26277fd93e1bbee5556[0]  <=  I845063b254fc4b71844ce1e01433e1d8ad7e176fc80530a73ecb26c31bcf8bf7[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I7032c41ce2651dbb03999e2120193d71ed608e40ac2d51329837f3abc0a976b9[0]        <=  I51b1e937ea9e8b9d8f3d8c8c66d7f69b172137911df42ee5fd10dfc5d32bca27[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I51b1e937ea9e8b9d8f3d8c8c66d7f69b172137911df42ee5fd10dfc5d32bca27[0] + 1 :
                                             I51b1e937ea9e8b9d8f3d8c8c66d7f69b172137911df42ee5fd10dfc5d32bca27[0] ;
            Ic72616171e7fb8489fa12cc29be1f74602ff8e4bd28ea085e938da615238a0fa[0]  <=  I51b1e937ea9e8b9d8f3d8c8c66d7f69b172137911df42ee5fd10dfc5d32bca27[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I9a800fae8c9498d12065155e7e781ba817ee2b03ea6540813400bbe438f4691c[0]        <=  Id90613f9d2194b97066ad1f5247ec5becce3f39f02d165502d84b92178a02948[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Id90613f9d2194b97066ad1f5247ec5becce3f39f02d165502d84b92178a02948[0] + 1 :
                                             Id90613f9d2194b97066ad1f5247ec5becce3f39f02d165502d84b92178a02948[0] ;
            Ia09db6bd7cba6c6e15cac4c6ad0d4c98235a7437beeabca1388fb1b4dece5d67[0]  <=  Id90613f9d2194b97066ad1f5247ec5becce3f39f02d165502d84b92178a02948[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I1dca7dc76f83994b077209eb2742069045e743b6eb763805cbddf87e6a8fcc34[0]        <=  I38b86f50ae5aadaad749bf30610fc173dbfebd9d3c9d91147b1b3afe8d7f1004[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I38b86f50ae5aadaad749bf30610fc173dbfebd9d3c9d91147b1b3afe8d7f1004[0] + 1 :
                                             I38b86f50ae5aadaad749bf30610fc173dbfebd9d3c9d91147b1b3afe8d7f1004[0] ;
            I15ab76f6e4824af9b3b4f5062e8dd3c426e1ff0c5f68e4733828c710eb7bca54[0]  <=  I38b86f50ae5aadaad749bf30610fc173dbfebd9d3c9d91147b1b3afe8d7f1004[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic16409f8fa42d6ac05643c3943352c03f19cfee0c3068e96d6ca3630b8f2cacf[0]        <=  I12d2f80160672a05ea5c1aa8b8b52b7ad7872b05584cd462f2fd449b06326ea8[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I12d2f80160672a05ea5c1aa8b8b52b7ad7872b05584cd462f2fd449b06326ea8[0] + 1 :
                                             I12d2f80160672a05ea5c1aa8b8b52b7ad7872b05584cd462f2fd449b06326ea8[0] ;
            I12b276cd6b0aa86ca2e28dbb1f4008ab140668e16e4ef96604a6d1741c7f2f95[0]  <=  I12d2f80160672a05ea5c1aa8b8b52b7ad7872b05584cd462f2fd449b06326ea8[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ic66f776d5d728142606f048e3cf27e927f094082fe1dd31f90e757beebd5b5e9[0]        <=  I08cb7d15d8198cd0c19dee6c97c2732b1f72f7e00294bcfb0887c25cb0951701[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I08cb7d15d8198cd0c19dee6c97c2732b1f72f7e00294bcfb0887c25cb0951701[0] + 1 :
                                             I08cb7d15d8198cd0c19dee6c97c2732b1f72f7e00294bcfb0887c25cb0951701[0] ;
            I01577c8c0e65ca47449450a8b2455ee84cf5c48bb26a0799b5523258a039ae40[0]  <=  I08cb7d15d8198cd0c19dee6c97c2732b1f72f7e00294bcfb0887c25cb0951701[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Icfe7c47d401f26676f3f8f13e34894792fff7a3881d754de5b4ac1130cfad989[0]        <=  Icf9ebe6aa27457ed3d8ac986d9dc8260bc590e8c778585764d6021c62b1f9d5b[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~Icf9ebe6aa27457ed3d8ac986d9dc8260bc590e8c778585764d6021c62b1f9d5b[0] + 1 :
                                             Icf9ebe6aa27457ed3d8ac986d9dc8260bc590e8c778585764d6021c62b1f9d5b[0] ;
            I63ba87cd2daa7c3c625d3ff5bdaca7f2115fc2d65e13972a22b2c2ae5b746d4a[0]  <=  Icf9ebe6aa27457ed3d8ac986d9dc8260bc590e8c778585764d6021c62b1f9d5b[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ia6852c630d3d698cbe47da7b990ed04d4e0b995b3d765ff6a8146da11e42dea9[0]        <=  If4d6db4bdc3cf9677389d183b78d9ce032dbeefbc9c6374296777d351a8d958a[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~If4d6db4bdc3cf9677389d183b78d9ce032dbeefbc9c6374296777d351a8d958a[0] + 1 :
                                             If4d6db4bdc3cf9677389d183b78d9ce032dbeefbc9c6374296777d351a8d958a[0] ;
            I576afeb6020cc0a8e35837b4b96968ed04cd444999558626adac849848fe7c6c[0]  <=  If4d6db4bdc3cf9677389d183b78d9ce032dbeefbc9c6374296777d351a8d958a[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I5e5d78a5f1d49833052eb3e84c516dea9f05d6d49879c593f5e0b9745f84fde7[0]        <=  I15ae50aec5944edbaef4ec461dfb5ab01f597a46233c643d7139247b8bc2f6c6[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I15ae50aec5944edbaef4ec461dfb5ab01f597a46233c643d7139247b8bc2f6c6[0] + 1 :
                                             I15ae50aec5944edbaef4ec461dfb5ab01f597a46233c643d7139247b8bc2f6c6[0] ;
            I3b8769ce28405c0bb978c458bd6272f10cea5338af4170ce4e93a8932ae8dcaf[0]  <=  I15ae50aec5944edbaef4ec461dfb5ab01f597a46233c643d7139247b8bc2f6c6[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I6454add174b2968c545e831c5bacd6b95b351b7d68448b3fa9c2e5476a8cca35[0]        <=  I6dc76307fe143582b214c945a6c0a35a4545c8bebb622615b3ff784edeb2d0b8[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I6dc76307fe143582b214c945a6c0a35a4545c8bebb622615b3ff784edeb2d0b8[0] + 1 :
                                             I6dc76307fe143582b214c945a6c0a35a4545c8bebb622615b3ff784edeb2d0b8[0] ;
            Ib4638612fcabc0a2c2f2bba5a2b9eb71cdea23575641b3f81fb6220fcaf284f4[0]  <=  I6dc76307fe143582b214c945a6c0a35a4545c8bebb622615b3ff784edeb2d0b8[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            Ie062df11427db764a0e09705579e134d08f4ed2a027e913a43495db5d5fb9051[0]        <=  I831951ac212604dca0a254f80af9c1bc9a941f743abf321cc91063922eabd175[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I831951ac212604dca0a254f80af9c1bc9a941f743abf321cc91063922eabd175[0] + 1 :
                                             I831951ac212604dca0a254f80af9c1bc9a941f743abf321cc91063922eabd175[0] ;
            I16ea389c88e4591f7686eae3f1988dd5361bf893895697c0ade8627986a9fc5e[0]  <=  I831951ac212604dca0a254f80af9c1bc9a941f743abf321cc91063922eabd175[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I2a2245385398379002074dfa174bde148f97bb3bd83073505b550c0c0bbd1e65[0]        <=  I0d347b21cb8cd8b8a0fb2e002b97a2078bbdf1c6e71a0e4b9cb022e2a0db8de3[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I0d347b21cb8cd8b8a0fb2e002b97a2078bbdf1c6e71a0e4b9cb022e2a0db8de3[0] + 1 :
                                             I0d347b21cb8cd8b8a0fb2e002b97a2078bbdf1c6e71a0e4b9cb022e2a0db8de3[0] ;
            Ia17edf214ab782c25bbab97f6bb4e04b2fc46d41f9a97fcf617418d54ab76a7e[0]  <=  I0d347b21cb8cd8b8a0fb2e002b97a2078bbdf1c6e71a0e4b9cb022e2a0db8de3[0][MAX_SUM_WDTH_LONG-1] ;
           end
           if (Ib46a5934f2d38e6813d46ec1b5be874d1f79ab6b3193199e03e39761d9af3a0b) begin
            I862f2564a9e7f99bc8370fe12c1a5e57612d564f1606a21f6a468d558c23fc5b[0]        <=  I9c8cc6c27c1fe245ae54ee4a9dbe2f5fabe4c675abb8af6a49a61e6076233e73[0][MAX_SUM_WDTH_LONG-1] ?
                                             ~I9c8cc6c27c1fe245ae54ee4a9dbe2f5fabe4c675abb8af6a49a61e6076233e73[0] + 1 :
                                             I9c8cc6c27c1fe245ae54ee4a9dbe2f5fabe4c675abb8af6a49a61e6076233e73[0] ;
            Ibcfba9f1fb81d976955a1fa7101f0b0db16c344c82cc5ce81f50dd3aa2928d37[0]  <=  I9c8cc6c27c1fe245ae54ee4a9dbe2f5fabe4c675abb8af6a49a61e6076233e73[0][MAX_SUM_WDTH_LONG-1] ;
           end
       end

   end

assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[0]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I96fb06aca6108479f7e21e1835a091a9060c2925cc6320c8ed71a0a0092bdeab +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[1]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Ie000dee1e3953811fe9424588b71a7dbc88f41ec69afd16e17e8fabf141c31ec +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[2]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Ie873b138e19cd7f7e8afa8bd8f8c4610b65d0fcd647e76d880d25f6fe36c54ef +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[3]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I8ab1772a3bc752331b0bf62069643cadb48bc13bbb06ad3eddc68ac603d73654 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[4]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I4bce49360270b653e45b914c493ca8e5b74beb0b6b85838bb3b54f1f39389fe3 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[5]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Ibb4ff9ffdb2771ff640bf958798f8447a0dbcf15ed0ef9f82068826ec621de77 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[6]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Ia4691d32d9e84827a250e0b3d6ea8142c24c9df4ade01c19583e6cfca06cd990 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[7]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I3a1380b85cc7f797ff92d02b7081d1ec3ba069aac74162ca059c399daa10690d +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[8]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I14919dedf2b4d4caae8efa1726435d1946f48e1e9b1052133bebe8affeb3556d +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[9]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I852a201bdaecd968b6f9c9b6bd64dc8035a17fb92ffc806a690781666354b069 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[10]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I345c0aef41ee2863a96a076a78d92c7498f50ef90e82e75565df1d1f38a08161 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[11]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Ifb94a220081758ce91634fef64be084898a662f7c0e8cc9f86859bf3852b3efe +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[12]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I5f1b294a0702ab37f94304ae67fe91abc04c397dd682d371126a7ceacf7c43ec +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[13]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I81aa911c9f6f4bd88314aa3c5310efef6c40219ca93521bbea3c1afcea7bb48f +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[14]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I97f674eaee005fc7a54ccb648f5a0a67cec041e895d62eacbcc9a37068b912a7 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[15]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I7628fd0a5ee3ec547c1b4798a4d76de651807424cd18f0b3b8a3bea849e6fe0d +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[16]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I1d8a992801d3f6a457848578ce286b496d4e2a69937344bdcbab4e8b1af1fe4e +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[17]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Ia28f68b737aaaaa6b98aa5e9696b937e564754edef217740c414c16fe2e485b6 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[18]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I099e314496f03784e5504a35292defa79dc063aa81e6aa8764802f7fe3a47114 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[19]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Id4bcb557769f043a7275ab01d6d9794d4cbbd9309be38f58acc307a1e693f347 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[20]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~Id1bb830ea0f92a1c0ed0addc915fc85198e4744c4bf7369b4ee1f7131f5f8542 +1;
assign I72f7d0f07e7879c5e77bcb27964b5ca3d3a2afc4df135e64cd081608b37a8dbe[21]      = I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75 +  ~I31009872a3e84f78bbf1f12a7da708c45e3b708bd943b6f4561ad436164b12d8 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[0]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Idd9957e5b52c4d33e24910559d8203415afdf467bbe1c9de950145282c7eacf0 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[1]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I6a09910e62aa0cf665f69be80c9ad61f2d31115012314b8188cf79fae365626c +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[2]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I3d6f6b104bd2ffb35ea6782748bb777ec7eceae47ef2e1d18d37d1677d56cb80 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[3]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Id5055b759fe480d476c4bf08c420a5dafe9e65cb03c6d6991c1d225af0a51d7b +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[4]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I93e543ef3d58bc8bd48a279299dadae1d7f4528c3d09d7106b969e15565d3a15 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[5]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ib6ff050679c6366efde7b9809fcf42051f107c18863bcea79d41b5fee0603e9c +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[6]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Iba81256fd46cc69f1367fc6ed7b712d2695e099c52b476f9b39f0a13404dceaa +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[7]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I608b794037b45c46a29ea01e378b63a1f267c4b489b0866fe2f6090936fa9d44 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[8]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ic48347f5264e8e479996a8dba0171a108b602be1e1d24b2fcb43cd2bdb82f61d +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[9]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ib62b5b3c80d193b97bd6b5c0d5678e424026381949c3f24546d367df930cbcae +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[10]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ia7900b5a01cfc1c4db79ca653f072956c13e2040cbd94cf07de2f1d969222fa8 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[11]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I1aa136009f34c39a8dbc39b4444642cd09c9cd2f01bd6310287d4ddc9bedad85 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[12]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ic195e053a186bcb0e653c0ddec75c57d1b3210c583162dd90978858c98fa53f2 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[13]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ic859d34db6baa83e73a8627c251c877e93f15653973d0634c42a8ffc9f628bae +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[14]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ibeb23788ce301c724494a2852312b38344c27416a5604c0145fa330ccd1f290d +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[15]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I5ccf8e87b0b8e8ce9bdf4b3329e4458a628f2568184f82b998ac62ea28bc0307 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[16]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Iaea7277e745e05f803325e0f19dbc5a54234878a9a3cb2cedcc013e3942e9cc0 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[17]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ic94e7c887d7f24b573b470820c36fe8a0fef750e2c46675f8867d78f2100f1f9 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[18]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ifa0b8243f5ab6adb88a70fc1245e3480ea3fb3f3af846fdefd0613ca91d7b122 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[19]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~Ia00cd24df6e6b22b466e1492500f1948b3ba3d70bdca407d1c22b4dfaf374eb7 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[20]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I8b41f817a4008df0994e2efa6b33eb847e82b031082f90a767467ffc03cfdb93 +1;
assign I2d1d71329abe9d76c75b65d1cfc8efd3b92d68cab8c97c3553ea62472faba3dd[21]      = Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6 +  ~I8d91c857f2c8154bb09d456ff73ebdf81e3b7d9bd1c57c2e6b8c2de74e55cf48 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[0]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~Id0f930aa222bd91b8a7d5f80a38d84993a63fa1c6aca3d37ed259294e08869d8 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[1]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I58598429d44ad951f91139a213d3b0bdacac6d71f1b9753886dfe1d39d0024ac +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[2]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I3cca3cf08c967f80e7e255a590bb9c442abc535cd529f7ff304f25d5519dab04 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[3]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I42d1b7202048c81ca3a8bba0dbbce65501cb7a519fde37085c68d01db7edd635 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[4]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I07bdf8f629cfc9c094023be167a717880dc3a42099b01bffb431036521cd6019 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[5]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~Ifaa925832248fd0e2f5841096d9618c2fdaa3c63a3130b57f493782f96473088 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[6]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I2c22aed0ed8abb0cb8906a35a4d44cfd7cc68b2924e474680a2eb6cf7caf5582 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[7]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I31ca3705bdc7e063c61023d93193b3ced40cf440afd817d0d730f6c8d37f8b92 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[8]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I789461a909fa4abaf3840dfca4f63bfa63fdab389e149fddb7d8ae2b876dc912 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[9]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I6ff3298d93471156b56cfbbea17c8dc0405bfe8654e9f830bb33bc6c9a649b3e +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[10]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I9eb30c75f8d71ade925633d7c8bc6b948ae519cdff33ddb885761bf72a8b0869 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[11]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I5456c559bdce4d65af540e4c71c19e44227c62e5c129b7de968ac7f311dd76f4 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[12]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I98e4b84e98742d38b206ac059ad123966ee63903c616b9c31b4ba9615edb9f40 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[13]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I40d7eae63827c6efe2ac480c8eb9f8a8f77bbfa845caae02d137397c9da822a9 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[14]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I30a9d5330fac5c3ec7b63cfab0edcef0eda61dddb23d2aabf733b9982c12b4ad +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[15]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~Icbdf29918b91006ffdc8b68c707840ee6bb9c27779dabd372e2033888743409f +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[16]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I7f6b89a61d6313029102fc48e92a54ffdece30e9eac1191d840c488be69d8223 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[17]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I9471414594b824d60836981bf4b9931c135520ad1ae7dea177e0bc591c2572c2 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[18]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I0e9135a0817e96971dc8c4fe6eec717a563c44738f7e38d5bfb2f4dda8c77876 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[19]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I0847713503570d7ab3efee12577ba27aa81869a22b14ec8a244fbd4665d566f4 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[20]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I7b529f16d1499766369f75cde5a356cb12c06d21f42a10932edc6d54146735a0 +1;
assign I437a80b5f5d16324e086f21cde91b88bf11bc4fee1b943d83a425ef259fd3a86[21]      = I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee +  ~I1b93b1b2c5f55e2267a4deb4f75ca91039d6893af8e082ea85b7a5e9354117e6 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[0]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I7200758287b0c7ed92552ced989756e1d49b5418181b9e36421da7e2694ed3a2 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[1]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I96e7a523360a0cc0f3abfea09a566658e5e9f3316c3c412f99fd6340d1b64235 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[2]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Ic4839247bb24d460ee6d963d31fc390e8d9d679cd73f058d94ec34a18ceb39c0 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[3]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I23ef4f4232fa0d8813a25ddca38a2745fb660c05dbe9ddc2cc33c47d45b3fecf +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[4]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Id5e78e4ed6db0562ed51d1da1f34242f54def8255088c3a1ccf0221ee8fa153f +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[5]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I17cdc222663e370d6ef2539ad03c45a7949d9606583c17568a24c528a3e8c12f +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[6]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I65e452247faa2c9d6b01dcbbebd5e8c31884c88e70dc8ec76d55aac7e77e2d46 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[7]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Ib0641eb8fe554f69ebb57e8e900f995c07bddadffd25c01781ba234b87af4a94 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[8]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Iee9c2c6a9b8e84402eb1e0de611c1cb8ae1e802226f2c07833bafaba74f1ac15 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[9]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I443435c78145236b927711299e8bedd0d29a743e3784ac22f70b2284b6be11c1 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[10]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I4a86387a3136768ab52d320fae7fe63c7c74bb5541d18889faa263c71b2bfce6 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[11]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Ia0c4bcb29e2939b889fb7a5a7b62b49a3eeb3ee6f4555518c9059cb34dfebc7a +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[12]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I3de9fbe37d08009f5fa66bf7c59debe7da836dc078e212968afdc608b100e3bd +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[13]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I7c6d90cd79e1b85ce9a5452570cfeec8faf9ce3e6bc886f66495ec2a66fc8c7e +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[14]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I57d80f41498f8d7b91410dc02e646a45a3f05d45e9b5871ae95d6432ecd2af56 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[15]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Ief90cf0b0997823c3071eb46b636e384077579beae3d85d29e639a7719763396 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[16]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I295d7aef060ca978805bdf65138e5bf134551eda9c396a22165a77a3091dfd28 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[17]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I73a855a590363c762c34008e77f73f961950c0dd71b795acab3adf40c4540453 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[18]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~Ie38c638da580ca7d25fc0754497163d0369f31a6cdb4bd26663a759b74efd588 +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[19]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I2c635a0b11af3be4774428af79ff5cbe6a32ede6ad03ac197ecbb3ca2ba78f8f +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[20]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I34a89a8aa68b1657dc7137437574877b170659ebdbcc93a772989e2b8b5be31f +1;
assign Ie7b77a6994898104117c58bc634f3e85a3969669f097fc26118efdc65814258b[21]      = Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493 +  ~I9f9d895211b42c2c9d491349dbe7aafbad775942920197105c34837dba6563a0 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[0]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I11c6d693bd6c019722571e1aa6eea0507f351a89cfc6d16f8fc51997981aea81 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[1]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~Ib53bac100fd49f57a5185ff4ad973dfe8eaef6de1937bb32d9246dae9459442b +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[2]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I7ce5fe43a760b5a43815388233952e1bfe5d8b5a7c002f26ae2d462129aad434 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[3]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I3a2c9aabb8b064f82bd6f6571bdebdd704abb7526f4977a7b98613f883fdc62a +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[4]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I52f4d169be660862052b60924958cc9a0eb99b1454608fc48d47192452f8b390 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[5]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~Iade009d6c5b9e00f5459c53b0c254dda356081e6965366db7b7ac42a992e3ae7 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[6]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I52dd625c97050874c15b1980a389843c4a7a890d73f6efb003c4324c029772aa +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[7]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I11bf8ca77f64484279bd3f36febe1c6869fb79b4585a800449a0e5c683c6aa18 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[8]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I255a6c7b69c31d60711a86b1f0da51040ab60c48952002406e028a200a835049 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[9]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I24bc395a7644f2a2d7702656737c32662f8c2e8a7e2b2d4c1bca200dcdf49219 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[10]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~Ia84166c5479fb08b9d5bafbf3446230d231e77cb1a3034b53477e2f0632ca74a +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[11]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I544bba815490c8592dda0fd85cb612828256c09ba1431bc2632b74cc9cd2aa29 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[12]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I7b8225b7ff4972426858a8550dc67a231d85fe94426bf0812906f1aee0e2d097 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[13]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I3358739f5e55263208e661a339d6b29f188f07ef07e2ee7a63a24011a4f8568f +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[14]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I5eff39d324b6a8910fad41786d651086c622d331987e649ba4b3baae11ca40ce +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[15]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I4a5c4f290852b8c1baa90ae00400045825f13c24b546dc4a7848f91824185f7c +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[16]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I9af65d3592633577409561b2069e30c73196d1a4798cb92f4d2f14db8771895c +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[17]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~Ie2261f6d4e2c2ce04997cd365593486e02a7d85106b9c3b568ccdfcda7a9c352 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[18]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~Icf0b2747a9e17f2d2672f7a17111c6bf54bed7d8fedcb5260f25fdc4280ae727 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[19]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~Ifb6bf654293ed3bacd2a4ffc883b8ca5e4dedea39e338bd1a30b21e8f8df2f62 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[20]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I0f4ede6017039c42f04051822cfc539cbcacd77427efe92d393ade1c10a46462 +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[21]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I23e0423ae4012d108a4e6a495814e0e6f920fa6dcab900bb35cba7b95f590c9b +1;
assign Ic0597480f1b25983453c2c9444467d40b143d832c9115cea4ad437cc2999642d[22]      = I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac +  ~I571233769cc63838bcc3d61e7a5e95805c3f4116c0053dfe86831eafff7c32fe +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[0]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I7fbf7b7f7a1f0155cb188ee4219620cb35a2fcf98d2687cddfa2508273b70154 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[1]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I4f56f225d6fa40e0469f803c2f72ca27e9c45768ad2af9af9ad10e529e249aa0 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[2]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I634dc6f7c843c6e4c63ce6a21b9cd7a386600d1155c0696988403fc1ab790217 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[3]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Ieedfb1902d1f76f95f5f971b578c2440fa5de47dd78e9dc70c35698f813048cb +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[4]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I88272c473a90efa576a83d0c277090f5814599e5aa192b878cde74215909c46b +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[5]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Ia3e877a9f66cb7582b125e56b7c3f79601eb8e700f54e14f967a4d9df9b5725d +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[6]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Ie278ca9a470ffe4ac78bc335aec472b66707cf02bd91256aff2e7c73b5d2c6b6 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[7]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I5ef535b2e573d96fd518cbd837132928a2a0c6a25d4eb3c360f1cc0aed89656c +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[8]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Ic486b9953b158eae95a2d8914f8144e669e056675946d245c8239bfc249a16ac +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[9]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Id89c8a47964d1e4aa4bb9e96a79092cf7fb55eee5808d6323ecbdecf8926adcd +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[10]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Id1e80f29821e7ae727d759f44b21e84843025c938468caf7c8adfba52f1cae43 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[11]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I7530c712ec14c8fe97d1699177ef642847c5c1ce6185d1eab39b8416b562b454 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[12]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I41b365f8c613bf86dc5e2ed41719ec6823046127babf87a083503ebcfd38ae75 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[13]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~If9bd4d7f3740f15bdf597de00eecf1cbf2e3b4efdbacbbad889c0946a6b34a24 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[14]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I31c470f2adda0a23b85c3245646a168f2478bfdff11a434c1455be20db703c64 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[15]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I9fa9c98579041b6735eb78f7b3727824dd61991c6a6d91a158c6ac65cb20b05d +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[16]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I9fc6fbd6f2f888b9750fa59a966971aa6ba6fe4eee8c8f3ed4c3ea60141a7d23 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[17]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I8c133563a8b5e359a6a45a7f3b4e939fc84766f9fa09634d18e5d2101d0c0645 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[18]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I84238bd7e53e0dd7ba07efd813661c8cd1648b76c44665dfe51fd07dfaa9b249 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[19]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I6c3a9695a1c1d22809b1378e82cbdbebc1ca78428194df50cce0a69d6a159398 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[20]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I4d032ff7482be75de7d2b816ddb2bebfa9e896e45fdade2b5f81b35c003a59ac +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[21]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~I6b4d2a32c92c22b1cfe81ee6620c69af1850621deea406d75f098da0542843e8 +1;
assign I061b92250e8f4b07f7490d2d8cf732e80ab3137330e3727a22f0642dbc515ad5[22]      = If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d +  ~Ia0964979ac559942d1da1c41ecb3d9e94c6c7c0da3d16177cf2379db8f37aa65 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[0]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I236cce67d0aea9f9c8d5ea3c39cb598d55f734b44ad6e3972e7f6b91d56001fe +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[1]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Iceb8741c9680982b02ba9fa2dd76d3b45155ca5f688b70c41d66f3b3690dce42 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[2]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Iac9f4a2fa823ae63e73b655020376580991cd4b2b3123204a757afeefe35a10f +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[3]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Ifb57457918458a6aa9c5df68dbb83243fbc49b3b7037575f43749dfe1bef373a +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[4]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I91589fd8a2ab91f079bb41631c44926b2c6f83b82448d758d97578c314d0b76c +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[5]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Ic20b5a20229313d70c01a5f53e13e96095c1d8695144668e66efdc81efdd8374 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[6]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I53e90d4a2bbfaffcf92f2e9fd80c491e61990aa575337df13d24211a558315a0 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[7]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Ie57b3acbbf1d1593e02ad38bc0e07bb84db2655f9282adb3ac5edc311e882641 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[8]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I632095e999af63661b01bfe8bad0078cfc2e74217253d3971230968c235bc526 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[9]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I6a66a98136fb7fe52fd830d869dc53a3855a545aedc1d16927f76bc12e319060 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[10]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Ifea15bb5031583fe42f92f554866179105e46b1eac3c6b691958a998c26ac2da +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[11]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I8b2c2b27add863ad56639a306f803b656ee8f91170e649d29aedc5321181f857 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[12]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Ie3290070e785df28e64ff4df124d14c370c9edb924d5f35b059a6c82e8373f91 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[13]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I02ed3128371185efeae1e27046aa378006ec78d7c458dcba137f69c29c4363bc +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[14]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I8dcb7a5498da4a9d3e4a76923e84c88a30ec174503cd435864a066ff0ff464ba +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[15]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I94024b61447a332a2c36a75bbf305f3fd80606bfbfcc4ee8c5783e3910e9840b +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[16]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~Ibcddbd4e851466c5ff49f13244c2478ab6c089e6d8ad294cdfbdc8451ac6a895 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[17]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I50ff347e89fb452beb071f112e4a51e074cb3d66bd903552db23c17670286e7b +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[18]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I8b5ee5d271abdbdc518ce02f900da21e858d3e2530585fd859690a1a71502434 +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[19]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I54e64fd01d9aff7ddfc4babeff6703891da38578bb141d250c4ef5949d818cfb +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[20]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I448065f71638c5abddd1eba1fcf567566281d5b4b23ec4ff2d2208d32a506fbf +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[21]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I6ed6ee11f6983e96e7ccc4e4be6ed8c4ed166ca9075b9cd218f26f018ad2140f +1;
assign I34b3868f00019200d860d678e890c83dd4d2e08c2a746cd48665b55d1fd91308[22]      = Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e +  ~I0678dba3dc1a3400ab26e223257bf71c03f0e8d284810653b5e507fe964427f4 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[0]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~If34d8ceb2732716c923a7f250495970948ae431d5f1e0a025618c1070940ec39 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[1]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I60014273d45dd5019a1b82bdc0a65e44d9a16368d996c8c9ff312fe27e236171 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[2]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~If16869134ec7e59b567e29a1125f0d27eff7a3c612240e25462e2ee84a7e0104 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[3]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I8d95c0be0c84d3ee590f8e77065a6ef224e0a75b50aeadea980f9ef4b8d25001 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[4]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I28940d6e8fc5937055f8f50c0d65ac9fd892bdc9f0f2a571808f930c8ad21717 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[5]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Ifbf3cda7e0639ad343a64c5b3d2f45017f1d280bf72c96520cbf272104c90ad9 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[6]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I4aabce2cc01e829bb9c3d6a984cf2b5bf9230cf3913db788c47a932ddf71b869 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[7]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Ic9dc8459f6cd65f223a6386c82f754469ef74fbab59ded4fd1370fb69136c847 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[8]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Ib22de4dadb6e63ea49c52cd8bc86dadfd7b73a002dd8e726a9cf1b7b299a8c46 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[9]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Id6c8c2ebab66fb903f108466c8d15060ed1328fe9a979858569c39069bf050c7 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[10]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I385f4177f3a22b6fa4a6352d164c7d54c94b980806080c51d00a65f030966110 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[11]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Ibcf016cc83d0fcc2c731aa53147c199b32b3dc7a9f1a255e1a0e31615077205f +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[12]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I7e7be31550be1cacb2acdb27d5120769dd7a0a49efb833051ceb83c8cf691e21 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[13]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I26d08096b43367ba37b8f6dcd919bf4ecb9c660a39f2c0ae29f655e42b88887a +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[14]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I2c200a5ade27683d4afd55e06371f9880a7bb99259e2ccda5c368fe46bb385bd +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[15]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I92d28f6c97dab90de260df37f619e0a9000db48e278327a5c5d1528a34bb6dd2 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[16]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Ib053c04dd4e330e6784846706317bb6c8b12f9b36a57ee12807bff7de8ba7f0c +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[17]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I0f71479f871309f1717e7a1a2372ebfff4623c315cc31914588df3896740a074 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[18]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~If49d6a59c1d539e369406ee4e8a2ebb30199f46c335584e62921f98fd811001d +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[19]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I051f072f564eefd657cb4d59c1c851b56df2e70861d875f3b4c9b95e8945db08 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[20]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~Ifc8302f040679d23faab1ed8387a8a3aec85aba86ba9a78d3ca903126266af4e +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[21]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I2747ce9b7349ed89e3265df62bb0d0e612706d8c1b61e30a2878094662da8ff1 +1;
assign I2a4de2c850d1a5eedf0c9fba85c3c801fa74d3cc0d590b033b5e3e8e4e1a0a5e[22]      = If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c +  ~I3619e836fee4be75d6700a0e72e84df3a5a61003227363b8c4d348b8353075e0 +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[0]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~Id658b37d70ac8e3a324133f475a77c7948231571aa66ea0dd11b6460fca011a3 +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[1]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I737ae96fe290087c8ae686b90b2ac94df2185f7ad8b4252a6ec850278ba5ea9d +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[2]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I18777be7a1745485d18289e0b4a6e43e8a2e6758be0967b8cea04a3b0faf973f +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[3]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I1c30d2957a73fc51bb7044b869e28e0a8f6e0378a6098ee5e244efb43ab6a690 +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[4]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I69f7964c2f630ef03f49c2a6cac12420e0998397470245e6afaed2546b33775c +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[5]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I6f63c71eab6c2d7e3eb41fd78c9e18d6362d2dd4100c72b43d3e4b9d06663165 +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[6]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I23c91b29deaa2df1f4d96e343f6fb852a2b594937a4f62dc4be1fcbe0347c439 +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[7]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I8411087f9f6fa41d454a74dc89e5152e5e8edfa501c8753bd0735cec3789f14b +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[8]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I119a98150511650722429eab31b5785e99128641bad59a3cb31e42158a648c48 +1;
assign Ib801a0abc10b09b17f39a16844603b6eafe0cdc390325b728d8f9ddef2d5baba[9]      = I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7 +  ~I28a2b1ada19dc69ebe4949a75633b2f543159d2d1cc169f3bb6070c1419878e0 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[0]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~Ibbbf3f4aa7f74c37a0e8ac8a675ac9a9fec748ac720e6a78e9cf937dd089b8e3 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[1]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~I59a4b1b33d114a1b5bdd708e1f856f4bf729c6b86a4064967ca1faf779189164 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[2]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~I9b13cfb3566db96edc7c018b88f158faa57e4db029e3982290989c6fc08163b2 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[3]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~I8a1ba53134dcd1141a6f03dbed0f18ff7be9728dd9a6d6b138ff266c5307ba24 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[4]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~Ifd2ca31ff3eec501f34892055a36979681d27574ed8007e4df5cc0109b71bd89 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[5]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~I6b2620e847ea73b8618ac7bdcd8236c4278de3bef0bf1511ee9779306438fa38 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[6]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~Id2cf59876d070e0f34ee834d2691f7fbdb039bc9273329e2ce8eddfe736f0a45 +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[7]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~Iae213c2ac7729f8efe23deca256bf56f030403ef6ac00a3bc181414b6a3aa75e +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[8]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~I08e50de7e2aae48cc03a9959d08cab30d3c1c2ba8c4ef0799645787b0c09473c +1;
assign I49eaa0b83c0670e3c2f65b3306309a805f6d7448c9e6eb8d4b36b046e5cd2d24[9]      = Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975 +  ~Ibf22dd3f14f19c3fc769966f72e8ec980dc79c2991f69d03ca2defb7f720f880 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[0]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~Ibdd37577b403da9aa72ec3f4707379b1151c0b15edbfc4fd304c4e35c1672da6 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[1]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I8e23f89e84e219d5351bdfd4aab58f61c1cb310cc731164c6e0dd2eac37b07af +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[2]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I3baaba73f51f47e6a3f2310f692de9f7b9a871c65605e14d204d6965153ff4f0 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[3]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I82d316ed1475017844ea73f32085b755d17c9fdafd8191df2e363496e1950869 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[4]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~Id9e3ea08b52843b4a9426b735967bd4ac3d49bd67ab8fc85688b0f55e6df186a +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[5]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I77e34c24ea46e99b6bfc0f960d428d6ba3ea4f9261d5a183d83c386f259ab431 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[6]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I930ad334ce972f0b5dbddf698f6101a196d8072e90d8144b31ce3f4b48a73e59 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[7]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I4c0096e7bbf30db97520f824e05dbc28e6d1db344202349993fc68cbc95d6585 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[8]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~I75c796f56576dfba821e867b0de1a871ef35851371c3aa422532bd287f02ee11 +1;
assign Iae754c2901ee4c433c13177581d9ebab0bf346b31680a855929e9a319f615e43[9]      = I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948 +  ~Ieee1d2436dbda6f58f19df70b691a4ff28d37db8ccc12e04413e45f80d7124e0 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[0]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~I65b0824920910c82c7d677c2dcf4216e86940b3edc0b3da85d8f65505f58ad48 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[1]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~I169d92aaa7eb4f8516e38745955b91d8f6e0ff43cb212186293bb78884282978 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[2]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~I492e47d35231729b266a9f31aba61a3ac2c93a9786a20f6a152d342cd1d0b911 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[3]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~I2624a2d841eeb09774127e5d709364f803826266b46f0fc3122fcdcf0aa129e6 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[4]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~Ia6414b3aff6031e10856953f6b15ffdb0971aeb680d784a7199386be15624ff6 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[5]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~Iaf94ae58c1d9c9206d02651cd03cf2e02bba505f76b849158530a38382396ffa +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[6]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~Ia0a40c2a77389cda4a8333aeaecf37a2595fbda87854a43162ad1299544bd9e6 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[7]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~If692b993dc571ec401ce86f38a18ea4f96a797b00c04699ce83ce875b7c31730 +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[8]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~Id5a74d0be90678a7b69691c10e4ab75b47914e213e67eae2f20d4b58e8a8d9ac +1;
assign Ibfbaa1c9c7233bd157bf60566e8dafec44bbf5dc9a8f0bf459a69b9f1e227c78[9]      = I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f +  ~I47b54f01ac82a9eb80a681633a06c4e1d432d358091e9d079f74484f40ab3e09 +1;
assign Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[0]      = I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85 +  ~I6201d3c2d85bffa03f368b5862fba1b2e0ce3735fcc8711cb8107adf16ccdeb9 +1;
assign Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[1]      = I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85 +  ~Ifcc25cd8dc442c6720ac0f764b432530aa63681953d8ba16b441892ff5966bfa +1;
assign Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[2]      = I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85 +  ~I256cb35fd6d4e6c6e1c1a9b42dcbc307f858e5f9525acee9fa7af42c820664f2 +1;
assign Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[3]      = I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85 +  ~I67183da8c2763243a285b7cd41d838337f98eb6e59feaaa0a9150bcd6c29877b +1;
assign Ib3c8ff1cf0daa408bf3966437b1b52d059a5a685fdef802597a79d14e7ef37e4[4]      = I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85 +  ~I730fa6d01ade8f1439b29b955c5cff62700a90e523a4f4208ca2f9978e59afcd +1;
assign Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[0]      = I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd +  ~I37084afdf6695d3b8fb0530643c8b03deb2499f4f68ead04e3b5b79aa4467f73 +1;
assign Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[1]      = I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd +  ~Iee510842ece3717ba6eefc3ccd844e97a9718788683d4c7ceaefa6ca0030585b +1;
assign Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[2]      = I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd +  ~I53d3de58d6308b770e4a8884447a5f0b92931c8d83c62c86714b6e539b498894 +1;
assign Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[3]      = I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd +  ~I1e8142c7ece070c02ed90211fbeb423bc2a4ab19fae011793be99c68ff103705 +1;
assign Ifb23b085bb1c5f0456cad8d85841933550057b6e834945d41edfb611b614241f[4]      = I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd +  ~I425913b12fc3c865d95f1caead00d8c49de08765b634aa444243f4a03a53d0df +1;
assign Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[0]      = Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03 +  ~Ibe0fac26b5e106fc1753aeb842e8a04067fc91c95e358b1caa58db8192381837 +1;
assign Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[1]      = Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03 +  ~Ibadfd4f0852067e83ba6f0d57699585ae20eb542d1ad8f2cce3bda0d043ff2e0 +1;
assign Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[2]      = Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03 +  ~Ife27bd449bf6acad3f06d6e337bfc29c612ba6b3f06927e6f9699ab24d1e836e +1;
assign Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[3]      = Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03 +  ~Ie130bec82505842b184f5dd86865ab095110bc65e59662767e152f427dd7462c +1;
assign Idc979d57521c293e4359a88586d474b209e740a9304f4ea296f27a8f7763c08d[4]      = Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03 +  ~I2abc1178fa35959d8eb41342a7d7289e29054439c7bc06adc61f3a1d2e55bd6f +1;
assign I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[0]      = Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e +  ~Id27dfca888552262f492b81fd23b881938f66eb15f7ab21afb210fc6056fa09f +1;
assign I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[1]      = Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e +  ~Ia96c921ce4e0590c903d02dc69790c6af52898da90f4766121fa7b31e0ce6190 +1;
assign I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[2]      = Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e +  ~Idf239af48228dc01198fdd7240b8282cf247cbc6969403dd994aeac0e5f81898 +1;
assign I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[3]      = Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e +  ~I6687de5f8cb258492154a67fd3a3d5ee88d97a4db1c6c273ad158d5205ae3b48 +1;
assign I54a796ce62a764ac810b48aeddd21f65ed4b966d26b7d68a838c462b85d08f02[4]      = Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e +  ~Ib924c4eaf872874debc3b6ee65921f0381331e1421cbfc3bd17e8caf273049cb +1;
assign I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[0]      = I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5 +  ~If53d34fa90e564a24f6e116baa8a7934ec4c51c5f0bce8160f0f389391792fe9 +1;
assign I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[1]      = I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5 +  ~If0fe01f34db565bf669e2df82579abb4d3629e8bb001bbf874b9b76f8f780a37 +1;
assign I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[2]      = I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5 +  ~I61f7e06790f5516eba113bb79388fb515faa1b3a3bf06598a07f534ce2845618 +1;
assign I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[3]      = I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5 +  ~Id6b81456b5d3050b4e1fe80ccc8f992cf56eb0f08a1d29ec1e7cabe1baeb0872 +1;
assign I9ead67c6c06b3a745eb43ce8e7930b2330d9edf647ae990150985bd7ebbb3e4e[4]      = I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5 +  ~Iaa0b6d0f2fe24db548975f410ac5b79f687b7646169247f3891ce9e4644ee0fa +1;
assign I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[0]      = I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c +  ~I45ade5cafdcd254cc640ea8725da6961717fd6c50f747242aab6976ace4e8f10 +1;
assign I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[1]      = I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c +  ~Ie2e727d2073eda2be7642a6a2937cd3c4e553d8bb6ec56d914231b5bfb12405b +1;
assign I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[2]      = I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c +  ~I1aadd9b378df1ab58a1b1af097539d1407636833d9c2d8b08c8f70be326fe199 +1;
assign I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[3]      = I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c +  ~If83264f9ff9f7b77429559aff8b14fce54040210c6ba3476b77824c28b95bea9 +1;
assign I5c888504c3a7151c09b930f7cc0be203e201b0bcfb2508acd13c6f721ed26460[4]      = I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c +  ~I1cf0e3016bbd2d8e5debffedb198273a2d019ce75f2f8352a285d17264d262f0 +1;
assign I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[0]      = I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55 +  ~If9628510f239b2275efec7ce187b8eb7360beb042a425934ac81632815361368 +1;
assign I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[1]      = I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55 +  ~I7d0cbdb63988e88f9f3f69b35029cb2078b97b6cc9008644b2721eda7fb6cfad +1;
assign I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[2]      = I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55 +  ~Iea2bd90043dd35ae24830a90ed10d12869de66637ab0237a1ad459fa916b57af +1;
assign I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[3]      = I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55 +  ~I0f54db0f4bdec3ff62a8f1b5f4974982e3600a906dcfc79789fb9fac058c353c +1;
assign I35669121bfcb264925a80de8432ba33859173e652c8c45d316130a2e034b9bc5[4]      = I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55 +  ~I9a4f77c8ba9a40c1b543070a42451ed37c0f22850a4734cdda393e69c7b54733 +1;
assign Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[0]      = If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75 +  ~Icdea1f407aaefacb918babc28247d540a8a52d513d26d7fbb5e81a41797e7555 +1;
assign Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[1]      = If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75 +  ~I83ec3e2a8ec621acd2afe475255e144f2158e1941ec685a346b75fc471b9cb76 +1;
assign Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[2]      = If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75 +  ~I25600d0eb62c066eda0baba4269851387918088406d117377eb8bcc2e080e426 +1;
assign Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[3]      = If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75 +  ~If45b8fca9a85788040c10a47569139b44384357512af96ee7bd8cd98d88f8f0f +1;
assign Idee00af7413553c8fe7955516c783565ac9a66c62588a1e05723f15cc052636e[4]      = If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75 +  ~I926233df0c5e8461173cedabbf49fead4b0ab577d82f2585af3a1fb6e3130e21 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[0]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I979c6bc2b8486315e3db6888ef068b88396857d05a62470d4f3c33833cfde130 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[1]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~If2b1e365b8ee6d4afa8536f5c2f5c80d31e86ab6729b26795614d75a6a18ef42 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[2]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I50e7a3df23a8147b9a87cb5e38d44bce7613b2a717d1e3a8bda1171f9522997f +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[3]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I3d6bb14416567aa7b8883b3d1778b55c251a22ed42b09bb3cbae6a5210cf11f0 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[4]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I54b0a17c9919d856bb3ed7cbbd8e42fd4ffa33ce8c32d45e4be1e28b71426ee5 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[5]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I4a6a17ada186c2bb60e521443c0a5a0248d03242c4ae01b751fcce4abe853065 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[6]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I33d759e40b55a0d83119f5c19cf87e6e3181c7e3eed94eec60fb52f9c376addd +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[7]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I84920b6036437109dbc48865b69f249d82da5c7288a7eb7744ea7ea567e03657 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[8]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I78f0dcc6533ef218ce6959768639c983d2119dd518e988eb3dcd6f0b4de98c82 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[9]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~If64a23ad02d1da21fe63cb33f95d37c576739eb181b0fe50d7a5101817b4ede9 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[10]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~Id4cd4fdc9fdb1198c2894543e212f665c925298f1c92b4da9c432eca9442963d +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[11]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I2e15c5739b990462c8a17b590fb7d60ac9c7e6648b79e75697139f55221fbcc5 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[12]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~I294ca1e2c287bbe18783f7043149078d4fcc1c59e24792d75655fb29a36e33d4 +1;
assign I5103d7b356a9808a39fb545d2912ed75756cb376686cbe8031d04a1a51b54248[13]      = Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8 +  ~Ideae854591637828f033505e4fc9dee34d82369d02f7680ef6887c597ac1ac82 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[0]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I597d0e1b64b5d47502804c7ba47fd0c17322bfdbd4d332b11f9742713f76855f +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[1]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~Icad68e9babee274d9a5b79cf432d9e2a1938e06f51aeb564af6936972b3f8e54 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[2]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I15b5266ec781a5ae11540d23bf8b1a0b2eb45d94ab6f367a872885ff3207d5a9 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[3]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I5c1a09aa19ef4bb254881dd92543acf840270aa36ad4e0f5f63a6182a4c93a1d +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[4]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I9afcfde9391d485e865b08f9b8ff69cc2ecaace5f5e26e27b7e1775b625722c0 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[5]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~Ibe932d914d189b275138de8d6f3ffb914940d4b2bbecb574fba3c6aed885c44e +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[6]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~Ie2abebb2c2604e435cea102275e0726254ad91df1973aece477e1e5315f82d0b +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[7]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I8befad7180232073f2f7db5a3f546a5a1af79b21cc9cb00a13e266db4eebba48 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[8]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I3a9293b8f323c7e097a099fa6beb33ca299723796aec9396365d43334eb55e35 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[9]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I52698fa0d5291f0dc20fb5f24c33e968ea63f47765bb7d231720330b624b2fae +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[10]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~Id8d0e36ce1faa76feb8cbe0331f2179ddfc066b70e93e990b5d5bce17f505440 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[11]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~Iaef8ec1714d2faf3d3b947db31b7975161077ca31fee04842efc1f7159104d30 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[12]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~Id8da43222903044cc48243a7bcce7864e66d151673396879258ee4af7008a706 +1;
assign Iad2d1fd4a26298ea65c068bce2041d41648a657025ab57462d26ace980c1f091[13]      = I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68 +  ~I8eb86c8d64d83d4ac46667af42b6383e4d165459475ec6be9d547a70ef0248af +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[0]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~Iaf205cfa67ea9b2c39d6705da465f081eb75c326c1d80e63e1331a098ca9a4ac +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[1]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I16ffb13aa3dfd9da5da39d9b2246d5ab46fd0fdb7c02781abf4d8bd754bbbdf3 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[2]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I9a15ed1b2fa413056071c97b4f003717902f38d29805752222c45cbb2cf58109 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[3]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I6a10084ceb62d383dbc5871a208fc087b23de418b2c780813ae950bf4e594c96 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[4]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I63f5ecb10fc3ed9bd8bf79403afed8ab1a70600ceb1e755de0d44af98495ea88 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[5]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I377aa224e1817d2ab5cb02a5a290a723621782607fcd59b319d8cec1b092bc1b +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[6]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~Ib1310cd21337a1faa061ffd12a2670171f582e03471ab315b90de9f8fc30959a +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[7]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~Iabc9fc6e9581216af19559d8e709ea0842cba4f29f3fdfb05bd71d6d9f7594ae +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[8]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~Id165331f616d7e8f347cbe46daff955009fef6f8c0310c64c01dd35990231279 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[9]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~If17c7df712b5dd40132ac60628bd514bc70092122a0cb89ba7d4559439779fc9 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[10]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I9d7506b5ed3de0e32e821ce6ddd1c28aed177910ccacc4d4aa2a8ee57212d162 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[11]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~I734136c95a40c62745d684fc7e8cd1114b883c6209df11cfe01b9174cffc720a +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[12]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~Ibae97ff31fce14dd0506fdfe7407fd6260f7cf8584a01da77312b1aa48594be0 +1;
assign I5bcf3ef731433466e20a7f327403b22f6c125166231fa7b045115a5994b6a129[13]      = I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b +  ~Iea011619fa5b0fb7d22dc4bb4ce3fcc4856dfc7286ff393fb329ac0d7e348207 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[0]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I954e0367a6f3af96a7e033da51e7256543d7eabd37191d4b03f3077567cb629f +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[1]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I1e6d7d9769dc32e1e014951538f1cd1014e9d07b675e6369e88ad5a6fd400787 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[2]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~Iac4172f940fcbc93db2047b26fece588f3fa63ef255ef404beb5e6ea016b2ba3 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[3]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I0e9a7c6c53b89ca2685615c270e8ef3d3f51fad8619953972e1037edfe633834 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[4]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~Ib99b447a19aa10415461faaa8d8026b0073582bd078930f2cdf0f531259d9c50 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[5]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~Icd30277c9d839d833f27f571231dd138497796d3e7818460d836a48b87e34d03 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[6]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I2862bdd9be64c24d98e80e8b662a7c97c70943bab3d49cc8d39443abcd5c2c3c +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[7]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I4f73c51d25db7485bf4a0d63f95f14fc0661431870ce704f70cbb787eb336f09 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[8]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I2647390c3800518f2251794a7ee4aa2d71ca9589534cf73eda0accbd2b3342da +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[9]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~Ie05c1da46b594d3c94aac179f6c98334d0d667cea08108719b44541b7b0a2049 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[10]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I1bfa3da571b0e3d943ec7b9a8c641283e080bcc6502fa8317ced3c0a6eb2c4cf +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[11]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~Idfa7c6c8248be1a2f8a95c6c74a71be3126e039a31f4e16e0b964476c6d47953 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[12]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I5c43417b1bd96dfedeb36f6d3405fc7f6b73c11a55f21ebe6ffd675e991a13c3 +1;
assign I69cd8bc4d72be249c7d35da67425e793b67caf3e00c2d983e9d1ee15d26a440b[13]      = I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e +  ~I71f31c9a9943d9fd422d00aa01888aac32dd8b34236bdd9bdf3e660413a3512a +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[0]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~Icc43ea934f0c07465170977b52d2f402fe155ef77f3ca27119fa665a1d918694 +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[1]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~I78abc91706fec0893eee10a69916f7247b718169155038bdc0bb6f8661ed1c3a +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[2]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~Ia428f915c49f84567006696ba3f5c783035325755b4fefcf74d65aaae1f3d3c9 +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[3]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~If270910122bcee1c18cc592dba9b38c026f792d8d1472400a09edee9d7633e22 +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[4]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~I1517acf28729695d689aced1c7eb358d9acfc4453fedf95a76fc22c972550c63 +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[5]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~I8ca8dfb7a3a8ecb9eac34d1d1ef4768d31b86a757cb7b9ce61ef159816ceea7f +1;
assign I25438316397f42f06fc00bfa8bd5893f0bd54f3296972d59f0a975310549dd64[6]      = I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a +  ~I2cb1ae23e53b89ca0fd3d1df98b32d5b9e478e9eb579b0875981a6b056e8ef4e +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[0]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~I1a2646b8251f83855c3fe8f6172f36500201ce43b9b5ba2cf0f25fd5d540e89c +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[1]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~I1d9a8ff2514f112838c7e4f568303dfcac3f86d94003ec4f1a40a35b79ee8ef6 +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[2]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~I83c8ad082be8fe1a71adac4f41a3bd7019d2df299d19f8e5a293367e49b04fa5 +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[3]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~Idc29625b375c44e890e371217aaa25d5fda337ba8177fcceca881adc72292a3b +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[4]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~I6e88f83ef5bc5f950a4bcb904ffede2603201e72e362aedb8db04412f7bc2bd5 +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[5]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~I7ff25e517e328eda581e7637a2114a7cffe873df520114410c0487e503c01aa6 +1;
assign I7ad97f2a109ae874c27ca94ac967ffafe0acd0867eedca16da50277b0f5cd9c4[6]      = I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0 +  ~I463662fa980f8a5e4be086aa5f37db53b1d6ea8dfe11725b8c407f779a168998 +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[0]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~I8db02445666e4aa12d7e495ba28ca0eae6ef411094d30330e91eb9eb03b38aa7 +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[1]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~I8c971b4c1be575fe328c0a4a9ecc5dc75f08d36f65aa58642976d971a6c316d7 +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[2]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~I09e6d011dacfba2800f9ade6a495076a67e4acc6a944fd649a7c382422e8fa6a +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[3]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~I76599c709cdbb3f3cfe4071b96fb7dcdf8e072fe85ad5c8e7bbabd4f6182303a +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[4]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~I0d9bc57dbbebd429ee5a5e5dabc1cd0bd9f4de95a920346b9e61cee83969ba0f +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[5]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~I91716015389a9d3b1d0cc77327f439e02e54be0d3524b2cdbeed886eea673b10 +1;
assign Ic2e15de888b0562549dca800378d80b2124f50e63779e906eec6193d368f42ed[6]      = I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4 +  ~Ibc3e77c4d6cb28599b7a21c7992802beffb168f54d8dfa650750ffdc6730df29 +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[0]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~I34f861f0a748b0ad1550db8ce40149dc638194b0089cf22e2380a39a49f8c902 +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[1]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~Ibadbb4e272ab1105914763e2790898c8e37a553a1b6726e8818431bf5209b369 +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[2]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~I308f551a8479d066b2a4b473206e8f407082cf83b37a376e6b0e1454f7ea2635 +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[3]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~I58c6fbcd5f77398c3514e6a850bb69d9f57880a387f10132aa63079c0a1f4857 +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[4]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~Ia9d25b6cb880b9a00c9bb27bdb80c08988eee46afccbd578659eb98301fbb8a8 +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[5]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~Ied710d5ba03554d4103468029a9d895c25c10765b6e3d73bbdebc54d7cc7d8db +1;
assign Ic7327ae923786e056a6ded84c0a7f2832a5895df97164cdf0dd3a31d9a616d25[6]      = Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e +  ~Id7dcf87d2a40e82e7f01327d834d5207ae5873a7e5133c3dddead9d0cb9703f9 +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[0]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I982c94b61dff8249f2f3055f60da6e2c2b0b56c403f151168b28a5a211aa6428 +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[1]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I710a57e6c5c8e228325430ba2a5fc32ed9da101d76ccf1d8c9f3397859b39ef3 +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[2]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I2cb87b14b006ce6a36ee5439eb18a4287c5b9ae79748faee259c0435d0dac81c +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[3]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~Ife00518e7b24a5de694b56a32211898b3c23d2dbd2df91a4197216c23fb5aa7b +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[4]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~Ica9ef16b19711ccdfe32e34eed347b590635f1ba7983272eb02f980f80642254 +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[5]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I9331a9d6610ae5cb77aa3d477fce0c0ad7378a884c86c4872a1573f2d8a90d8c +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[6]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I48d9ec419ebe83e2a5a8281e7beac36acc9e554b86b154736dc51ff940f5348d +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[7]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~Iab97067540ba8c9551711cdbff0c6aa3993534d3e8b352bda090a0997c681afa +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[8]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I25c667a6616c9a94f6618166c99298b28d897f9ac8276bb85816e4b42582cdfe +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[9]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I2d2137ac29a7c23160dedc43e9caf010f72f7d08b057e49fcac89984e616fa5a +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[10]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I11775c069ab4acd951a3ca47bfa65c7632a6a8a369bb103d0bb719806dfe0c57 +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[11]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~I6e418efd4b385b2a298c1c53d344e35f593e8380d1c27d7cb62cfe35223121c8 +1;
assign Ib1a2d00f903f9c963d847ef4406c0fa8e029a3594642e401129570720a2b6b41[12]      = I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a +  ~Ifd66abca1532f04fc777617d91cd2d5f4d4fee35c3f075e91639a196780168d8 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[0]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I6dcc482b16866339b78b922f9a7ec0f4a0ef311c353e6a4e107dfcc351abbb23 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[1]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I8c8bc477ddc4000dde6459d7cbc4ba665fd4ecd97242d9f9fe97ca6825bb033b +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[2]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I54da11ab334a3942047eb5953935aedd00ef1a24bb5361fba51504632ae61831 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[3]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~Ide2ca364c5742f786e5408980fbe12322ebcc2920fd99ed322112d3623d9e372 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[4]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I6024b75d70e3da7df4e532e712df56a8bed06352ba0a545ec355f59473929d41 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[5]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~Ia79355adc994f77e150b93a3e38c8bd6f0a5848a212ac64559cf1210ee0d11d7 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[6]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I1b68e82cfc8606d3a9325ff2da047f345e2f34b44eb428bf2a3bdcf42a6e869e +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[7]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~Ia1d4bd5d90332afbfaaac3cd0d8f5fcbc626ec4adbb0b0f16fc80923925f703f +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[8]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I87af49f5f04df14686aef62aa27c16723af3ad05398f00e29788666b27784de5 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[9]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~Ic1211f3a0703e281ce073a20afbabe9b2a698d1cf74f07f099d21fd89ffc8908 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[10]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I2985f4f17b726f40ab6609b57a796727fe46605944c5e25c594caa8dfbea9f58 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[11]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~I6f7aa66db409365eac05a200d0a0f1d2b25e9c37ba4a7db3b58a7298af0fd6e6 +1;
assign Ie5202331e0f88b0d4e0cd13ef5ba2537e9eab88ecb140231b24757adb3aaca88[12]      = I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2 +  ~Ib1e319af12dcd98c09841e8b06e7af86f2569bd7afeb1718bbbd26e30f65c464 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[0]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I30e28a0e32497e3137bb689fdbde46389bc490300e15be88612f28eff07976e6 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[1]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I0b525cae7fe005cf25a07cb0b1486152d726fc74aa55f03480f10af97379953b +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[2]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I3df4fc0f2f099890a34d7b376328da6460d429e2516a5f8fd1aee5a8fee835df +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[3]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~Ib1b15c9e15e963cc4f2e9caa1b6b132e338947224b705b51ebe710d7e0f661d7 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[4]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~Id364040d3b9f1ebf34ae3fdf7465d955b49d7a2f4709219f76229766d6df98a4 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[5]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I7cd9dadb64725f4217f1330c893724a7537a616ef41d9dc49fd2794125e0dc3d +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[6]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~Ibdd77bf8b31352e365f7e6440a57247a8ba62e667b000c1347165bb39f3c7c2b +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[7]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I35e7fd3f09acca79a1003b0a4b7ac62c4a2be93bcf333abbfb13a5eefd7d5eaf +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[8]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I7e269b2e2d9ec70c47570bad75bce0ddf53e85e3cb4ba87f784ca520c5ff1084 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[9]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I0c23517b9814053cd1f89a8b80a64fcff6ae65937dc97199c0b79ba8f7a34ff3 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[10]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I73ecf8ab6430c6343bf7596e671ce01a3e3e7499813ed75c583a7103147b0bb7 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[11]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~Ib7f659da098e577e33fc0f5da1c03f6d3e68b3883ad7888152d2e8684a6177f3 +1;
assign Ifec47f4431982de6f772ddaa617f274fdee595185187d6d5004b6e4f4c015f41[12]      = I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc +  ~I3386ee46348e8c4359b1ea2153bc64afbe76f2b6bc9a312629b8c52762a22873 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[0]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I8c2fe0c8cb55f09e4dcdbaa3960acfd815764161f53c6234273dffe4558644cf +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[1]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~Idc64cee034c1ee132335ae593844b2c46e3f1b1b2cda8699940df311735a32a0 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[2]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I1c7699448a10638886eaa021495d4c7cc378fe1e9b0aafccda001c15484b9419 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[3]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I45b03b0185f9efbc11c707a64fda9203cc82ec2fbaee7ff34610c74d7cc1132b +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[4]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I3097f16921e899a99f2a2b013a3f6d339ac9672fa5e17655ceba4de2d506e151 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[5]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~If0d62663c8a08719b83a27c76fa62525eb14d452d4ff0f33e94c67f58d7c86f9 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[6]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~Ifedfb1db4b16b86149f5eb8b0adf06499331d423c368c0077c738a190a1814f0 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[7]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~Ice24cd0bd76a7d12a0199df195b34f41f7f72f037177656693b3154d102ba729 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[8]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I6148a04ce3733485aeb6c4d20b6117eea37a510aba76ac29e82d44980bec0934 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[9]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~Ia6391e6b0ad4d9fe4136b90a57d121f2b5f16ed4662429f1b85677591fee37a6 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[10]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I5dfc39b913b8e0d00491e3f7f45b6b467a517b5e87baa065097e28e6d695500a +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[11]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~Ie538f6d2c778992e2324a9adbde215acaf7b8dc3a72a9230d4fba2332f3cab67 +1;
assign I92462043de59ef8cd5a4e3f5495d197a534c0f56bea8cbee271a47c20aaa636b[12]      = I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93 +  ~I03929e638a59a35fc0168772ca06f7a502352e03525042ce6d49cf9ecb671093 +1;
assign Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[0]      = I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d +  ~Ieb5e001b45961175497657da7a0340c2a15b6d8de1b72ad68ac3aa7f96a47af0 +1;
assign Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[1]      = I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d +  ~I6d58dbbb9b18e4b347b34e548c70a9bc0d819986fb3a6bcc3ff8a67c1fce9c9f +1;
assign Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[2]      = I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d +  ~I82772b528a8c156f2932a23a720f8446f3062e9605839897b4652bb2936fca1d +1;
assign Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[3]      = I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d +  ~Idb259e613b71ccde839570ff2e7f21a9cb7bf676ffd4aadfb08d6a963bea9640 +1;
assign Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[4]      = I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d +  ~Ie9b1b4412060f1e9acccc1f3ff897bce33f24fea3bfc91266f9e42c1f38aaaad +1;
assign Ic5010e56c6be831bf875c0433df8df328c7d095cbebc4e0f4235a75e4e0d812b[5]      = I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d +  ~I259a9b6041f341013e6ea0706c4e9ef9a77148bc003b3f0cf9593ebd915b30c1 +1;
assign I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[0]      = Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6 +  ~I41a57b30ab1dd9c40a723f99315558a47412465aa3fe967250572e8373aa7180 +1;
assign I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[1]      = Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6 +  ~I42968c25ee2870f891f69991ae3ad8bc1c3acde2f8f4d6c0cacc48f562399c37 +1;
assign I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[2]      = Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6 +  ~I44103a07ffcd818c0d9280b96ba08c32f96edc83a981ec9748ed3d6e9c061d62 +1;
assign I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[3]      = Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6 +  ~I1c886223618a03ba9e18de68462ddcc522338cd26d24b5e126da9da1df1339f4 +1;
assign I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[4]      = Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6 +  ~Iac242fc0dcf37a86cc334319d77aaae46dd223017f2a6489c4e33314eabc9874 +1;
assign I8c1f83764e266b4a8346df1eb751a4b183fd832dd758d40bc26c11f2f21bb2a2[5]      = Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6 +  ~I3225ba7b6d0e0c7a94dfbc8e074ade02b79a66f6aaf97580a451c2d1781a625c +1;
assign Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[0]      = I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab +  ~I25779b63a47c05d4588d4b33fecaff61647609a62fcc90f0f541c6b30ea9342c +1;
assign Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[1]      = I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab +  ~I05bd9a1d7818f4945ddc448149dee571e80dca8b6eba7ab79b17b6f84d3f35f4 +1;
assign Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[2]      = I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab +  ~I17eff5960d8d41f0832a48fe9a3ae0dfeef1bfc44b73eff506fe1d3813398d15 +1;
assign Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[3]      = I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab +  ~I1b02edd5d00090446500b1dbf66a7e674de978c068b81ff0b0fb7abb9ffb1654 +1;
assign Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[4]      = I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab +  ~I2c865426b0f044469b391bbc13f977fdd19dc89c908574ba289388e382d55cbc +1;
assign Id1b1e71a61168a04061cd1ba2653890422f05a5c290b3fbce314a2b7084fec52[5]      = I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab +  ~I2e557a901de23b8442e8002b3560bbf9cb8592b7bfb7a6e2f8aad12843a5a041 +1;
assign I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[0]      = I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727 +  ~I469f4965961eacfe3dd0cb82fce4905e19e6695d71bec95956e8209d2ae39ba1 +1;
assign I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[1]      = I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727 +  ~I6e148041c3612c795f1eb1513a9eba29e0509f02f94971fed189dd9f03d54a4c +1;
assign I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[2]      = I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727 +  ~I2f687e6270528a72aa2f9f9cc0a5a6368f8eef358270329cc40b56abc0e4a35e +1;
assign I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[3]      = I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727 +  ~I661bc8acd80497efe43e3d6fd92bc4107b1ca63eaf162cff5695b35f8d4a7e26 +1;
assign I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[4]      = I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727 +  ~Ic72f2f8a61b8ecf8960d476bcf8fbbfd4389e932377679286e7182cc12c418c8 +1;
assign I4573af005ead82a8524b5e12d9ee1dd4c746a991c3b94073f79d2eb37606c726[5]      = I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727 +  ~I823e337e6437e5ba36ecaf0b1ac6b7a4e74cd2ed7019dd5447355626a8877d89 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[0]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~I1622b11941b00f6d2ecd90320158533a66501a6ddb78defb4464a937f132c232 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[1]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~I9ab473d34fac3327f03768e14c7bb20056aa8a3dd31520d385552eb6d214f890 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[2]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~Iedf1b21de2a0eb04c4a64f9eb34e2b0b3a152d90b1938b61ca45c880eab16ab6 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[3]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~Ibe3e6de02f0c30287dd89b07be5254ff70d9683389574d02f1423e792bd2d534 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[4]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~Iad8ee4f6cd13a9f415cd3519de0179a66cfc993a840b3101cee554b55c0e7e7a +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[5]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~I15123100f4377e14c62cf47fb1fb652badc3bd0e8f0ab4b970a0bece065a6380 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[6]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~Ic0a892c18037ef674c8d94cdfc94cfca47d977ca2da9e678303255b96575f022 +1;
assign I6ef9e0513dcaefc5fa764cdb40985d7ab354088717afb046ed454d14016bed9e[7]      = I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733 +  ~I2c316e8b8cb6b499a7a8fbb513b3067829197cfacee877c35874a2ec686ada4a +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[0]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~Ib3a2af9bef5f5d8d7228a3b49a5e0d4a37a33117e057078a552588a24d46addc +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[1]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~Ia042bc20eb6866de0ab9ca9154f0db63f7d4ad84d553be858a0be88fbb8f7f33 +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[2]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~I5b4ba308b0fc2946fb11b66aa5c24c7b5cb2a21955116b97f3790de65cd2a064 +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[3]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~I005ecc3a38317079c7bc5008817e11017c33671f77364ad9a07d0eff1e0ebf0b +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[4]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~Ib63856036797d30e60f13453da509ace15e3324c25bdfdea5aa495d592e2006a +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[5]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~Ia9bf10fecfe62530ea6be4687ecf78a2ac08c6fc6e38328c2d64a80cb5a3d72b +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[6]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~Ie1447c9e1eb4ed110e6b0353bc5dd2cd14ec645355c3cf897df6f6c5808475ad +1;
assign If8a5fc5985382d4f0969cfe75ebce7d62d235e3f20d33c73ee5e2aea749b5c8e[7]      = If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521 +  ~Ic8f640e7a0c71ddb20a985259b5e48746d28d2898383765c3b78c577f281d27f +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[0]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I3b1d695a626aefa8e5b146c7f7f26a8da119680783da7afb019209ac9fd719aa +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[1]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I1d91c7e9c2f99df4e0523b7e01b6fa6ea3930382238ccfbc07201b7d3edcc969 +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[2]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I7c1e9623dc53c8aa8611b46c0375994510a97c4d49d0b091964cbe4671acf1d6 +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[3]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I1b5d096081c0190c0ce6a674de1afee9ccd766a9cfab0637a0aec33199061bbf +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[4]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~If145a331c8a8abde8c26d2571cc8b38e1eaf2768a4658d350cb602bf8614a521 +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[5]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I86e764dc3320206d9b52013c2d735ff4d27bf6e4a82227486e64b4ceb68dfe8a +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[6]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I4a98524c02346f4b9468666ffaa9d996b9b868a5a8730264d798d7a66b7454bc +1;
assign I27dee96027b352ca164b395f5ac99c551e425f929a355ccd40d7a581e9ab8340[7]      = Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1 +  ~I1187dbcc72f33b4cc3442982af526be4cfca1b5ac65be943d4ec380421632117 +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[0]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~I73ce2860dd9aa9ca2c0d541a6ae1e5069badd35988d922cffb6aef0038cde662 +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[1]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~Iea2dd4d33966d53ae739a16876ac2cf04e1d95374a5af68e59a5703dfef2aa79 +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[2]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~Ic0a386f5301913434a3d6aaea1d56d6acb3484fababb7b8831d09563bd8842cb +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[3]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~Ia8a4fca33add1c3c58b04eafe9d023751882f409c5d2905f77aae3fef8c2b008 +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[4]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~I9cd4ac82c1e6f2dab27efa85314df34a40d8747959eba18330bd424a38debece +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[5]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~I9bcd5f3f4630ce7a24ea4479c9ddfce59ed809dfaad9d767e80295c41b332f4a +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[6]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~Iac7a05e270cb898af4ba32c16445d0dbdffdafdcc5fae209f09367abcff9d6b7 +1;
assign I5ea534084bfc283bd814fa7611ec5d4f3589d86e3c89408e86240a48704d42cc[7]      = I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709 +  ~Iad7f008b5f08f3ba94a0832261fb4add17f0897e3c7d54a250377b813e284331 +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[0]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~Ic072a2fb2ce65ca734c05e747f12ad094cc5aaf9267dd94dba345b5c7b11dcdc +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[1]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~Ic20328b806ccf89387180fe6d88ba762051c6bc2c7f82494129e8c3600108804 +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[2]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~I11855780f53e8711f8eca9370af31f472dffd126c02cfce8154a959f33c68af6 +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[3]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~I39b8420e976cbdf011232d83446a5cb92c2ba58577792c9c61dd71358205e936 +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[4]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~Ibca01267ba9d7e2fe9f8df34a548836390ba12b9b782f16ba40965c00735213a +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[5]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~I105a7d84244a0d9143b9b2a3c64ea6964f7e1f43b7f8f5cb15d579885bbf746f +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[6]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~I1b0f11f3bca53713a53e2ed18fb81f5a25c7151c874be612677f5204bca28093 +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[7]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~I434991f7c09dac3a7bd42fce3073dcbcf8b1c6579822074548ea94fdf1ef4eaa +1;
assign I2b9680d8e8e6258ca19f1204c9e4156671222e8a6c43008566922ec7118b301a[8]      = Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d +  ~I7fec897140c79264b7b7b7f3ae228ed090ff69351985c07d317ff9c0cab1e58c +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[0]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~I82bc7aad8e3adf5b7bd03d9fdac6eea60cb800e4502e3af7bdc9d49139563fd0 +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[1]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~I218ab164221d559f1e8bc2a13f06a7593eb4133134762698eec270be5d4c3906 +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[2]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~I4135dbaf658fb73b41800cd275824d1c9f410ab1b6e555b6c4c8df12f96c5861 +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[3]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~Ief38674752576e92e90fbe2a7abcfc952274123875a95657dd42c910133cccde +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[4]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~I783b89f0c1e5463646e0fceb976f2b27aac523a677eff6e597e434672b0daac1 +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[5]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~Ib0ee967a174d7c841ebe71e144d6303bfc80a6083ff6ad745c76d488dea66d9e +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[6]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~Iea7b69c43ca4b3707d3bfddf19b27616b8686df915734ba86d3685127bfbf39a +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[7]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~Id36acaa2c9161668c95e2cc3e6e852e9243ca7f486ca6c2ae4d124b1a8ddb522 +1;
assign Ia3ee76fa1278f1d1bf056ecba0f557559e8e58789ccef81b4fcfc007066ef447[8]      = I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7 +  ~I325ec6d7bab5ccd6e9c4a7e9b02a3b8c30072df123bf6318bd97f1e8766457c8 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[0]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~I07c37e958136be68b3d658649964c73ca78160582248da1d45eb9ee82c1f679b +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[1]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~Ie17e17c22c7215d0482ba310638db13a96c0943216f9ebaf53c0c29c69971b23 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[2]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~Ie44aa17133d02266160c8fd6f75716f8bc4a3775356cd1ef0f495b13145ba864 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[3]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~Idaf1699bc7916d99a2a5ce0174383c189dca6d7537734b19dc379bd634d0d209 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[4]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~I64aaf806ebf0ead2a4836251dccd62a394b984823592340be94f4ea02e12d766 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[5]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~I152b3a1e710e5a39bac6338591c6597ee2a38fc25555f563beb7a1a967bf4e94 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[6]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~I9ede22dbb56f48c045a1b5a05945124fb97b6ca7e355dd8d9dcfdef6e623b953 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[7]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~I30e30c2bee3bac86dd68fe8364f818ab63e91d65c4fa1ef45fcfd03c9df87cc5 +1;
assign I7d846286fe4821fb2bd7a5ae312d3c2deb4e3dd7d80503748b61f145f4f21ff2[8]      = I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499 +  ~Ic0bef9008769fe36d726cf80506004d66e7c843a046653201c9bc2c816115c28 +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[0]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~I252a77c3eaec2d6accaee6de3ba5d0b354636e2a2aef4992eca0e2a74eb4d25f +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[1]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~I5fa628cdc28fdeb96014a4d2c2d06b092136cf2a14a0420bd5d3861b83687413 +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[2]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~If258ff7e66143201e30b3fd451e1b8e2ec9e46596c2653ec836617c093f28018 +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[3]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~Id160a3b60a3c7a3ad93044461ade9ccf0b7a627efa4b1bba84a2ea0d4fbdb551 +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[4]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~Ia42e25bf722566321268c83de181d196619f062381c7fdb381ab5f6aeba6589b +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[5]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~I4f96b4022f127e7d965786f2cac8ee6afdbee96980608c876c6b699495f80b0f +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[6]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~I6a2505f0de03f3e2d303fd207ee819f5a1777b650930b87a235ab3cca5de6e87 +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[7]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~I8600d4c5861319be0efba19d9b66ad483aa7bf648f2132c1a339157c43920c18 +1;
assign I508435928f736ace1c0fc789654f335ea84aa9b035556fa221a41e83c3c6e4b0[8]      = Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b +  ~Ic551d228c593c4304b4ef79a965ac1d9081774282af09d79cd587ef9abcd6003 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[0]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I01d7d3d20ba0eab63d519ae054b6c22c5be4000c846a6a4883ffbbddee37663e +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[1]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I4177cb2b0a83442a271f59bf4f758851d5146ee00d76a1177c9a34d4208b7c09 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[2]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I5df828301af902c72794032c0e55d8e7548c9b2277b2edc77f53796ff8e04804 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[3]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Id595e96924941a80a6ade8778fcbcef39b07a62fa1d7350fe50182fdae302556 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[4]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Iefbb3d08b0b2fc51d2f6b60b25b8143f3f88a705e770396e2f6d050632ded97e +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[5]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I71c3a88492c33461f93d43680f11eae8ef3e9402a4b931c5d31f959a2f8c147e +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[6]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I7a7bbb1d7d9b77199c0b29fda08f8a63112052ffb0a502a05586ced336e13c62 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[7]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Ie1657c5216d7c6e743a23819c08b7c7f2fc8a56793e1bc67fa5c5f3b37976641 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[8]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Icac36c9706c9e063b771faf556f6699e280687be228aebf6ce71f5ae775a9754 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[9]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I8b3bb7a4701d3ef22c71a9631482e13afc2ff80f40e2f0ae75cb2211af5ce6d9 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[10]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I6a24b9c3ea194d09d619dff007c4c6f53a3cbbbae5c9d3ba718bc3546eaad989 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[11]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Ic7af968d25c444d210ebbc7ae563688f4f8a48f38035ce5bccee100e10555047 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[12]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Icb61d0767612534695d9de0380a1febbda612604f373afa55f0339c7a679e99e +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[13]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I58d2fcb7085fddc9250ca075b010afdc2d019c4091f5d115d9520586224a1ae8 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[14]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~I4e5dfe1c7112e24769a5e6aa86584c09ed659fa5d05af38d18183db31189a3a7 +1;
assign I58a903a5ce0a1a646e4cc2b6261735e16215bbabfc445bd6cd2184b845b79ad5[15]      = I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29 +  ~Iff97998b0778cb649d03228ed3acc81c1b3a97f6bc47041c423120b1311112d0 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[0]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I422fb05bbac12ca5df13eb7c0c3fd96a4e819de9669ccd64d40060b5db3f3421 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[1]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I782d29ca9e53ffe86cec8809d7d413c9c5ebd9edb6a0d76db2d0c321312d224a +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[2]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I0705e6f1954b14f35dd7fa8a64370c2f9e6e39b6e265857e72946815d1f994fe +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[3]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I3f9e2f1be98a5d14a8b79b252e9b5a2b3a09304f27a3526a4a66b365b682787c +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[4]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I134dfd9d579ba8b2d72bf1c47119a086fcfb6b7d591cc2c5558e451f57636d0c +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[5]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I5f4870fc880aac0f84130a26e3cd493954ea49eb3804dd17a91b2ba1cea599f3 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[6]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I918037e81d2f9c05c6a8b94c64724b1d0ec8afafe5666df433fee3e296171f54 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[7]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I136f70cfdde5473f8944efa2b1093ed76f82dd06a341413ee2a56054ebef5fd2 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[8]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~Ic02dae50f30bea04d63949eadbcf892ce936efc5373a6185668a20311dd59f4f +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[9]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I54296c97ecd9a699f171f4d7271c761aeea50255010a0a90d2dabc16a0cbef79 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[10]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I50a310ea41e0637bf28b5f56cf11560bc936e15c73acee063c60668bfa905fed +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[11]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I25d2b0d3ff7f684e508a62271f3d29c729dc46478248627013dd91075f8d2146 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[12]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I7f9f83601cb61fece60f94c3120b43ca0c737ee36b8c67ccc917d3a428d8750a +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[13]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~If4fa37977e1db59d1bd7a30b2b0919c997b6e25e0438e01b62dc273d10497867 +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[14]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I66291192ca8d81c8e3f667651d5201cb41b6872f73283d13c6718159b008d8cf +1;
assign I91628be289f2ea3c66e2de4015f77507a13d90a3aec13c62756d603ce8d8f8c6[15]      = I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171 +  ~I4bfef3f43cb1a77ce8b2bf4b26160a161e7f28308b8d2817e6e2840f09463e37 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[0]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I0aafab9f9205eb4a8c16e213e116d949a5c625f7cb2b0f3d124deb80aad2c6c7 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[1]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I9095fb177f965807ae5a73a45c76b1c0b6300c6800b17259e5836adea5a78ec8 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[2]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I3780e5266741d9a9435818f002588f4c44ae518b77a30ede57a3823e1e1e5867 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[3]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I360ab21cba3dfd419f0ca83f85d9633b918c3d24a00214399b0465d7106466ad +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[4]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I2c061ca6ba4299d676b5c6f1e1cc920bc1104e7ac730d207949b952d1a98300f +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[5]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~Ief44fc6df0864dd0766877e0d673847250f53ab137cd9029916ab7149446f9c2 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[6]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I353e1673347daf260e61fbba813cd14f83c52ce3f6e5168c0fa6308d41e93590 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[7]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~Idf77a6217d51b2439f71afbf5956a52a241f2bf8722f54cb166d83c3b45f6721 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[8]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I8ea9b55580c15fa584fb934e010debd92e2e893630de456e85036d583921011b +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[9]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~Ic36cf3da50983e4168cc0a31ec0a86c171714355c0fab18398b8daf57bee1a45 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[10]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I7469c1791d81d0924eb0faa6303565dc78fe9eb371fa13039ff89b92b7f51a6b +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[11]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I9b8a4dcee9668bb71803c25e0ece0eebbf704eb29cfa7b91c47cf48d61076803 +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[12]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~Icf4d3544466d430d71abf2513cfbc16b575af540d369d405ed831753f304673c +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[13]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I0568efb50e0bb85c39c9ac6d2ab3474ab38799257dac5693085eeb0d74859ade +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[14]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~If072f43c0b06c41c30d9bc40dae674ad9052e5533b1308adb97cff2e03821bab +1;
assign Ia662d2d00de75d083bb4296ecffb2cfa770b0791f68a783382a7585ccc92a3c0[15]      = Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4 +  ~I2f05dd0209278c1e661998552da73728c1521c024a7d26f4652d4f151c6e5f80 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[0]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I17dbb17fb2770beac552dafeb238c5e8e7a948c35c7c543508e652cbcda01dee +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[1]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I68ed84b705e3c00d0fb66182d6eeb93f43999532d713f81fab39a36259e0e7da +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[2]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I9d1a378e4d5703b65f197cb76a1982cc10e0c17654eabcf10d9df091086d8acd +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[3]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~Iba503643311c9dc3366b9bb843dcc1ee2f0243c4cf78004a660fca224b36c5f2 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[4]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I05806fb5d45e4d6f569c12116644b625b7ba071eb052ab97525f06fca03dd88b +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[5]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~Ib2630bec8f9f78489ca6cfe0bf25746b720aa422b9d529d67d6dde2d045d9c3c +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[6]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~Ic57569daaae5eb0e66117615c8c6043b5f76b114b5c34b0df50445f66a22849e +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[7]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I5cbbcfd1cfc35b3e78d01b29831195106ebd9ba5907f44dee6761c2b047c4a60 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[8]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I6dc5ebe003a649f0e4106dc27f25387651d43259f0ddafad10411795ee48b40c +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[9]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I238a5c9cd1dcce0d745817081a4b240f74de3de6f18a3abcc42cafbb19a0ad69 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[10]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I53c29303c76ac3c1c02fc9a74eaff9595153ba06d67c08e07790c58e53b674f1 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[11]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~Ia92993e9a66294adf7a4dbe1ea88a9e8be6367da1c05b8df343b3c7a38bfd8b6 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[12]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I329448311438699d3d590bba6ab4bfc9cead805f96015b77617f42d957bde7d5 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[13]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I717aab2686adb8a0688009c23d92aa4475e240ec0747735e6fee5e196a50c444 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[14]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I13a54b612481fe0fdfe8b52909179bb82298c2bff4f10adc4f41215fa4396311 +1;
assign Iff23dc8747d5acf836c4d52c6a7ff3fa7228207ee6ce2c58be2cec86ed4c2e5a[15]      = I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a +  ~I26a27b64a7aafdbcf4a6d058181fb84e0e16767f4bd7a9c45211c4c1246d3b9e +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[0]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~Ie46448d24890ed6ffa2736abb97331dc3ed219b9324bc0e8453eed6aa2a4806c +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[1]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~I8ab86da421b01a03999daa91e41ae95ff58c6bc38566a3deff72633a5ad1cc18 +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[2]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~I20ddfee724da47731a2062b2732598b429c42f7d22bcfb300dc084de362a2bdb +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[3]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~I8d8dbd62189397b5e9189ead2126a615d5b6cea393901e21cd89c255d6672615 +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[4]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~Ie79db7f22cab9cd57482ce0141d83d5c1ff720a7c3dca2c3664feb4a1e2f4850 +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[5]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~Idcdcb2dd5e2f2aff0d7b362ddb4ae1ee4db08edc2c3df3589a7143bafeec0bcf +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[6]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~I525b9b85b14df7a6533a7e54bdc9bf40a303c890a4a410251c8d556d38b33125 +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[7]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~I65afc937c55081dabf16dbfd02eb03c97204efbdcfbb523609571bb32d537d5e +1;
assign I9ec8029eec0d58725b53d483303572f2a356f90188935f47572b022855052fef[8]      = I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d +  ~I45a11cd2f581121ac03fe112ec78bd07c070673712fe6112a3e4fb4eba298e27 +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[0]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~I9342de9fe82f2273da138f99da619acf144edf1f9c33682fe3b1a09d0121c4d1 +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[1]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~If6cd81d168d83d5f6a7ca18051bbbcea5c7a9e017cfffcf72f31f73275c3a4d4 +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[2]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~Ie2c7966ff2c1e84a7ae016f31b0f8b9ca7aa42eec03467c7e3dda37dc34f070c +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[3]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~I468b28bee4fe1c0d20fe7abd9338bf844ce0a2e322ed6b6de11e2ac621572c48 +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[4]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~I08c55e08731cbdc9703e607b481a65177e7e1e242fdab9bfb014964bb0d1d22c +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[5]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~I6c252caff8f1ab047efc25a950ce3e3ffb47a5b779e37a667c48bc1487528218 +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[6]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~I2ade6ee1b52da04fce9491cad314947a07eb9aaa8b0a430db2f96e2d290384dc +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[7]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~If6e953221a61b86b1fc339b69af853f6ad538b60770f2f7b880d7aa15bd625b3 +1;
assign Ia571bac3304956cb869bede0cb5ae998034063df4940cb228a6ddf5eebeed62b[8]      = I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c +  ~I6c6885b180013a16955ddefa0dc75c25ac85fb76059df9bf8b63af72c8c1fb4d +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[0]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~I907aa3f6584035b934017a601019d35f353b3f99c7573bef60fad167f9d9ffe0 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[1]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~I7ae7cc2f052d37b650c0abeccd841b1b18abb4049c976fbdbab72ea579a5d206 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[2]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~I5c0776e9826af1a98810296a7cb86adde5b1b41c434e6040bc6a5a30172d1bf7 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[3]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~Ia244be7d571a1e41348c37534a23f7cc942b689cbcd5dff8c10043325b80e322 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[4]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~I14730b2825dc07428388347472491ef3abe06da3bcea9b7dc9c919079c22325c +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[5]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~I22670670d7018cb361ca0ffd92516837302d5528c26915b62d22505471ab7384 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[6]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~Ibc34c6979b8f5adc5421ca8603b6dca91161055286758ac10d0c612263077758 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[7]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~Id39c55c4f0df8a0d8ee4f8b47f3de8cebf5343bf75521edfe38a695565eea926 +1;
assign I492ca88a98edf3e13a5a4a9d97befb487bc99e764aae9127c245742b4e9532ee[8]      = I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757 +  ~I06a5cdf2e430e40b5c08ab617356f6b4b0389236041b77e2a57d9d314bfe77f3 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[0]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~I22c3d90c4ad5f41054f9b3dc7ddae143f567182c7fc695c5cd087f126ccdbcf8 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[1]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~I533d6897ed500a803f6f6468e36a2a922495b3effbeb405b47ffb7a5f4d82c89 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[2]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~Ib8d3655f6360b2b189b79353d38c9c9989af811109144d45af0f8b68a3276149 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[3]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~I6b264ac5221269381b155a30c051523f4488ecdc6eb2cf60da80a8b84c49bd96 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[4]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~I5c3a945e8bd4c55e9cb38d19100b13668bd652bc1162d16b30f1562a6595a032 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[5]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~Ief691d56b56a000651b0a4c6cc9f26bc44da82f4a6382550d96ea4101b81ecb9 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[6]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~Icf55933dce8b9f95a57d7d019c9b29f72e08454428013009cf0e4d2c5b6edf0b +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[7]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~I5b0da0701e7399ca2e668c1602f494f41127e4c90e6fa91632da0016e7b395e9 +1;
assign Icc8d5f39acd6cc0b25609a772b388b0d5955fbcfc6823df61ff6dbf6a515c7d8[8]      = Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84 +  ~I6106f96669a63f337b78a6bad5894881230f0ab6467c23ec877cf27a5bc76cb6 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[0]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I566a76fd27d46125a614f5e0c72dff06a0c1d836c7fe4a2c4086129386b34dde +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[1]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~Ic754ed4f2d29b948b422876f371df4f89b86976e25183ce1b9f664e1a9b19f56 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[2]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~Id7310932ca8964fd49adc052220c04855b028e29fb7a48521a36e2dbe1d6d5f4 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[3]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~Ibae8222f76059e8f61dff938a64e23080eb668880ac50ecbb50de852472a22ad +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[4]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I09673e64aaf6f35dbf4aae16ffba969d08a800d32ab25413bfcdbd540d7b01f3 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[5]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I3ae1a42457a669272eeff1bc293c80c67239ef6b725a09eacb82b06ec84edd65 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[6]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I5b4c4554a78c551dd34a93ceb225237a2d2540a0e05311c4595bdaa5a4cb14ea +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[7]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~If27288056468d3ef3052303952f2e4be67796c40d6224383047d71d996f98cf3 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[8]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I12dfae8d4c1a0612c6d65c6f5493247af5e06ca1d8c72dc28f9ca41b0bbc6ea3 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[9]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I295da244d8dab1563a5947230e49171eb905c3758c289526ff6d3e0c3efcebbb +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[10]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I89cf2ce418b6d96c0e2b9c8e82167a47d40ade45a8f08255a1b849a9df9e6d06 +1;
assign I5922f57bca418d81ccfcd880043190142461092836afc7b0386e31af02d05fc8[11]      = I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc +  ~I47ba4d6ad7b1889cb52ff7a1d42176e166270e39a1d2875f3a0cd260a1fc92ab +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[0]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I08240dfbc0f698324c1ffdb8e769016bb8b947fb0b8dbb72839375cdb4cc47e1 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[1]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~Ia9ea47bb0829c979af002fb7aa0e22072671c2876bcdf79365ff2b3691172149 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[2]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I58df4f7ee4282cdb7bb80c9f1d907ff37590b1db22994f3a07b521132ab80087 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[3]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~Iadfdcb3c0764107a2b0deaaf039babe6a08f1018f3718f5539718ed6a5aa962d +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[4]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~Ia2417744c8f15898d5d951e15cdf8c03d932cdac6acd27e32045e0fbfbfe4f30 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[5]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I6d70d8c6d44eb58daff53226cbb59eb647b6dec6bed37021a64e16ac5318d484 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[6]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~Ice3b06f04279add8283c8173340c2bfd4b4801d85610179943f070aef508a893 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[7]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I4fa5ada2d589c7a90e700745aba8e09edcfb0252f532e4c74eb0809c712a36f0 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[8]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I71c6f88cbabd48d41f42f2b16170c8955b79d20b8a8b211e174d1c1473567ad4 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[9]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I1e7e130607ec849c80f9e687f0215ceb767a2650626f20ee44a6fe677fde2299 +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[10]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I4c02563233638e273f05bac3e277c702b38c204fda200dc5ac163662c77a429b +1;
assign Ia1a3594990d0ada8b6dcfc4e896995d6d48665106f3d0ad4208fcfe6ae10297f[11]      = I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54 +  ~I85d8f259f770b22a380d6eb5ace0281c57f0952506152be05f38482c47334988 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[0]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I989259874d3f12b373358db47fed6245f192edac9e7df00531ea7ba75c360d4c +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[1]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I2ef69d9eec4f925b598115d569d2d85a4545871f2ac62635f9b072ba718b595f +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[2]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~If8cefdab8d831c3db83e1ef615ca534f34c58b9903520c7741cafbc84e28d207 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[3]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I00e5abb30adb527f6b32257212dc21f9797e9793ebbcc10feae9e524188539d2 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[4]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I9349cba960e03e6068aa27e997993b0c466e040a1ee9e6053536d3346c84214f +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[5]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I19797110801d39a7970e6d8665215c967071ad9a1bad12c33401b44f595772b7 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[6]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I0d25b3618b50ff21e3f301fe44087368e38fd6b37b6f6fab004824aa9df51f0b +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[7]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~Iba62c53d136b455b7d575b868f2ebd2dadc6003981aa2aae72863a0eb812bd1a +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[8]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~Ia6f2e4979fa9229a647a81a4fa3f8b2af809199049d2554ea15fa9a6ba2f90a9 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[9]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I83d70d4886f48dce0888e203c2c333c76d35f0c73767dd9443ec8fa4790ecb09 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[10]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~I3f92074e96f2c2711248b1d770b4ad718a565a323e6fe4ebb379e6494039af47 +1;
assign Ia333b5543dd73697b7db6b5197d8224d0e9c027dd62dfa50dfce241b73a59fa7[11]      = I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99 +  ~Ia478acf4034b69d392277c3d5c6683346547ff26d418b3a6c36a3f9a56e3cfe0 +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[0]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I06186aec49594899011a9d7bce163a3a43ec094d7c92033df033594ed5eb43ac +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[1]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~Icd8ef17fc44642a3c86a1cb62727eb607e3a4e6d0b021406b9b710ea5c96c06f +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[2]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I2a3d1a32b282fd624497621815c6ff85c904f5f3fb50f18cf345c5a5d7a557ef +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[3]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~Ibb57ab5a5468d08c8b299ee67b535b83995e94d6223d0c6d93dba8580906e319 +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[4]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I6fdc128e94d85f0f7f884ee1ff44fdb6de2ad5b93d83c3e36ae235afcd3d23c0 +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[5]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I2790277776fa84c3edba2332cf538f8ea3a40c1b06cece7463a3b4757b1fe213 +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[6]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I068f00aade8307d2a2e2ddb37d7429a04c2f6786232134a041e62733cadb03ac +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[7]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I07087056bd31363bfb1f76f8fbeb18d1deafd5e4816ca1200d362c0797a77bb4 +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[8]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I01c264f9a89aec9dc11fa16206ffee1c8fb03bcb279e9e9f53fea1e94e9d8b23 +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[9]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~Ie42f89c20abd223240a9f93a89ce650ed2f581e1ceab0587a4fea2ddf9f4f98f +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[10]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~I44ba42cf2460fce5fde6d8a9fba799517336268d29b5817597d819a9eb83df0e +1;
assign I59155a6e4e18fad7a0d3f6031841cdf21028c2f571a6379c035d80a40d265e69[11]      = I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec +  ~Ie4fafd34aeca2efbfd3bfd3bf45f73ceea27b613ed242a43666d85f3680ada44 +1;
assign Ida88a2dbb8109dff5f061f3ecaf9586a219f6355e92312ffd580a09126c72376[0]      = I7689b1f287170d28fc72712f5ff2fd209108b000a63e268b12da08dfed6d60b0 +  ~I65cb4f1288affe61a7cd9981878d8519db25d724cecbb80eb3932ccedafcd5bb +1;
assign I73f2fe34b7ee9a375ae43b6d3cbd515175de303a77f64ad277094e9bb8e45177[0]      = Ic114200c11d550dcee2bd668ffd91dbdd193a00571dda2d6f99b4985ef999f83 +  ~I577e642ba232b9a606abfddc4d84ce4354744e2f953da3b285e417dbfc5aef16 +1;
assign I9f9254e3af43fc1c116a2d33bee39fb18594b7696e59d5aa4c3884363616a5d6[0]      = I2090cbe74e266e4385d5075f2913013cc38b26c5332d982cabead5dbe52d7775 +  ~Ic68515eee7d422be9cf8950e48b81d743d5491851d5a117d1f9b70d1d9b55060 +1;
assign Idbd45e6a4aa2cf66d740fb7d3c41c5d4af78bdfe13d321e6ee7eceb153e03de4[0]      = I7802f219761d40fb4b24650bdbbc6faea69cf01618fbddae575028e96aa7c627 +  ~I0ca47358f982879bb85bd78f6bc19192a5ed8c62214073342b37b040aea331b2 +1;
assign Ie3a6f677abff075b84cd72fb72f4b4ad16dc2a915b2d3e06d8136c5073549499[0]      = I9e11bb32c337ed1d87274c3040deee6d8813fd3f6795de87aeab9f93686ee409 +  ~I1606027ef88387f2150285b55cef89212359f49ab1a49fb71e457a3dba0c438a +1;
assign I6444b0cde8c0fcb1cc0b51c11d3937bd156b26f21a0eca3cabe0c6b0e696f7c0[0]      = I08382faacfb31fa012c97cbde6527792abbdf2c9124d886540d385dbf39e24a7 +  ~Ic09f51154140ef91861243d7b35f05961565b368264d44c8fd5d0f85bd0fa213 +1;
assign I1d41ad001c01e3dc84cd02ab5ba24e8239e273f81dad37de1fdf873305e073c3[0]      = I5c8ffe997fea9d77126fb36c6deb4f9b9c9b38e6aa562b574011ee5915a00857 +  ~Ie28425115106f4b2405fad6fb2994a76e64dfa60e7bc165f46ae67411932a1cf +1;
assign I75cef0e0547fa056ba6e20b68cadef6bea875e9b12fe99c286e8d79a40c9043f[0]      = I6f9b56f1fa7e83cc6acf75b74037938bcd08ba89ac2cb3dbf4df512fc9d521f8 +  ~I64862889bfd7d2a15503bc07af594be59cbaa8758863f78311d6f15ecadcc99f +1;
assign Ie4bd6fa32fac971db980d5dae63887ea1f4b75f375f1953975e4ead5b727d37a[0]      = I3ea241ea179029fe0c486fead3909ff2c05b2d47e4484549d1d521a4f891a9a8 +  ~Ied4424f3e85f3fb92f4e40bc63909f4e77698a18a1d0ee651e54e4de06ee330f +1;
assign I40f5e53051d38a2da1e0c992989c7740e6a7be23273e1412d01e853851b97a0b[0]      = I6f9fd1c4756d8d1250b0ed96355e2739d3bcdaa3603b7e1cb5cb0dd0ad5985e5 +  ~I6c850d46af2f31f4e3d31c3fd2b2d9c7471ccf817b452a4fa2602485f5e7f164 +1;
assign I0e9c027df8259f9e499658f9ee700b50ea04b829312da04e92f13edd2af302ad[0]      = If084c3e6863c87018f76e95d715c83cc83dd85ddf7664f98c6ff35e8a0ea40d9 +  ~I1a1a9f7ee74e17c4a0d7064ca9fae938002b1b685f3cb6309569081b0d971aed +1;
assign If5d8bf4cfab249bae208cb278b5fc90873cebd7a677b1d1e22df49b576863146[0]      = I7fcd9ade547e48c042200e4bae7d4699b326df8a285204b7e23eee2a019cb01d +  ~Ib5929b32be13a8436b74dadded1f26d3742e1424b6025d1eacda112bf4749a15 +1;
assign I03501709a4343537388784e4e39cb9c1b52beb3749d09e2daaf1910dc5b1e2b2[0]      = I9207b21b45d4265cc52ef02ed257ea78cc5a269d98165b2a7714a25b1c477521 +  ~Ibcb7809e1db6cb82ba62be017c5b8685cb6f988f85a0d29ce2459f6ac80498dd +1;
assign I46aa1767826fecc6fede490a807238d69235f3cdf96dc753215e008a12454119[0]      = I4322d4cf469c3caa560e48f6eb1fea264c42dd76b65977c24c676681518691f8 +  ~Idb971d0017094cf8b28e639623f85e6e5fc2c03a1da1e19a1ef87b959fe8e1cf +1;
assign Id749da645d127d8ff383558a6e7ab4a5c2a59f513cb7808fa4dc4e9f6f14f2b9[0]      = I924625bbe810db6c8d5cca4407571d5819d0f7361e2d7f1906bbeb822457aae4 +  ~I89373d12365deb440d5337a2586fcdab81347ca28ff6f261a12e35a235bd23c6 +1;
assign Ib15e62b641f64f20a1d3baff39f2dc6a403616e09955f5d7f47ba4fc093badc9[0]      = I3a01e4ea96fcd387a6bda68d7d07cd6b4e89ca653c798f08ac8402696b42a371 +  ~Ib8f9b76d6cf7a74f0d437f634ce888096a0d6d81d66dc6c60b62a60006b661e9 +1;
assign I603d7bbab10dd31f19047e4a73046c804506ba70d1504351984be41bae1d180e[0]      = I96114d8145aafde7f8f5666ca2f6dcea9ddfe9796f2e3a54556fb1b23fb1a331 +  ~Ie55394a5e3d49de60fbc4f33b3f9813b885da2049376036c935e8cd7c85010d7 +1;
assign Ia7b80ae8cf2697315846253262614611c079c53ada59bf7d982596ff8df770b6[0]      = I006672e4b2c9c693fe5b05655ebb6f31e96ca8e2c92eb488cd28e5a940e49766 +  ~Ia6240db37d8e82731a264e5e3eeabb88e632dc6445647a26b4abdb142ff44c03 +1;
assign I58250efea716c203d1475c4046ca67a47a156f9e4709d26d4b05a29ed1578337[0]      = I408f22a4a77906024a2e6ceb970b39ba9ca76300fb2584bff35e37da452c6613 +  ~I4dfaddc409bf6d3698f255e55590182c2c8c067e0766311322460720dbd0967d +1;
assign I50cccb280c7d65372645e94b4a4d472860f246a8a6d89c02e4feee7dac903e8e[0]      = Ie84e7eb709edc06e55ae27284cb93a0c656ce8559679c49a47c7f03f0d64fce2 +  ~I1dd3e1e1e78d9e24a54fc937e7a25fc0e2514eabd1c1cc662d81ba73aa44680b +1;
assign I01d4a1a1123a68c80a967604072ca420c79d4e205c354221591cdbcaa24c4050[0]      = I84fb24aeaf533382e57c00dd73683ce0e4f5f33a0e7a3b36f2ab00732891682f +  ~I80d4a0cc8b63f2ce0dcb344da5a47c95cc28b5f93d5bc6b77e9b875cdd58db99 +1;
assign I702778e2f8308e720ae6aebd003938631b4a76341308834c90d10eeb3611ce3f[0]      = Ifc8b49d8467101e2eedcab4b6ad6a73e4f657c0e995ccaee5dee276a5ae916b2 +  ~Iec19b0b63d20ea69dbcb23411a298bb6e833ee523fdf082f9343a695891a990f +1;
assign Id2ba36bb60a1673c62e790e5ad15a4fdd49bc397b3cba8e6251a88e63c249091[0]      = I001fd8ecbe068f57df7498db3f519cbb5a65bc5af187f1d34b5eab3df45447d9 +  ~Ib612f39370c6527c5f6eedb0eb5e7676212642673e940402586e823ddcbfb4c6 +1;
assign Ifb22aa4df653a2afecbf1dc570c526ccf003e19a0f5972b9bc5ba9458e316ba6[0]      = I11745815606a2dcec9059a24625e93a31b0f15d9b81c97403905e00d3fd64f43 +  ~Ifa501efa24e47050960fb3c383458a20f54abcbc5ca45bbe2d15a037670cd5cd +1;
assign I43fb6b8f15f49b741ef111f2b4a57e5da84af4d6f3ce9b92e0a2bedb18eef4bf[0]      = I37a341bca6a12362e49dae8435798cd8e7550a16cd506a7f852f4223088bdb4d +  ~I8f088dd043a22011add21694f90df62fe1d2f6670cc72cfee805c9fb49756c77 +1;
assign Ibc1b6326c8e2b05aef237f6ded855eb730c445a3cb6c7d49293ef68b6ec623ea[0]      = I8ab2f0a2c9cf1f1e0401a67f3749b106fac7d45293bb9648325f330e3230517e +  ~Id86d515c6d081de87b9ed3c3521ab079e93ee082d8a0b396d44b3b70cac06b9b +1;
assign I3a8bec62f5e0501c90baaa2f6f7288929d91d107a2197e1c574428638cd020d7[0]      = Ic6ce7ef3f9390c17ef23e718bce985f168504ddff0d66e2babddf08b37dd2819 +  ~I4f94812066080b656de1a2807f5f669b2a81085bfc0470f9868bf5945856b451 +1;
assign Ie8930f54b7806297e3bb1082b70d74d5eaeaf269112a0d5f82caf5c941ff7a2b[0]      = I26c16ba52eb0f661ca599263265d1d0d7e1f155b4afec85407f3ece6fff3c391 +  ~Ia92baf4463c96e210b460ea02d7775353edc6d475d7a315b594b9798cfd17900 +1;
assign I948dbc4fe20518395aaa5356bb504e41a80332a8adbba9ae4c6d8a4ca0704b7b[0]      = I31afedbc324d4ddcd04b3ef766154a6414cc6e31eedb0ff24b40698430e84927 +  ~I9d4c230c86454c5c5f9ec98917ffc8d23fd19105ef93ba860ac2650bcf43ba4d +1;
assign I5140e483e7397c66b8d4835ac2e465f125e62c4feb9835d7a5f5ea7849def4dc[0]      = I807fdac75cca555b8d81d1b4d7e53ae7cfa0e4b83bcb260cadae218faed4f781 +  ~Ia4a28d520896fadbeabee4130dcf862a9542852d87be480b1df2b67817f0ce65 +1;
assign If049a08cd46a811753b3637ee0a96207144b0a5eade57068ba5712c3ba23c8ae[0]      = I0f8a9c8deb02bf990a6ac2ac0569f9d0ad9f167d7c18dc70ba544912aed4bf78 +  ~Ide9498000905141bb106efc7e2184bd460d0e59a2270b10d42f981cf3bd514cb +1;
assign I6b404c4caf16f09360a848f09b33c16a69029ab05067f1bca94eba5e69701d37[0]      = Ib3e6663aab02fdb649843c552944b6e325240f5010acb414c311ae56e78f8459 +  ~Ie9a6b0e499ede3f80403e8f9c795ef4e93108ee8db755e12fb931259f1699712 +1;
assign I1efde896c2d2e97d2b635b34d6ad30d31a8c855ea5975dfadcf5ea136fa3d063[0]      = I41339bac55a76a05186d632423b1fef8173940f0cbddfb64c83282af5cd04cf6 +  ~I362132341c8e8a464a2bc93e7cc5b1d9d7804dd93965614dc340b48fad5c92da +1;
assign I860fff7ccba78c970b447509ccd6de21b521bd8458673134640ce16c6f1ead4e[0]      = I28fb4df9f762474ad496e8689f21d13bcc5bd4fd79190892b78409a06720e2f3 +  ~I4b3c222863418745872c878545e419ee8f9c531f2cba89d28f0787992b0be8ed +1;
assign I9786358e2588e06550a490e47029ce233b6d39273ad261316c5f730a7ee4bf17[0]      = I84ce9c6711b257cb8cf2f09bcc02e0f03490605e543ba12942207df6fabed5ac +  ~Ie39e570f1b5dd9f1ae893af78d81e458d077fcde2aeaba432209269b79785582 +1;
assign Ia01e9ec22c644f28b2be05c8002d4f576e816688e30965ae9f3ef78ca1272b9b[0]      = I8f3d31b6843ca54e80e8f61be651cb7788b43302b001d791357fad349785eb1d +  ~I50ebc7f8f7cf324814b5885b2b18c90bf5007d8030744263d6e66880d836eea0 +1;
assign I0797e7fab1998d109cd09e4aa801cd2dfe57364a83e9c84bef81be8f59ca729e[0]      = I6fb6112b591f6f1495935e422361833f041f7231996d88a3936b5da186e4c48d +  ~I326b57b49d3fcfe654c4cb9ebcd6edc0ad7969e3b531f498e3c31270a5c4aa70 +1;
assign I035ba5b524312fb6136ca853695154f9334f6336e5acf5884beebeff72197c7d[0]      = I959de6064e6c31bf0d18c2d6b4c274ebd5e9fadd996fcb32e695047831716951 +  ~Id3898be2185f86831f58bd16651edee3d1bb21fa07b33a1928740ab496404178 +1;
assign If058a896104351e61394ece6dde5212381937b7d36a4b63f5e99a268d5c7722b[0]      = I0f46fb1c05f0f882ae878e86285077da38a459201c305e13fb4925ba34eaef8e +  ~I2aa77512781cba636ab96a5d09527e1ac34623ea2bb6c6a8d742bbcf6eff499a +1;
assign I29e36792da89f6ea79232a191af837f9da3739332265e00d97d40b09ef384a58[0]      = I99e249a8eaee9127d347ab629dc27a21d5b55d2826c354eaffd9e6fec47b1043 +  ~I225543794992ac9aa68ac3eeea38d41077ab5512b9f3b95fbd65a839294088e9 +1;
assign I5e9d25157a8f35aed3b702ea5120ad81de73bafda0cb5811bae0fd0eaf2d11e1[0]      = I2f779bcb2996facec77594ce5efd7c78acaa443f2b6ab3a5506ae96dcb986b23 +  ~Idd1dac44a6f35d558d400160a087fe7628ef80ad72c3962df2b3a3809b89bcdd +1;
assign I57f4038fbe1f52bf47fe1cdbb52088b800609231fa2007cb1ff941817005a0ce[0]      = Ia765277dd8a5fbb2a65aedce2934fd6c4dc9daa4e0b316604f6f137f19fd5d25 +  ~Ic039114ea8ac4120b09973c79fdc044251fc66bdeb18a498dd6ed7265cdfba2a +1;
assign I592de5159deb6cf98840aff691c78457fefe7ee33d85506cd1dd400679207812[0]      = I1a47d1294e98ebbb0493fe3cf7743d1932eac70fe9d2754367a51d9a49448d12 +  ~I21b3fa431ddc4bc8eacfb17a90fdac2bb32e4d0f4d0118715642c37601a1f883 +1;
assign I262ef0e0ef60c8effdcfb37ad79058672a12fe1aa6b0099d00f1067fb709c255[0]      = I71c11e07942c42d17f5b85b1da8857e91f789966944c1e0948bf5f0285c91079 +  ~I1c6d953c9a0e96d328cc4b515867b2ac21d2947a85e96be19f38e67a8b15001c +1;
assign Ic69f5c16ae27a74a97e7bc6fce24e0c868c1e1e5b6a348410853d40bb11f5d91[0]      = Id810b154e951f2b2d0b8ae826f31effa4f39b3a0396d446ebcceedd7225c5018 +  ~Ib823a58e9d4db87e4d73a81a772a02435af32a11d3c2265fb8a16021cfe4503d +1;
assign I0bba5d4133f73c77eb3812cb20554c368cfe3a6ddc34cc7405b33921fbbd9a2a[0]      = I2a96d9fee197ec3bcdd50abe43ee0d3992f5b03db5cdc958771ed812bf3a0b4e +  ~I3427390162b0952481e5f0728a20075c9cfb814431ecbb1a4014d407ab3b3afd +1;
assign I98234b1225d9d3d636129139d51ebd098c46162cd51cf3530b9c8f8c0f12684c[0]      = I280a4a7c5231cbfe245c071a856f7d1560c4154e9f9a4c5fb6895baa2f4f5871 +  ~I35a9ae1cf23d8697091de65a1d0678632bd6889ae32408d7658e542a756e95ca +1;
assign I31906081d1cabbb8c066a2d5377802f2366fe4f3993b4f749f59d89ed1fe0388[0]      = I01562027a6c7a542ae356bb1d0db0dc55b2094f3470a1894e67a3b7fee9e4361 +  ~I37e54e8ae28cf1a36cb9101d5afd4d523ca9a6ae244efe641c547a4114726bea +1;
assign I735b667ac51f343a3a50cbaf5478e1095cf20f38a650d24285dbb38ba66abbbd[0]      = Ie3eb1aebcdf48fc8f41590f0e9524e989193fd14fae379a200c20d1fd3755db3 +  ~I9544a194d3d75c6c414169ea2536e111c09711ee602eb3462c4022350906a21e +1;
assign I4156cb61e9e7e8947b6750f177dac22866e9f9ad06d7e45bdad1304988857d6f[0]      = Ic585c7a7014e8bff08f28b2d432e9783bea57ff5b456d851503a2c3eee80a768 +  ~I1e4bc72a55efb8462410905dcb2c9a8412e2533ded854d23ca648e0e36802960 +1;
assign I45ae7cee40ada2a73a62a90f141788d37c2a24f503646ce743ae4ac3e43b5bda[0]      = I4f0a460fa116f5a45cd0c435e594ccc7597b449cf5205391a2dc6e977f4bdeb1 +  ~If2cec64e868d25d7fbad45ce4889c6a4cac0084aae00d2aa8963678edbb88875 +1;
assign I5ae0ab8d5ea922fff8bcc268c8f3bea87f11b7d6b824787e972c00a9db0be916[0]      = Ib7f3bef766d8e66cc9002dbcf3538dbe974b70de4d7a8a3d9cc3bfbe815841d5 +  ~I73ad61911b0822e313aab2c484d1699cf2655a42a2bb0a1c9ab36228e41d0f7f +1;
assign Id33bc2a3f235239565a24ba23a93a90e564b2ddcc7559044ccd4f2e6aa6fdb6b[0]      = I027d6136f1b64e5e2f94af338f8fbc0ef9fdf8dd0a2d58aa0eb6879557361681 +  ~I218255d96e659dc8f60cddd40cac94a56d93556ed609b60157d88b298ec95f0c +1;
assign I86a468c8931c4e794856a1c434471a885c62c94dbbc95059bb67ec45a9a722b7[0]      = Ic62f1d181b6452f30ab2146b4e43113b2ca1bf21962f686be46f59084d39fa0e +  ~I11284a18d6115421b4c76054c1a580c41987dec66caa7d5bd9107bbd4ac8bc2c +1;
assign Ibc857d78e207a3c56616aab90400d7f0b57c62f4a5e421ee4b5b7ac7bfa1c31b[0]      = Iecddbb8ccabf830117fa8836a6eafc8dda6fa463d9c907ea25d298249bd066dc +  ~I8516ef195e4ba8f6e29a02ab5ea349a26bb68f6ebb4da847d56c03c942e9c20c +1;
assign I275f7df80a91271f558b5ab22bb6a5b46f01973b93cccebe198f0f3c6e2f2cbe[0]      = I5a2b6e5bff0ffadb36a7f02dbb3cf48ffd37e6e29ef09200db12ccf9fa9d8450 +  ~I2411dfbbf605c7590bc678373dd20b7241356a433756332f9a3445ba8dad57fb +1;
assign I8cc2be0175b91e2589ee8980b860af09aaa4a81cedf23de18f9ae69d0514c369[0]      = I3a9d955359963dadbc16853d82bc2495f84c37d8cabb868a144c5f24d9edb2c9 +  ~I69d896cdb2303b99b73c4d6886f2686381230feca86c62fc064a85e4d11266f4 +1;
assign Ia6661480da7ffc0644e0a42782e89f84535952e5f17f2ecf3f1e4cfc56c532d5[0]      = Idaf457dba6ceb8f056ac34d3bd84bb9e9554c0d55db8928b9b48692c316e6fc5 +  ~If6ca882e537cdf5f458a2e11b7a11f057a3d2a00923825fe236afa0b0e1442c0 +1;
assign If4a3892f82907488395a090155f489b67d9808fab6c5f4cfccde65fc41d3b92f[0]      = Iec8531839aeb35f1c356e474abfc871d1ce889c4aaee1b37b272dd9650fb6981 +  ~Ie35443efbbf821e07284652a4b37347c4cfb959495dafa4fd2f81ffa2edc56db +1;
assign I7b2b5024c5f6f54ab62c8e703f603950e46ebd179fc35e2db34ace053564af4a[0]      = I6a320bd601e721d94d7ac0aeb59e2c81a0a9737d2f7b49d668369336dec2ebfe +  ~Id6d0b1fe00e5324e0ed7c37d41ee3e848f9c7dcfb4a85f5da2b82ed4d8942b21 +1;
assign I709336ccea8dfb4b988c870e3d5c854d77a7acc5ff842b9c2c7490be8e10b3c3[0]      = Icd9be4d5172c268eba385d2cf858caf3450d81a87bb90fde24fccae0d1637d99 +  ~I0a309e8aa7f7e07abd837c99be6d8bb8c29dc1679b449111a02f49442d5cb432 +1;
assign I6ad8cd22867ad477cef7562ef157f85bcd0aeb6ff72ceccd15ecf5c00faf12d6[0]      = I64227cc72d5c6450ebded626fdcdfd149c8e29dcd6839ad76b2b9a932817fdf0 +  ~I416c7ff28cd1d182ba2e08c3882c04d5073a014f7b9b41e56a3850cdc289ffb4 +1;
assign If4a806d211914f82ca329f57517b2d1b1a60a8381bddbd3153e78418258d819e[0]      = Ic754b281b704937ea08e702dcb74b7175f8901b29809052424f867a6685c1d41 +  ~Ie44d1a587dcdbb709546c6c567988fb0a19c276a1df7aced4c09a029196dfd4b +1;
assign I282657b255db6edb8d72272a04f6c69d5b8f32795992f902cbedae3bffba4a4f[0]      = I861b39dacbc8ae1c9cb21a407a53608f0d5adf148148ddb8c3ab1cbce25e2497 +  ~Ic2b8d811fd01f5cd88dd60bb1b89b33163b3cbeae48d04e2316f15500c6a1a40 +1;
assign Ia3f8a8cdad50f5772d19748e82e1e9e0558a1d7973bc2cda424ba8d383c15d62[0]      = I994137ceebfa9f1bfb6f3342c02ef25b1a5e881f6fcf6c2e7f274663b5b4a3ba +  ~I85ff9ab4f9a4a3301bb8fcdc7107202263af0c37f091445efb5fa163a6b47a51 +1;
assign I9ec9a8bbe81467bd2ec058114005f308873b8eb8a8c939f4002003402bc6c486[0]      = I5193db4e129f33dd7cd8691b74f52f030a066b583bbe2d9a4a6e9962f1c43280 +  ~I39ab1bf4bdde9805c5bc7695c4700975d5a6094c40e107b82477192005d9ce21 +1;
assign I2a951c202348bf2bb4da1f79c63a8515c95484c9a16ac1fe9b857fee59361511[0]      = Iecd0fbf7643812e36e8d17ed6782ecf4b181df9d284988b1f416de07cdfe6095 +  ~I602591ae56f1a42c64e50378841e065e79aee138622a0a571effe20cb48645a3 +1;
assign I009b4951ca9d1200c6e7787f401228a9af483223fbb4150aca223cfbb80c8b7c[0]      = I390b2f0e16e0de51443f9cbf8ae301009d17581f5e20ec4956a8e95ede2c0822 +  ~If37e9ed3af8a31c989dc6ad554207cd464c591b630ca1e5cf56b2eca57a18d8c +1;
assign I3af56e36e8422acbbdb52c77327e09618a7b89e21e35787ba522cb8a322ed0bd[0]      = Ia733b3c17807a98828719894627b0a1fb161ffee86fb28c11d92f5b185a6284e +  ~I80099c7b01770cc5f7edb3a3551d8edfe9dccbcd2a12daf8ebbafdfccd141bd4 +1;
assign Iea773cc6750944ca9d0aaaf2dbd818c485ce25a1e333978a68333b521404516d[0]      = I6b87b44befe3363656697619cf3dd967526646ced0f90813c24c960ad4d57d5f +  ~Ie479ccbabaa8a00009152557e4de08bd240fd28f1b131c674dafbcc2505711f7 +1;
assign I5e0342048fa50ff3b98e175c5c8aabadb97e925dfbc34fb7f68376b8eaa3cb1f[0]      = I29ee4a3cefb214cdfe60e6907e63799323eec92930d4a48797c96a7c1f3e3a15 +  ~I6364406b04427fe3a4cecbed48e12a67cb08dc632b2914b0fe52fab0ca541c0d +1;
assign Ie03375db3932197354d4fdbdc800b2b7134470f1622806909963ea424d5fe6af[0]      = I748cf7beef2ac47341c77503d0042b6e1570248031f1d9880d0bf14969378379 +  ~I610dd39f1d44d84764b0acd6b3fb1219fb6b6d6ca92e1b226ca76a389bf6c937 +1;
assign I529cffab52c15bb4db9614fb7a0f353e2867564b31984bd2c5551f5a5d407fbb[0]      = I559b90a32f7cfdeb35bcf30683787c6357460614330553ffd4f5732cc03507ed +  ~Ib9f9384ac4ec4bad29fbb4ce683ffda7dcab311135f02b6336e6209f5742fddd +1;
assign I3bd4e85424803f9f3607ec830b6c73bf1d273e7de387d11359eae7f842fb1551[0]      = Ie6d770decdaac3d75cd6c9eba7edc89898bd152a7c75f43a464a47c9994c9a87 +  ~I60980f76d468775bcc8a7052681fbb6ef4b2243e5e30e5365cda6cf598bd0bde +1;
assign Ie54a4e9ee8bf7646b7e69193c8121ff42b4ab2f266c49916322dec059c92684d[0]      = I6541e01880f3c658b3404a81e96fd03b861ba4a26ec927e9c2c64aa9973dafc2 +  ~I892a754f0322d92126d4731e8066760a24897f93e2afb858ee1393604d2cbb26 +1;
assign Ic07553da54e29d977820e271e50502264b236c156bdf4e3a654cd948a6d4f726[0]      = I184fea1e133f0a5b9b8a88926ebceffbb79cf7816941eaf9a326764d876c924f +  ~Ib0f8816eafd3b950f67cfbdb6a44c59ab7c0918979817a4a998d8305da847e72 +1;
assign I8ba1954b4d7af696e80f659a70d18bea70c37a8f494827a2778c421ca1dd8ac9[0]      = I78d3ad872172f1089358c601e00c98f526455a961f30bfd6a966e8d8bb6bd098 +  ~I04b55f2c45002f1f1f7a6176773a22730dcfea14662f0badb102ddb60b84cf9d +1;
assign I2d1936d0e3bc9f6320f1311cbde5d8e855ebeb68cea0b8c3dcf77f3dd63ceb84[0]      = Ibe18bd1138dcd8295a35b807d811d5b05b07df9efd2326d0cae0cac6589e7bbb +  ~I5edc072d158ac583bd1cdb2449086d4f0b17e36d724f4cfde79820788ce57f31 +1;
assign Ic0b3a57afcb2e31014f5c80d84c8eaf5f7f20d57abd8e863e6ffe0b8146108fd[0]      = I68fb3ebbcbcaf18cb81eeae19529cbcf7fe4175df44bd847d87ba9675ffa862c +  ~Ieb128919ed64e331affb6adba798c267e8c3ec924a7ef58f50b1bc0b29702c23 +1;
assign Ia7f87cbac38cab3ef1ce6466b6b419127464ad3172cb03af43e0f75b9575ff2e[0]      = Id2154e04af88ba8cccdbe100e1c4e4bccbffee35bebd3d43f9229d2915bc1deb +  ~I90cc372cc2f3b23eaaf2cb32da95ee715af64ca2eaee77195d9813647d2a0d08 +1;
assign I27a670adbcc49dd11d8a6647a3220c4ac80946eae616e3da78e7a35f5f522502[0]      = Ic95be152c428a61c5e57fa5a5e776b9341efe9f2d08c73fe0a9d2663b0a974e0 +  ~Idaf65411d995039ea730b6ee4b5ae727325da17dc79c8664270d60f063828453 +1;
assign Ib913fea37f6ef92b53b6ec87dde4020983e78b263662b92008f7241cc029189a[0]      = I6e7d06d6c6a765e6994847af070c889f9c7059754ed634122e0204f750919234 +  ~I977557441002c273f9b9b8748ffa9edceadb342e028ceb581c3bbce9af103a74 +1;
assign I1b653b0e5ffe67c25c7a73b1e2fc591f5e57174285113fe2c43ab123799c556a[0]      = If0343bdeee565245554859329a0188f1267cab02c325fbe93d4df18606760025 +  ~Icc10ac19a64065f5923ecef4f1353f13c7796c23f2555f8ae6566eb538d77677 +1;
assign I068d321d442274e43788076aecb6c24130003e03ced4df86bf13a33d2ca5e1f0[0]      = Ie090cc0a910baacb33f7e858eddac0b221b9a5c567ebde9bba44380b06e8dc29 +  ~I725c369a5013eeb6b581209bc8a921fccfcf1754137191e26757abdb72ced94b +1;
assign I975a1d7b1fe781bb19e80aba369e5146327185746eb5088542eba76fbd88ddbe[0]      = Ia0e41f1ae6bbe04c95f97b4d03e31d86b4399463bbd9fb5bd714b9c2b58bb23f +  ~Iaa02b7ddfffcecb763aa916a2bc4c3aea58027c89b515c40b72214d9dd44ba21 +1;
assign I6668b8618eebf7c40e35e5a06aa3b131a6ea1b668bc36d9731036b61087013c3[0]      = If4a86cc5d7bf6b2552861b330822e6bf86fa60debb5d503d86e081b720f3432e +  ~If8737fa82b71d9b0e7223baabca7405e148621600bdaef02e65cd7bd175b2d88 +1;
assign I1b4f3dc17b05ab02ad55643162e80975cc4802ba8cbc4323fb017859b3617abb[0]      = I0d2ad8151436f1c3336aae018a92e8bd400452c12972fef401e7ab55030d285b +  ~Id85c2b905d61bcdc87d500d6ede3ca02d52bc3eaf278f087f27fe6f277c91262 +1;
assign Ic69eaf55d245ae896d42f0f702ef6cd804be0d02cfad9f883b3dac30786352d9[0]      = Id2881f7fc5d7a68a4583d24b1a8a9e09928ea1e5e3ec22fff19d4d59e12a201e +  ~I5923f41aa444bebfc18d13202747ff84e20a4753bc9cedf697b9ae8ec3418afa +1;
assign I8c815413903d61f8d5f9a8abbb8b5e6cb133bcf0e084f4a46ceb98fc67f67515[0]      = I8733749031c60ed31e2867dedeae4f9ddd4da169ff086c567288ece5da43decd +  ~I4ac498dc826a9dbeaddf2f013ae7116e92dc772ea55987a4661f18e56a4123a8 +1;
assign I6abdbd209c6b52b3d4c69e83d51d89be9b3b8e719e4f4e15f50afdccb21ea02b[0]      = I9180b03e001160fe9a51818e7641c427a35e0b2cbeda9e6bc0e32878bca05815 +  ~Iaadbb1b235a85c555a6f37d003e87a987b7d9b07148207555eb717b7332f67ec +1;
assign I6f2bfa7344a4516d6e0b959405ab2c16aabea8d70a454d4eab330ffb6bf9ce2d[0]      = I2f00eb344711414f5f6efe7eee64b5690b4610385673a7186711075eeb319cf9 +  ~I6afb533ec993de4f9b04007b355a9cadf08488ee6ca02aec2d7916a4c98a7fad +1;
assign Ie7eedf6171b2af8aa5e550f07c6913fc6e02bde23689f5ff9f035b89ea7f4cfb[0]      = Iea8f3fa357088442ab8048febba14f1e6ae367c6b1a854ce0b2c4861c4a2ed27 +  ~I01313177417c899543a67763ede925dea3ee58ef4a31714ad15a7a3746bb5be5 +1;
assign Ia298bc83a87ee16d194185dec24955ca32e85a919f168cbfc79e0724038e43d4[0]      = I0d3923859952e0ab6d926924645383b83904ee287f1783cdaa7f314b171f4171 +  ~Ibd0ba147d1a08acea707b8c60da14ebcc4ad62e67ef26634777b5dae38af6d61 +1;
assign I78dfe767d8265759b3b1488f6788812b210a952cba86301b7afe8acd0b194947[0]      = I45f444d890e00116a19e16e3c50c555419e910e2413c0277f62032d6ff66ca15 +  ~I1e92e18a915678cc96aa493a00627dffecbd341dc8e022615610061e52c1ac3f +1;
assign I12a747458626b92b4c562f72f3e5fb63a575053284698acfde64b482d44a98b7[0]      = Ic67dc4f0898ca883d489eab901e11caae2adbe1c1c502ab57f5366cc26d4d335 +  ~Ia7b91fa4a1ef16f859ee162b91daedc97927244dc19aaedede898049daf85a19 +1;
assign Id27fc6b236852c780351e17ad6e85bf55621c84757b3014ead5a2b9ef31d2ce8[0]      = I89150482cc550af995633308cb14fc4aac6984b8c5bb09ed4018e5692f8866e4 +  ~I9918d91748722a47f8526008bc3fd4c498bc80205211d5c92acbc511fdb667bf +1;
assign Ic117e33adf22ba594c3e3c03966b6bb0c6827c2c980f6ba1ee5f6ba40da372dc[0]      = Id4c7f10c8e46d38df8e36571905e342a0b283e8badd00d3e4081890010c25f34 +  ~I95d109e37a87827de1455b5ec479dda78a0218cb9db245b80710cdb1e8ead67a +1;
assign I223d1009ee5643d0804f1d58bbeee2c3f61d8b120ceadf46556e379e45ccc061[0]      = I3c6ebb6c57609827961bfb1e39059b0805cec40a48787adfc9b2b138a5012c9b +  ~Ia0c7162290e415f24699688e45850c243397b5cccf07daf0398dda04810b0690 +1;
assign I60bf67e044d9694caec17617c4d9ff59b9be7698c17aa034515ab1cc94d6a5ed[0]      = Ic8177ee86d033bd8ab95b63937a4f80b02ebbb66d4c16d84c8822d133e7cdd0d +  ~Ib9dc17b2b9fc7c228eba40cf625a49a27ec16f8c8a91957de14fb6849ea49212 +1;
assign I7da66be74fda28e419201be145b24b82c9b29d1155ed00f78e8907d584e214c1[0]      = I65cdf21d7c52f9a1fd2d4bb265a678e8b543e0dedd9fdc5cf9e12ecf756e66ae +  ~Ied32ced79448b3f92faf0dca1673559e07372ec338e8c51a750be1c6975a298e +1;
assign Idfaa10639faa52207bae09b46b05e70da4e285f83560fc415e3915d0a0e8fa4b[0]      = Ib047d12eab2012f21895617ed9bff57a0678c2c85235301fa1276f99ecc8625f +  ~Iaddb000276bde734c13ec1395f06c1b3bf5606ad5cb138579d711cecf26ac88a +1;
assign Ifc9a7a5a4da00db6f00362e2b2b91e1ca59a65e8e35d66791a13468302dd081f[0]      = I4864402239c958072b187da428e64688ab13cd5a3ba940785ac5086f81c50e92 +  ~I211ada7f9095ced6b3d20f8f7f67b56cd2e73595481ed5d4c08175ca874d16ae +1;
assign If453fce64c627db639d688b2260fa70ef90f802d31cac666fd4cd757cd574682[0]      = I8d03bb3beaf84d3f94a15648cd5536d5f14020daffea4160bbd12426018140e3 +  ~I0d49182fe7486bcf54c8f68904b4b90436de6f3bc42fab67a4e47f61154e22c4 +1;
assign I1eca2d1c9da79ade1c32a3685553f133098e1e40edd1e8d9c299a961627aefbb[0]      = Id3b64ab87f29683b9210364e13398a54c486d0b8b8a7a5ec6f15c29cf752b5cf +  ~If79b91295d25c503f6bf5ca7c6eebd2ebf6807dd9990ce31e844cee0d8f89dac +1;
assign Id3b8c5a0992cfb8a82d0e9857a0a77472fe0435d93e37978bc77770999bc4b4d[0]      = I2f3b819fb1f865426e38d2b39a1a4a8ea0560e0888f19913e2393d416205f3b3 +  ~Iec1d04d20ec09595743b7a35860b5cb2ec862c20da87c6f899284069c60bdd71 +1;
assign Ia5acd518b995f7c0cb3e2f5303601027e6195fb82489331aa60c3fc8dfb21184[0]      = I23e7ddde350dba3f41b08c523c29dae580b57e09b8fd9d35af6ba3bd4b104b6e +  ~I2126b1597a95d7aeb7d20d4e0f4270e1fc5cb0fe6eb5003b05abbb7e5e9a2819 +1;
assign I588a95ce70c7581d9afef4d4a297b619958d34acc8bb75e4d61729b440945a89[0]      = Ifbd6430f8434621a650f4942f3be3669bfaa802cd912188e4139542d2a64a511 +  ~I72a115d9b3659f31366e1d73d6d9a0793e20be233c3ccab2b513fd79786224bb +1;
assign Idaeda6020813227d8f52db3ade5daa8152deb71aad3e8cd03094b66b7af5696c[0]      = I1cb9b876fadc25322c3f466b101084a68e5a283260303beb238d55ca788523c7 +  ~I469b0bcfe9cfc27a8596782bab479f30aedaa132a5cd404feb1fec4b52a17d3a +1;
assign I48f239b0c336ab3fdd25e5b7758a5e6c3c0e698832c1f4518d3d1bc6845acd41[0]      = I9bd2fc6de34fc3d410b3d5e30c2e9e811c7063afaa6888afd119cdc02e39afae +  ~Ib4c52550766a2cbe0de236d6783edfb1a6a7cb4c2bb9333a9379e1b75680dad1 +1;
assign I7226b2d9a70f4f716635a08aacafd4ef7a6f5fd31edaee6654bac5577e6398c4[0]      = I9e9c82e0f8d919f8e2e03046a1654698592da05002140ff69fdd551598618d59 +  ~Iaa72101e8c3e7fa248ac4d4336b3847c4f602b6db009e9cd74cdd25251d5178e +1;
assign I14a8ff2f5afad37ef2f9494e67d6fc7df5e0960766ad9f9c46964287587df5ed[0]      = Ic9fded9a702f4299431ec45bc00c9111907d62279133f1a5f62e5f6527823aaf +  ~Ic1381219782d18c1cb880970c062eb260d9d3be0b597e1465fc604c0c0c32c68 +1;
assign I0b4e726e030569d30af5272062eab7426f9a6c50a8e71353fc19fa3b0d576de6[0]      = Ib95adef89f659c6d98e43f4a9c43340a0acdf273ea6bfea0b8e99f0751c250e2 +  ~Icf0c3c82c9e458a347212415d3029f192c40152e8525a20b5c9bfed88ccdb32e +1;
assign Ib6234dcd7696dadb4fa7903f2da1ddf0a7f469668b59cde104d9fd751ebea2cb[0]      = I2f3612471464f3108bd427b6427c8fe79dce2b8e23dc4bb74cecb7e89a3b64a1 +  ~Ic5a87abf4c6018e9555de321c141d9754a7de91f1743d980e339ff9cebd63b7a +1;
assign I07dcbe17d78ed40700955c3277dc667bccfdb936125e6bf04e0e0ed08eafedea[0]      = Iccedefdcae7039447a6901e1cac8bf962a9f520d3b343c2b00e654c7e11a24f2 +  ~I3a27e4e3322c28e7fe85d7e76b7d5477f4d4f6acb8cdb876b9a54cba98b189b9 +1;
assign Ie14f4f4bb4b43f4c07d648f32e6470bc1626117d46a927a286a64d093110e0f9[0]      = I8252bcef404ae08a2a748c98d672c368fbe4187f26e788e54d93af9077f92a20 +  ~I11edfeb948852dab396975b53b12d09da7a5fbedc2dae9fe7c687768cfef05b4 +1;
assign I099c775595305f8021cc03ef225be27441e325455935c0545cdc553d0fea3d44[0]      = Iaa2493521eb50d228c5b0619dca5c86b89a165f9855552ce98021778cc196f8d +  ~I578437932d2d1156445b41a1238e0fd96ab5702bc3158ea337a9e37d14d6731e +1;
assign I9bfa196a8246cf5ae88343b221c084738279254b84fc66495e4669083ac05ad1[0]      = I69d7f0497be77c5b1457ccdc35789d454bbe83f7d9eb458527d737a2222c7796 +  ~I3c2c5b5cd798851c7fcb0d0e66ddf81a516ef9bdf4aa4ebd4901532bfb2a651b +1;
assign I9fb047739860e32f32c612e35c96205de22487ff301c0fc990f576bf205b98fd[0]      = I2c40224a96616b7749f39d78a0c07514232a019bf2c9ecd7340560f5aa5ce6bd +  ~I8153d6f17d832da24daaba2909a88f1609e523ad3b6eac7ad42521979aae96da +1;
assign Ib5aae92803bb8df9f7ffc9fe70a6f447be999b64f9d698828709487924cdd4db[0]      = Id95e503df18410329be5e7761b6857182c75f7d2b0268d0fc377a415c89cad3f +  ~Ic10ea001dcd0b864b987bc3080e95b338c1e91247bb90e884e161c926183fd2b +1;
assign Id89ea99f9b791029af271f9916f63681c6881dec4351cd30a7fc9e3ff1b81400[0]      = I5cca65d1f11141b49a1136898dac8226cb1ec1654c8b8846471f1e4c36bcf3fc +  ~I61efe7187a1aaa28235dacf68eb1e1dd97e7cb5900862790bb4d5872d7adbd67 +1;
assign I8f70e2b5b2ffcd04b7a84ba28ab51f0a9dafd95e4628df8b36dba0ccf87c666d[0]      = I6abf4748a0be2d4365fd1d9b53a44c3183015e1bdfb9a3f671eb5beed231eda1 +  ~I3c710fbd5e4dce0c97eb9da2d8e526f9d44d87fa75088c0421353614e6ef5da9 +1;
assign I21a71d60d8728a63954973b41b85f8ec46e1fedcb5208ea2397adfa9e58be880[0]      = I56bb103437d88864c0ecd5bea1ab5a0313fef2b904c52adb559e19bef8f716bb +  ~Ie02f677979058dda2291ddb93acd64f4461f6d75f3a33c21dac97129344f7055 +1;
assign Icc2b71964c3f1484faf865db6f25dadf0a84b62f85a86cae24a8c01baa1ce8ec[0]      = I5596d8fa3572e105a1618deba542906f0ba5acef8d7b0a48d0fe2e4eb3cf7481 +  ~I2b78100b50f7334d563daa27cab8078fa374dca0c438157d1ad44ed3fd9e3456 +1;
assign Ief6bd3a84efa60cd8d09e7f71dc4b3b882f2eeef86edace8634b6355a0ce5db2[0]      = Ic00f466513895a54a6974af570c7bd5aba8c0ecab5612798bf512ca88f27081d +  ~Icdfa68bdad11213dbaa576cbf43ca9deeb1f9f24225264eaeeede7d1aba5fd8a +1;
assign I21ed781b8a01923a17f646d965cd22caccb44b555b8f392387269b9a2ec9b647[0]      = I456f1fae558de9875bb1f76cfbb1840945f61ea1bce9c9bbcd0ead15d4b2803e +  ~Idb39db95234cbfdbbc89fdee230784c703e170b9e932643a5e1b811b24ae021a +1;
assign If070967e597fbcb6a0ce8a28166d084e71daea6fec72b92cad9a59d03c2dc531[0]      = I7b2c627cf9d530af8ad8ebc0d3dbc53988ea1819d98b5e36e1517e21cc954782 +  ~I7141b42fce475b5502fd33035bf37addde06271b2259e158ba03a66843b66075 +1;
assign Ie0c16d4ccdd2d7d6d9e45d2eea233e13674b7d5a1f8f41877267074f40f6a2bf[0]      = Ic61cceb25c811577024c75e771c53089a2adb9f80e6a622eb82f9d8e5bbb6c16 +  ~I245e922da0aa5470370db389d5bc9db33327c905528a1740aa015b7ccdfcc29e +1;
assign I731f6a3be9c5a884fe93ef383fd933c14af1cfb64cd73fc4381d91d4faa2757d[0]      = Id8edf0b11a998a6c5737c8877c9b203e44c777ca9ee01cce63f046a6bd375c13 +  ~Ia2ff4d61c4f4fdf29be87b50e206c308cf970cbad2638e86ba8c2be8d025b534 +1;
assign I77f33c069479b582cee609a1e4f6255628bb7f6f667e6536333c8e99dac1e08e[0]      = I2813295228131e78d6af31808dc1d9a6f712ddc60b2629d5329dc6ee2d07c9d9 +  ~Idd383630385363471e1b17ea946a61194a3cb287d833af386876c3b4ee66e406 +1;
assign I9288b2d29db5e8dbeef47da923a8ea2055a38ca1f37d4d8ed5d458408b154924[0]      = I6736fca4e33cbc58b4658d91a401b558b1fbf9b3496e1830a8d7b4237d0ef125 +  ~I3daa8702e9dbd047a05e5ea044d14b670c2ae3849526cc514be6a511c5c45c35 +1;
assign I8e09e68977d9f7456b662b0d7fe4575c48ddf88f897bbda3545f7b1b63d89ccc[0]      = Id66c49fe8c0d931dab1b901945cc3926c6e7e3d220480a28e0099a0656241a03 +  ~Ia695c63ae87e9a6742c6fecea648a214f5b24ea2b652bb5d83f35d9a59b94f72 +1;
assign I53ec51c004b0546b3dd0563e2c294a6c4b95b21301321aaf80c838931473cece[0]      = I1d8a87a805073dbe04ce0f76953a234bceb3e6027b2a187071b492f644843715 +  ~Ifc31b600cbbf26e78cee82cd354c17b872586c1a53ddd132edbd25ce87d8aa9a +1;
assign I3c0c87041c080ddc72a51a1b6a4fe12cbd62dd40515520e3924dd8cb63728a83[0]      = Ieb9ae0dc5ee16583e8d05536052b61089e8004344fa0e3fdbc88c5af5119f293 +  ~I261e70e693cdbc572e40e81c594f3dac624febb03465bfd0fb864d337e753499 +1;
assign Id9bb31b77b580b8375e799bc74c4829818ee16c05c6dad069736736dafa7a8f7[0]      = Iff41f572ab79a4cc8e83538b32d4861e88ebdd0a9ce51555053943225158c5af +  ~Ia6f7ae0adde8136c7a25f4fed69bbcaa376b5f28cbb4990afabb57a87ec03019 +1;
assign I5800b2a82f1442915cabe6307e4eee8c6b4071bf852ca93d4a7420bd0e6b1e24[0]      = I7f8fe2415810e04fccd129edfe956981aea020e4b24dd85d59991f4ef0131380 +  ~Ic40e94217a2d2c13f4b1ad2766ab1ae4e8ded0b5e0a3522dd51ec806c3e9feef +1;
assign I40886d5f08de09dc76db805b27c8ca792ccded54cd12ba2e6b70c30121ad9f79[0]      = I5eafefae338dc0fdd7610a7cc3093d323fbd397263d3c8b7546bf540e77d60de +  ~I78602c68a4a00f530bda7ba1dfa4820b7faeb0edabc636d6a2d8bf97005755d1 +1;
assign I0cd63486c66b03be7f8f629aa2577ef8849fa2408aa41a58514c75db95432892[0]      = Ie5d6a774e706204102b6a2d413e41c538f5e61284a19c7a47c42e356ea77d072 +  ~Id8e684d92e6d0b6e10b5e7f7ff9656e6fc67c99edaa59b49e453844ae33d23f6 +1;
assign I8dc1d4da11f5cf2226f4d8211654acb056d8fa751da8aab85dc14664d72b21a5[0]      = Iab62db2e5fab6a7735067ea4afe23d7904f71c5b92219a1ea7848fa358da3cdd +  ~Ic9d9001a209401fca8a3f28e39c4b89adc8f4e9d225aeffbb5d30893bea1a7b2 +1;
assign Iaa67bf8b75feef8789908b65a38dd8124db04184092d5a584054726339440c63[0]      = Icdf027acf32cc766a4ab1f19373a58cad87f74c1ca1791f66e958de6f18803ab +  ~I97f666707f6afacfc6156ef498941fe5feeb7424834b4a283139aefb5f50a68f +1;
assign I845063b254fc4b71844ce1e01433e1d8ad7e176fc80530a73ecb26c31bcf8bf7[0]      = Ib087093eca2530f923f55a4b4cddc83869730b169ab16bf26f6378b580da58f2 +  ~Ibdaeb96b71f9ccccfe79b1b3bab77122aa32217b58037d80a3183bf888b60c72 +1;
assign I51b1e937ea9e8b9d8f3d8c8c66d7f69b172137911df42ee5fd10dfc5d32bca27[0]      = Ice19f7340dbb41a6b126bdae27e69b813b5d6f73ba4db6ee79715328be678511 +  ~I574e4843ab81be7ad95cb7027fc3284a8780b07fb8a194a9c991997988d7ff8f +1;
assign Id90613f9d2194b97066ad1f5247ec5becce3f39f02d165502d84b92178a02948[0]      = I575538bdc858fc8c843bc6b68625f1ba5fd33a904937071914caccc65f324a49 +  ~Iaa4463f258ed92a2c85fef0790c47e725c555f37c80dbe366d973c9599a5484d +1;
assign I38b86f50ae5aadaad749bf30610fc173dbfebd9d3c9d91147b1b3afe8d7f1004[0]      = Idea12ce0edfa5df65e47f6496f2a457a03907e9d62de2cb3797ec2cc6c5adf07 +  ~I7102386e760e34e2d0fc4563b497acec7222bd171333a2169fac800df94ea27c +1;
assign I12d2f80160672a05ea5c1aa8b8b52b7ad7872b05584cd462f2fd449b06326ea8[0]      = Ib368839377e69cd28a997a22724c32efdc8820a04f9b5f93d9877bf398ec6e61 +  ~Iee34d958bf4feec1e5bde8a866a9919f29edd54f1bc51cc9c8216b71101d640b +1;
assign I08cb7d15d8198cd0c19dee6c97c2732b1f72f7e00294bcfb0887c25cb0951701[0]      = I67be614a904dd4d47457ba0dc7a19b2e9f8e4231797917ef3610aea55d5ba3a8 +  ~I64b0ef6642050de0690c95be2af9606797be36c1656f1306b87ce3e8131c4629 +1;
assign Icf9ebe6aa27457ed3d8ac986d9dc8260bc590e8c778585764d6021c62b1f9d5b[0]      = I7cd598a52037f986959ad3f02b4b2783a613170f53a7e49573c5da74f1cbf614 +  ~I23f31ebee34c7f4f9c46fba41d41df176a7465c074ad8527205a5782edab6524 +1;
assign If4d6db4bdc3cf9677389d183b78d9ce032dbeefbc9c6374296777d351a8d958a[0]      = Ide70b17967ff52e323b4a51db51e71445ad3c5483c745b2cec2cc338e5f42f6f +  ~I628b9674d7d6caaa70c54539241df2e7a4be0441dde1739b442513c6e4ded8a4 +1;
assign I15ae50aec5944edbaef4ec461dfb5ab01f597a46233c643d7139247b8bc2f6c6[0]      = Ib28a3a83a3be0baf561a184b6de18de0c4847ff892c403bb9da441f017dd5efb +  ~Ib066c9d790586949b27c4cf09dc957e7d28161ab00e8dc6920e4e0cc5ac665d9 +1;
assign I6dc76307fe143582b214c945a6c0a35a4545c8bebb622615b3ff784edeb2d0b8[0]      = I2416ae27b898336a36264980b371003c06275245f514135d0adac28d88379cf7 +  ~I57419941b1979cd06c4fa0e6be943f004dd80da502425ee5b6dabd2239139cd7 +1;
assign I831951ac212604dca0a254f80af9c1bc9a941f743abf321cc91063922eabd175[0]      = I2d58b3296656a43e75a58883e59a576c0bf73dcd6bc28a939582be7ce0a0ffbd +  ~Iabb5703a54942b1bdcfe2213d2011c659ec812f751dc75943b2ce511c81ffaf9 +1;
assign I0d347b21cb8cd8b8a0fb2e002b97a2078bbdf1c6e71a0e4b9cb022e2a0db8de3[0]      = I3f548241255df4c4a5a8b71a4352ffad6c3e5278c73de2b1afd1a1f1f1f94684 +  ~I798a6a6074b50fc61bd4e1b4696560abd2e515c86d47f85e9a3077cf6672acc8 +1;
assign I9c8cc6c27c1fe245ae54ee4a9dbe2f5fabe4c675abb8af6a49a61e6076233e73[0]      = Ic3ef9d69272fb936b5ada08c6eb60ccaa6acf7b139689e5cb44e0ab76c0ee24c +  ~I3f4a8ec7c554b1f0b9d3d2963b0e3dec4654bf07c5b836f8fd07c639cd19d588 +1;

// Iddd9818abacfde7afed60c93129175401439367a77e69ea93e0ddb3bb38e0bd9 Ib8d31e852725afb1e26d53bab6095b2bff1749c9275be13ed1c05a56ed31ec09 Id8198efa3604d164853468608c55efa148bc56e3564d5a30232bf98b8ab43aeb Ie6f0821795a2d09a9d5d9fee0deb445f74581e2f81076cf0395d62fcc7ecd5c9 valid Ib8d31e852725afb1e26d53bab6095b2bff1749c9275be13ed1c05a56ed31ec09 I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0
       assign tmp_bit[0]  =   (I2dd4b198298ce92cd830c48cf8f44e52b67c0a479483f6788cb4a8ed50c0ba75[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[1]  =   (Icb6f9b93ef17e227d2f57c3847914a8f7554128704edef38f04a510ac4f1dbe6[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[2]  =   (I56854af4b0a1cd696d29385c369527c4f33590e2fea9ff200cabfcd842fb39ee[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[3]  =   (Ie2cc2eba03b304bc797ee7dfcf2941bf5f6029158b6b59e6a727a0d4e4e30493[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[4]  =   (I5d86a7ee41468950b09236808805ca3b37ca38dda66c5b5776ddee52a1de4fac[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[5]  =   (If87fcf0bd1f2929b70124d0daf500408fc7488246a9461d240e042b81d10837d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[6]  =   (Ifa793dd52c6737ac0b26547f9463250e0e0009888ee0070476d9ea1a22482d5e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[7]  =   (If943c6cac01443ccf5d36654472b34781046267ce8c6c221ab9e21df6b8a804c[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[8]  =   (I3e949e90840b7faef8e7f89335f93ed69ca59bc0af12cdbf721d3cfc121b1bd7[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[9]  =   (Iefaeebda45a5830ea753c54dec1c00aa3b717016ecb29869a02730ca81b6d975[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[10]  =   (I82ce0231bfb8e48ebe9920240d5132d8fdf9cd256e6fad98d7e9e62f5772d948[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[11]  =   (I6d59da4a8a2a206a4fb2d2f8da999ec05b513961e0b64f0d290fba57c20ed13f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[12]  =   (I577882c167b8be35eb165d6d16362c8346db31a2e31b934b19b657f284e4ff85[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[13]  =   (I34a013e0933f2ed7d89ea8107ce411e3b282b83722c2ad8dbe23b3360f6251bd[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[14]  =   (Iad8c1435bc9caa462dd3d1f54247bb08239201f66dc04f81eff08b9828458e03[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[15]  =   (Ic0a514775996e7bee4c7519298a56e3219e21224ade2f3a3edce1ce0f05dfc0e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[16]  =   (I1b06aaf56646d33ee3adbf357aad375ac31dbee7f029d5c77ad8d81fc451b3c5[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[17]  =   (I898e5e5092570b3228dd42055f93129e5886d8fb2f65811fda38a53b218d741c[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[18]  =   (I933931f0c57ee6d824329af9a28541852dd6ff11b8aa3fe294ebcbb69fb57e55[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[19]  =   (If8073b9d62820d9420dd56a39dac17b98e9a12def959a8c03270a246d4ee4a75[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[20]  =   (Ib496ea4161d370d24cc568402af56dc4f77bb41266baa55ae1e007226fdf90e8[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[21]  =   (I89c6e079daf908bec178e0f6c167f9a4a60f081380b0fd9fb257eaac4982db68[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[22]  =   (I7cede7dfb957613c710fbc99f28e336af8a20812fa0516d3ae5412ccfbf48e7b[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[23]  =   (I5df9364f6b60d06e160c1b302cf6c07f1d571e149d4232f2efe541efdc0f597e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[24]  =   (I747a1d06ca9bb024ed3320a8a747ce84e3dc14139ff1d19b60085b099191469a[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[25]  =   (I2e94b59f6fddfe0e4af2ed2ce372850dde71bf7f5d464aaeba98efcba30c4bb0[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[26]  =   (I3b464fc2517fabb36a427e7776db9208762c633c49c6a2c607c7565daa566ac4[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[27]  =   (Ice54d60dcb0feeda686097445a5eb91a409b8071a7bc97c2289b90ec6b06150e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[28]  =   (I2f7567ea0c3e5cc97f5a8945d34879cea24c71173c7781b0c9b8901cd258732a[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[29]  =   (I3383b83ddf6f0f7a7f335c7b40343a4fc650d5af735dd76b069ed558989e35c2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[30]  =   (I1cc04dc513fc8b0a45c170cadc3a0058b0c16585cbc8d1ee94e2dd1f939599fc[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[31]  =   (I1cb1aed9639d4804432a1cc1723e19a3269ac404280f907951c293f59dbdbd93[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[32]  =   (I583b2703c5ded7dfa0602870739c5da95f002d944e1022898f8fe131fa1ab31d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[33]  =   (Ie8987dbe984ff1335571cf1a0c80dae7720dcf37e987c9e673ff672e7b3cf2b6[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[34]  =   (I88f33c361fedaf959a5e317983e9644c94582c2b66cf5fa7eb6ca9aa8fa5e8ab[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[35]  =   (I8c255e15d38c4a416e429af6cd261bf546dae73bd8f84c75c1f51688770a8727[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[36]  =   (I84402d152e33ff801779c4ca70de5f2e6bcf748c4a7994e04741c7ea42ebd733[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[37]  =   (If11993165e036ff50223915c069f0bf77cf1ec481e6a51eae79bcc2c0e459521[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[38]  =   (Ia7e1812156c29d63fb75c1fb27a74da10ecfc4c94e9cd4e636ec467cb24be6b1[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[39]  =   (I5b62ec069d6ed1348a5686d8a8b462cfcc2fe1454e7881656075769a6c7f0709[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[40]  =   (Ie60a0de83e4a5e351e8fcfcdb946cc117833349e91cf7a4f89fefe01370ef06d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[41]  =   (I3634d41f65e6753d4317d8a772ffec9531afdb61739b2dd8666972bce2b943a7[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[42]  =   (I0abe255d6bb02a97c26c66e5ce21fa6f6d06bf07f9fd7d16f56679b84e446499[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[43]  =   (Id69d5d8b2cfea2d697315c57128736c25ec2764367c57ea451395ab274c1e89b[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[44]  =   (I7649acb4de026a4b601e2f292b5e00ea4fb389c7aae99e424ac4a49c718b9c29[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[45]  =   (I6a5d3a3f286c3062d8c166c8e4e8110877844c75203d918f406cadfe1d121171[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[46]  =   (Ide5924e2a77ed02b93bc74042d5224812bc3f362a7d9519515c2b0eca72ec4b4[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[47]  =   (I3fc09dc8b11e79e40ce2b1ab330c4b6b8694359152e5b10c962992900dcc6c1a[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[48]  =   (I5089c05dfb338de662c99a38d2074b15622a4d2a13b038a97d0bf7d25c6deb8d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[49]  =   (I5ceb1be057a4b3ac28a0ce4fef635fd70b715e2931a06d5fb262ec4f2b6c4a5c[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[50]  =   (I06065ed8fa058100ac75c56af9874d53802b8bfe909fde6dacd769f2018cf757[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[51]  =   (Id21a1a1dc6fa4a77e4d74ec429279f61fba5f041bc599e6c3607782c03a51a84[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[52]  =   (I14f72ec3b7f8e044df7f37fd50d5e21badff32b32e34501722bf91ffd296d8dc[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[53]  =   (I37f868b41ad5beb13975a02bf8a4210f44ce26ed5436ec5050440a1fa42f3d54[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[54]  =   (I7dc3abe0e7d4ebaf67b15d5c5c6b5cc5ea38030302bf0bd7d75eb1a940271a99[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[55]  =   (I2dbbcd7d60e52e70a185cbc75f9a97843b59becd6fbb48f5e8bc63b289900bec[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[56]  =   (I7689b1f287170d28fc72712f5ff2fd209108b000a63e268b12da08dfed6d60b0[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[57]  =   (Ic114200c11d550dcee2bd668ffd91dbdd193a00571dda2d6f99b4985ef999f83[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[58]  =   (I2090cbe74e266e4385d5075f2913013cc38b26c5332d982cabead5dbe52d7775[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[59]  =   (I7802f219761d40fb4b24650bdbbc6faea69cf01618fbddae575028e96aa7c627[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[60]  =   (I9e11bb32c337ed1d87274c3040deee6d8813fd3f6795de87aeab9f93686ee409[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[61]  =   (I08382faacfb31fa012c97cbde6527792abbdf2c9124d886540d385dbf39e24a7[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[62]  =   (I5c8ffe997fea9d77126fb36c6deb4f9b9c9b38e6aa562b574011ee5915a00857[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[63]  =   (I6f9b56f1fa7e83cc6acf75b74037938bcd08ba89ac2cb3dbf4df512fc9d521f8[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[64]  =   (I3ea241ea179029fe0c486fead3909ff2c05b2d47e4484549d1d521a4f891a9a8[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[65]  =   (I6f9fd1c4756d8d1250b0ed96355e2739d3bcdaa3603b7e1cb5cb0dd0ad5985e5[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[66]  =   (If084c3e6863c87018f76e95d715c83cc83dd85ddf7664f98c6ff35e8a0ea40d9[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[67]  =   (I7fcd9ade547e48c042200e4bae7d4699b326df8a285204b7e23eee2a019cb01d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[68]  =   (I9207b21b45d4265cc52ef02ed257ea78cc5a269d98165b2a7714a25b1c477521[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[69]  =   (I4322d4cf469c3caa560e48f6eb1fea264c42dd76b65977c24c676681518691f8[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[70]  =   (I924625bbe810db6c8d5cca4407571d5819d0f7361e2d7f1906bbeb822457aae4[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[71]  =   (I3a01e4ea96fcd387a6bda68d7d07cd6b4e89ca653c798f08ac8402696b42a371[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[72]  =   (I96114d8145aafde7f8f5666ca2f6dcea9ddfe9796f2e3a54556fb1b23fb1a331[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[73]  =   (I006672e4b2c9c693fe5b05655ebb6f31e96ca8e2c92eb488cd28e5a940e49766[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[74]  =   (I408f22a4a77906024a2e6ceb970b39ba9ca76300fb2584bff35e37da452c6613[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[75]  =   (Ie84e7eb709edc06e55ae27284cb93a0c656ce8559679c49a47c7f03f0d64fce2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[76]  =   (I84fb24aeaf533382e57c00dd73683ce0e4f5f33a0e7a3b36f2ab00732891682f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[77]  =   (Ifc8b49d8467101e2eedcab4b6ad6a73e4f657c0e995ccaee5dee276a5ae916b2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[78]  =   (I001fd8ecbe068f57df7498db3f519cbb5a65bc5af187f1d34b5eab3df45447d9[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[79]  =   (I11745815606a2dcec9059a24625e93a31b0f15d9b81c97403905e00d3fd64f43[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[80]  =   (I37a341bca6a12362e49dae8435798cd8e7550a16cd506a7f852f4223088bdb4d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[81]  =   (I8ab2f0a2c9cf1f1e0401a67f3749b106fac7d45293bb9648325f330e3230517e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[82]  =   (Ic6ce7ef3f9390c17ef23e718bce985f168504ddff0d66e2babddf08b37dd2819[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[83]  =   (I26c16ba52eb0f661ca599263265d1d0d7e1f155b4afec85407f3ece6fff3c391[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[84]  =   (I31afedbc324d4ddcd04b3ef766154a6414cc6e31eedb0ff24b40698430e84927[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[85]  =   (I807fdac75cca555b8d81d1b4d7e53ae7cfa0e4b83bcb260cadae218faed4f781[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[86]  =   (I0f8a9c8deb02bf990a6ac2ac0569f9d0ad9f167d7c18dc70ba544912aed4bf78[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[87]  =   (Ib3e6663aab02fdb649843c552944b6e325240f5010acb414c311ae56e78f8459[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[88]  =   (I41339bac55a76a05186d632423b1fef8173940f0cbddfb64c83282af5cd04cf6[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[89]  =   (I28fb4df9f762474ad496e8689f21d13bcc5bd4fd79190892b78409a06720e2f3[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[90]  =   (I84ce9c6711b257cb8cf2f09bcc02e0f03490605e543ba12942207df6fabed5ac[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[91]  =   (I8f3d31b6843ca54e80e8f61be651cb7788b43302b001d791357fad349785eb1d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[92]  =   (I6fb6112b591f6f1495935e422361833f041f7231996d88a3936b5da186e4c48d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[93]  =   (I959de6064e6c31bf0d18c2d6b4c274ebd5e9fadd996fcb32e695047831716951[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[94]  =   (I0f46fb1c05f0f882ae878e86285077da38a459201c305e13fb4925ba34eaef8e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[95]  =   (I99e249a8eaee9127d347ab629dc27a21d5b55d2826c354eaffd9e6fec47b1043[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[96]  =   (I2f779bcb2996facec77594ce5efd7c78acaa443f2b6ab3a5506ae96dcb986b23[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[97]  =   (Ia765277dd8a5fbb2a65aedce2934fd6c4dc9daa4e0b316604f6f137f19fd5d25[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[98]  =   (I1a47d1294e98ebbb0493fe3cf7743d1932eac70fe9d2754367a51d9a49448d12[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[99]  =   (I71c11e07942c42d17f5b85b1da8857e91f789966944c1e0948bf5f0285c91079[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[100]  =   (Id810b154e951f2b2d0b8ae826f31effa4f39b3a0396d446ebcceedd7225c5018[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[101]  =   (I2a96d9fee197ec3bcdd50abe43ee0d3992f5b03db5cdc958771ed812bf3a0b4e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[102]  =   (I280a4a7c5231cbfe245c071a856f7d1560c4154e9f9a4c5fb6895baa2f4f5871[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[103]  =   (I01562027a6c7a542ae356bb1d0db0dc55b2094f3470a1894e67a3b7fee9e4361[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[104]  =   (Ie3eb1aebcdf48fc8f41590f0e9524e989193fd14fae379a200c20d1fd3755db3[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[105]  =   (Ic585c7a7014e8bff08f28b2d432e9783bea57ff5b456d851503a2c3eee80a768[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[106]  =   (I4f0a460fa116f5a45cd0c435e594ccc7597b449cf5205391a2dc6e977f4bdeb1[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[107]  =   (Ib7f3bef766d8e66cc9002dbcf3538dbe974b70de4d7a8a3d9cc3bfbe815841d5[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[108]  =   (I027d6136f1b64e5e2f94af338f8fbc0ef9fdf8dd0a2d58aa0eb6879557361681[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[109]  =   (Ic62f1d181b6452f30ab2146b4e43113b2ca1bf21962f686be46f59084d39fa0e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[110]  =   (Iecddbb8ccabf830117fa8836a6eafc8dda6fa463d9c907ea25d298249bd066dc[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[111]  =   (I5a2b6e5bff0ffadb36a7f02dbb3cf48ffd37e6e29ef09200db12ccf9fa9d8450[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[112]  =   (I3a9d955359963dadbc16853d82bc2495f84c37d8cabb868a144c5f24d9edb2c9[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[113]  =   (Idaf457dba6ceb8f056ac34d3bd84bb9e9554c0d55db8928b9b48692c316e6fc5[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[114]  =   (Iec8531839aeb35f1c356e474abfc871d1ce889c4aaee1b37b272dd9650fb6981[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[115]  =   (I6a320bd601e721d94d7ac0aeb59e2c81a0a9737d2f7b49d668369336dec2ebfe[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[116]  =   (Icd9be4d5172c268eba385d2cf858caf3450d81a87bb90fde24fccae0d1637d99[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[117]  =   (I64227cc72d5c6450ebded626fdcdfd149c8e29dcd6839ad76b2b9a932817fdf0[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[118]  =   (Ic754b281b704937ea08e702dcb74b7175f8901b29809052424f867a6685c1d41[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[119]  =   (I861b39dacbc8ae1c9cb21a407a53608f0d5adf148148ddb8c3ab1cbce25e2497[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[120]  =   (I994137ceebfa9f1bfb6f3342c02ef25b1a5e881f6fcf6c2e7f274663b5b4a3ba[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[121]  =   (I5193db4e129f33dd7cd8691b74f52f030a066b583bbe2d9a4a6e9962f1c43280[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[122]  =   (Iecd0fbf7643812e36e8d17ed6782ecf4b181df9d284988b1f416de07cdfe6095[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[123]  =   (I390b2f0e16e0de51443f9cbf8ae301009d17581f5e20ec4956a8e95ede2c0822[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[124]  =   (Ia733b3c17807a98828719894627b0a1fb161ffee86fb28c11d92f5b185a6284e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[125]  =   (I6b87b44befe3363656697619cf3dd967526646ced0f90813c24c960ad4d57d5f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[126]  =   (I29ee4a3cefb214cdfe60e6907e63799323eec92930d4a48797c96a7c1f3e3a15[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[127]  =   (I748cf7beef2ac47341c77503d0042b6e1570248031f1d9880d0bf14969378379[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[128]  =   (I559b90a32f7cfdeb35bcf30683787c6357460614330553ffd4f5732cc03507ed[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[129]  =   (Ie6d770decdaac3d75cd6c9eba7edc89898bd152a7c75f43a464a47c9994c9a87[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[130]  =   (I6541e01880f3c658b3404a81e96fd03b861ba4a26ec927e9c2c64aa9973dafc2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[131]  =   (I184fea1e133f0a5b9b8a88926ebceffbb79cf7816941eaf9a326764d876c924f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[132]  =   (I78d3ad872172f1089358c601e00c98f526455a961f30bfd6a966e8d8bb6bd098[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[133]  =   (Ibe18bd1138dcd8295a35b807d811d5b05b07df9efd2326d0cae0cac6589e7bbb[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[134]  =   (I68fb3ebbcbcaf18cb81eeae19529cbcf7fe4175df44bd847d87ba9675ffa862c[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[135]  =   (Id2154e04af88ba8cccdbe100e1c4e4bccbffee35bebd3d43f9229d2915bc1deb[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[136]  =   (Ic95be152c428a61c5e57fa5a5e776b9341efe9f2d08c73fe0a9d2663b0a974e0[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[137]  =   (I6e7d06d6c6a765e6994847af070c889f9c7059754ed634122e0204f750919234[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[138]  =   (If0343bdeee565245554859329a0188f1267cab02c325fbe93d4df18606760025[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[139]  =   (Ie090cc0a910baacb33f7e858eddac0b221b9a5c567ebde9bba44380b06e8dc29[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[140]  =   (Ia0e41f1ae6bbe04c95f97b4d03e31d86b4399463bbd9fb5bd714b9c2b58bb23f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[141]  =   (If4a86cc5d7bf6b2552861b330822e6bf86fa60debb5d503d86e081b720f3432e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[142]  =   (I0d2ad8151436f1c3336aae018a92e8bd400452c12972fef401e7ab55030d285b[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[143]  =   (Id2881f7fc5d7a68a4583d24b1a8a9e09928ea1e5e3ec22fff19d4d59e12a201e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[144]  =   (I8733749031c60ed31e2867dedeae4f9ddd4da169ff086c567288ece5da43decd[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[145]  =   (I9180b03e001160fe9a51818e7641c427a35e0b2cbeda9e6bc0e32878bca05815[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[146]  =   (I2f00eb344711414f5f6efe7eee64b5690b4610385673a7186711075eeb319cf9[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[147]  =   (Iea8f3fa357088442ab8048febba14f1e6ae367c6b1a854ce0b2c4861c4a2ed27[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[148]  =   (I0d3923859952e0ab6d926924645383b83904ee287f1783cdaa7f314b171f4171[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[149]  =   (I45f444d890e00116a19e16e3c50c555419e910e2413c0277f62032d6ff66ca15[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[150]  =   (Ic67dc4f0898ca883d489eab901e11caae2adbe1c1c502ab57f5366cc26d4d335[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[151]  =   (I89150482cc550af995633308cb14fc4aac6984b8c5bb09ed4018e5692f8866e4[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[152]  =   (Id4c7f10c8e46d38df8e36571905e342a0b283e8badd00d3e4081890010c25f34[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[153]  =   (I3c6ebb6c57609827961bfb1e39059b0805cec40a48787adfc9b2b138a5012c9b[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[154]  =   (Ic8177ee86d033bd8ab95b63937a4f80b02ebbb66d4c16d84c8822d133e7cdd0d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[155]  =   (I65cdf21d7c52f9a1fd2d4bb265a678e8b543e0dedd9fdc5cf9e12ecf756e66ae[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[156]  =   (Ib047d12eab2012f21895617ed9bff57a0678c2c85235301fa1276f99ecc8625f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[157]  =   (I4864402239c958072b187da428e64688ab13cd5a3ba940785ac5086f81c50e92[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[158]  =   (I8d03bb3beaf84d3f94a15648cd5536d5f14020daffea4160bbd12426018140e3[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[159]  =   (Id3b64ab87f29683b9210364e13398a54c486d0b8b8a7a5ec6f15c29cf752b5cf[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[160]  =   (I2f3b819fb1f865426e38d2b39a1a4a8ea0560e0888f19913e2393d416205f3b3[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[161]  =   (I23e7ddde350dba3f41b08c523c29dae580b57e09b8fd9d35af6ba3bd4b104b6e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[162]  =   (Ifbd6430f8434621a650f4942f3be3669bfaa802cd912188e4139542d2a64a511[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[163]  =   (I1cb9b876fadc25322c3f466b101084a68e5a283260303beb238d55ca788523c7[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[164]  =   (I9bd2fc6de34fc3d410b3d5e30c2e9e811c7063afaa6888afd119cdc02e39afae[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[165]  =   (I9e9c82e0f8d919f8e2e03046a1654698592da05002140ff69fdd551598618d59[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[166]  =   (Ic9fded9a702f4299431ec45bc00c9111907d62279133f1a5f62e5f6527823aaf[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[167]  =   (Ib95adef89f659c6d98e43f4a9c43340a0acdf273ea6bfea0b8e99f0751c250e2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[168]  =   (I2f3612471464f3108bd427b6427c8fe79dce2b8e23dc4bb74cecb7e89a3b64a1[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[169]  =   (Iccedefdcae7039447a6901e1cac8bf962a9f520d3b343c2b00e654c7e11a24f2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[170]  =   (I8252bcef404ae08a2a748c98d672c368fbe4187f26e788e54d93af9077f92a20[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[171]  =   (Iaa2493521eb50d228c5b0619dca5c86b89a165f9855552ce98021778cc196f8d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[172]  =   (I69d7f0497be77c5b1457ccdc35789d454bbe83f7d9eb458527d737a2222c7796[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[173]  =   (I2c40224a96616b7749f39d78a0c07514232a019bf2c9ecd7340560f5aa5ce6bd[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[174]  =   (Id95e503df18410329be5e7761b6857182c75f7d2b0268d0fc377a415c89cad3f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[175]  =   (I5cca65d1f11141b49a1136898dac8226cb1ec1654c8b8846471f1e4c36bcf3fc[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[176]  =   (I6abf4748a0be2d4365fd1d9b53a44c3183015e1bdfb9a3f671eb5beed231eda1[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[177]  =   (I56bb103437d88864c0ecd5bea1ab5a0313fef2b904c52adb559e19bef8f716bb[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[178]  =   (I5596d8fa3572e105a1618deba542906f0ba5acef8d7b0a48d0fe2e4eb3cf7481[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[179]  =   (Ic00f466513895a54a6974af570c7bd5aba8c0ecab5612798bf512ca88f27081d[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[180]  =   (I456f1fae558de9875bb1f76cfbb1840945f61ea1bce9c9bbcd0ead15d4b2803e[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[181]  =   (I7b2c627cf9d530af8ad8ebc0d3dbc53988ea1819d98b5e36e1517e21cc954782[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[182]  =   (Ic61cceb25c811577024c75e771c53089a2adb9f80e6a622eb82f9d8e5bbb6c16[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[183]  =   (Id8edf0b11a998a6c5737c8877c9b203e44c777ca9ee01cce63f046a6bd375c13[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[184]  =   (I2813295228131e78d6af31808dc1d9a6f712ddc60b2629d5329dc6ee2d07c9d9[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[185]  =   (I6736fca4e33cbc58b4658d91a401b558b1fbf9b3496e1830a8d7b4237d0ef125[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[186]  =   (Id66c49fe8c0d931dab1b901945cc3926c6e7e3d220480a28e0099a0656241a03[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[187]  =   (I1d8a87a805073dbe04ce0f76953a234bceb3e6027b2a187071b492f644843715[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[188]  =   (Ieb9ae0dc5ee16583e8d05536052b61089e8004344fa0e3fdbc88c5af5119f293[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[189]  =   (Iff41f572ab79a4cc8e83538b32d4861e88ebdd0a9ce51555053943225158c5af[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[190]  =   (I7f8fe2415810e04fccd129edfe956981aea020e4b24dd85d59991f4ef0131380[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[191]  =   (I5eafefae338dc0fdd7610a7cc3093d323fbd397263d3c8b7546bf540e77d60de[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[192]  =   (Ie5d6a774e706204102b6a2d413e41c538f5e61284a19c7a47c42e356ea77d072[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[193]  =   (Iab62db2e5fab6a7735067ea4afe23d7904f71c5b92219a1ea7848fa358da3cdd[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[194]  =   (Icdf027acf32cc766a4ab1f19373a58cad87f74c1ca1791f66e958de6f18803ab[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[195]  =   (Ib087093eca2530f923f55a4b4cddc83869730b169ab16bf26f6378b580da58f2[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[196]  =   (Ice19f7340dbb41a6b126bdae27e69b813b5d6f73ba4db6ee79715328be678511[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[197]  =   (I575538bdc858fc8c843bc6b68625f1ba5fd33a904937071914caccc65f324a49[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[198]  =   (Idea12ce0edfa5df65e47f6496f2a457a03907e9d62de2cb3797ec2cc6c5adf07[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[199]  =   (Ib368839377e69cd28a997a22724c32efdc8820a04f9b5f93d9877bf398ec6e61[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[200]  =   (I67be614a904dd4d47457ba0dc7a19b2e9f8e4231797917ef3610aea55d5ba3a8[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[201]  =   (I7cd598a52037f986959ad3f02b4b2783a613170f53a7e49573c5da74f1cbf614[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[202]  =   (Ide70b17967ff52e323b4a51db51e71445ad3c5483c745b2cec2cc338e5f42f6f[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[203]  =   (Ib28a3a83a3be0baf561a184b6de18de0c4847ff892c403bb9da441f017dd5efb[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[204]  =   (I2416ae27b898336a36264980b371003c06275245f514135d0adac28d88379cf7[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[205]  =   (I2d58b3296656a43e75a58883e59a576c0bf73dcd6bc28a939582be7ce0a0ffbd[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[206]  =   (I3f548241255df4c4a5a8b71a4352ffad6c3e5278c73de2b1afd1a1f1f1f94684[MAX_SUM_WDTH_LONG-1]);
       assign tmp_bit[207]  =   (Ic3ef9d69272fb936b5ada08c6eb60ccaa6acf7b139689e5cb44e0ab76c0ee24c[MAX_SUM_WDTH_LONG-1]);







always_comb begin
            I7bd679f7d7da9dc0742c725247978f1c14611083c7de896c4c2de108c6766fb9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[0]);
            I11abd59187e2db0058526cb1ea58af9061d439139fa151aaa74184499fcfd24d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[1]);
            I950415762b14dbc0817ccfb0d09d95d700be57ecc9f8011c6163f84336da6e43 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[2]);
            I9841a5dd86a1b359b25fb293e74cfbd88b34e11f22bb61170ecc921048620dc9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[3]);
            I4c8a0d23fea7158b5e99eea187df1d25395edf7df1db8482b41dab7a8bc25030 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[4]);
            Ia6f33a5c8baa6ea053642148b8e414d0b9d17a66f4e71f6e44e1f6c6e3e535ba = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[5]);
            Id7d51984757deb5794eccbf50647e7535041a18dc506aa16b4ba0ad36bc66b0c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[6]);
            Ib8b4f3fbd26b51974ecee1565c3d0c8fa7abd94e467a7369a62ceafa7ea5ddaf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[7]);
            If787a878ae1cab622e44a13190d301d15d0c7ed9271dc50e997c926071f1cd02 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[8]);
            Ifb337611e63cb9cee9828aa75fcb6d978249e65bcc8770d51fb4dd1644c96a86 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[9]);
            Ic3ea8409cfacf50e41b97c65b0440348d06b8f196001ba1fda6348071b47dd23 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[10]);
            Ia49277306313784711d5d8ff63e6a0a77d3fbae050dc1089c734c826be497dcc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[11]);
            I13f5f01dccbdf3df23c5bf603a9657e161c1e2368cb5cb48b212231d2fba7794 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[12]);
            I7c6ea337917ea8eb0696c514db7ffb66719763162bdd0b7e0ac764c1ae63d24b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[13]);
            I8fe688adfc161cafc0777f3c3ac9ae27372603ec55cb3865f90f38f9dbb59439 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[14]);
            If7c696b260799e0ccd86bb377086dd1be59c9d94754dc52605d659391439d3d5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[15]);
            I16ef3abe43350c9096f6c7e597c48fc86ed26a073055b7bcd696c34676529372 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[16]);
            I2f4a0e474435a97fa5d2d056d9de566288c0624cb094d71685934475b58572f1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[17]);
            I554ab27e696a028f48da8ad39e2db6668b57ff692603a9562cd7e8780bfa491d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[18]);
            I78d7fbedde9ab5751194c52134dec1b83ea8d48c4ad77c0b3eb952143612ab71 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[19]);
            I9b494d3414d329e4419da30566795e7b36627870c521c463cefbeb7b48196d3c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[20]);
            I8060bc4cf825f705f2218152b6a7a8600692076ba01123cae35feec231f128dc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e70c702edaeb77dc800fa14726f64f20e292558922ea4ee74f54774dd5dd040[21]);
            I435bc44b4b8aac5fe9ba3c30a74d51a42250154c16d5750e075057d1743ffd69 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[0]);
            Ifc131936849b96a3bcc7bed4c38ebe94d51c56feb4e96d25dfbbcc3670568a16 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[1]);
            I6d0d8fc19811812bc80267dd50fc4742e9efceded7a9428707fac605fac90368 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[2]);
            I15e7d6b702e93b31ac4e46f9ba4cf63da33641629eb9cd414d1e2c8cf54b750f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[3]);
            I26e6175466ec922073d5092cb4168f87cd1289008e4b99400c5b6c2fec3eaf5b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[4]);
            I97449b979933d41c6555a04ba5ba6cae73e44b040387a504f6f7e2ecb763ad08 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[5]);
            I272bc7cf289752b36b9811d4ec63f5c17cb40399f39607b00ba51817fad59e1b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[6]);
            Iff259e6b8d77d06a8354c4d1662328284ede633f1ca4ec4731dcdae94e869f66 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[7]);
            If4cdb00eb64cb9e80d78f3dedd797796f44f471b76f5ea3ddbc6f8521257e4c9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[8]);
            Iac435cdd22e5425837ad24bd6141cb357c302af7ee7637e1cc2ac25474cf7506 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[9]);
            Ic9e13fe7c29048953ae3698eb5d214d6b71367a78bf1042dd6b58064a6cc596d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[10]);
            Icf9f5e717c65afd1b3bbc3d6c1bd960155773ec7790543f56c86637a891decd9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[11]);
            Ife767fdd58724398b336a58803ca328013f3a8228ede0cf108dcae054001de56 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[12]);
            Ic55bde9a87033c380a5cfe5736d205c15099a2f2cf440f88472d7f6e65d360e1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[13]);
            I3af3a7e6138910d118e49b29a6de8bb8e6fbd1cfe13549eb0feea6cd07e6865c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[14]);
            I55e293b2d9539b16ee0f135097b8ec02fc9af54fc96ec3a3058af417b0d04e48 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[15]);
            I3088ff7517eebe83fe5804308d22b8c6190077f576f2e680848092e21116b94a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[16]);
            I8de3f6aec12696eef7d069510ff25e6e620fc4fdde5f92923a707116da636284 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[17]);
            I6996b52f42eb9075a634fcdb07fafaf45c5aa99193446869751c4859e7c1f963 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[18]);
            I3fe543ea18333fd169c6d6e692a5b42232e8abd2b14072a4daba9bacbe921d2f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[19]);
            I29d04420073229582b38d6b3f7d9d638351e92073269d5528b09b080e5fd5670 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[20]);
            I8090d844610f0d62cc25a9c72c2d76d9d6783a067de9c9ea9d5a1f5c48744c70 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie46890afddc5b950a96591b69699d8e74cca1a96d1dc4e1539c4e7210caddc5d[21]);
            Id60b432b19836d2e0919dc2e0201d162d7446434080aff7165fb949aba097f7b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[0]);
            I96248ed668211f13555b4a086e7534b958b901242794b9978d673726d56286e0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[1]);
            I78023336da442165a8be56b4ebf7b41f4bb48bbc2b05c308dcd344c8f36c476a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[2]);
            I05a7291b0f3122dd9941bdd5ce72362b3b0b1803abb126606c82744979184be8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[3]);
            Ia2952eb350b07a9cd76752e1a5f76814ed095eb0ee2a284f221b1c74e38d822e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[4]);
            I9f0d592f1a57b1d3e2c206ffe5a79185253205dfe7b20be53091145aa16f9719 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[5]);
            I62d2fe36d10e598efb7f38f4f57e4511d08c366d7df7f51bfbc63eaaf216035c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[6]);
            Iec33764f14e5b0a736fa76a2313325240a520c065b59c6cdd0f2fc5dc36a975b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[7]);
            I9e89eff507c5a2386876f56afb505a22f00d8c0f8a32635a00501ef8d56ecc6d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[8]);
            I0d6546f557347e1d72c176a40dcb077c9c4c78ed89975154f5bbb3875eb1131d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[9]);
            Idc5ae39b0c3c764ed6d9b7859b7627b97e24c2b4df7d97229a88cfc0c22ccd87 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[10]);
            Ibf4bbd894f269bd6e6eaf9511141b91ac61b5dd3e77b4ffd07aa88474f251ddc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[11]);
            I26ad8ce808bb26201de4f63afd861583af9abc55c7623bf15bd1808c0b0c2be4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[12]);
            Icbbddd7f07e1deff7aacc0e96a33556b62ba127dce877dea351b421ac8d00313 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[13]);
            Ib87cc4d1070a195aa8118b92d29d7c836685de2e44ba1b21388677c8e8a5fb25 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[14]);
            I8dc734304648fe3fba1dc7108e8697cb88b61a2ffa704491b2b9df8cc8354825 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[15]);
            I830406b0cd2e64515811ab932e9ce01d413f0a68ab7939a2fa14e4eee7d04a5b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[16]);
            I113d1ff61779dda7e1209787ba652b8b332fc5811cdc0aae65a304aa89d56766 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[17]);
            If50a43f14a383995b16d784cc119d01749fd30928019bea1b7aba0039c4c350c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[18]);
            I7dd3baf838ce22ecec10d3c1a3d0dd16582497f9e447038aa46bfd49571fcb4b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[19]);
            Ia55512c30a26e336794d389f3700b9153cea83619467b731571ba72a3a9374bf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[20]);
            I799968e729d7842ce09a838203458d89b96fe9d2d7a5de0cbac32eefbf834898 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42015bfc527d6282348e721bd286f2ef74770f2e1c1308c2becd0774080ec08d[21]);
            I2e17b8ef0d25ba5beb474e7007ce1fe5f99f6f7cbf24e5241761880a551f3c12 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[0]);
            I7cc2cdc76a638cf4fabcdbd60142d7e4fa11f11486c85b7add7d4f9ba16042c5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[1]);
            I03527e99f5c488d7864664f339e2094fced797e4b46101f3c2bbe0b892c2d299 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[2]);
            I9c110ac43d6a359d54082ce347cfc9885dba985b743aeb66bf25962b4539a6e9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[3]);
            I44089ced0a31e79af650baaa02274890b1f60ac7398745a0e4da4b2242f849c7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[4]);
            I1308b215c5082a0407de73f2273fc035460ca21b553479402290c244cdedad76 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[5]);
            Ic0561c97824b9d5b0d84c33cd05cd4f95b9cacab06eeb5e022b0cecd043c6a75 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[6]);
            I533b2cd0b272eac7c3f9005cc355cf85ce73803134a0fe0ec194628c3af0ed91 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[7]);
            Ie282d05ceadb0d075cca024b7311a5e477e903295d7928735a3c338287734846 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[8]);
            Id8832e8e711bb3e7fe9136084b9832a2677803cabec7f2469144eb3b6d4ee3ae = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[9]);
            Icefdcbf9ca1f8e02b93f295ed8dbc43258b29cbc0cdf9c9ed5fa60117263d502 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[10]);
            Iba1a21e329197ff5e399aca440cec6d6bd3d9593c332cfcba84d52d541ff1ae0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[11]);
            Ib5a93c88521f26a686316f032821a4e9540fdd8e93570ff35437df7522d34ab7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[12]);
            I91c159ee16a42dcacaebf8cdac4c59d45d2e93735cffd86620ffaf2b859c8795 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[13]);
            If7fb04f8e3e8eaef8fcc0486d12d1e37a887bcdecb366c1e8b53a3e1cce0637f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[14]);
            I6dd215113f113a81bfa59464b587ae7c95f02c1461664fdb818ce751c240b96e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[15]);
            I08384d6ff32b692ca710ac4170d45cb5d2e2df509bbc473af140dc50f51fe46f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[16]);
            I6159ddc580c73acd6e2391f4c6cd9989ebaa8947db61972e4fb97f1e12efd17b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[17]);
            I88f1c4536adedb4ffea1b595f5fa753329c4aa2187a3245269734a18a122e189 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[18]);
            I6f52a21dd933b23b7565abd508c69070b8cf652dc313689f62c7f04d7acb934b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[19]);
            I0421a9a7aa72d6f574071ffb4c65878f997e6dc2b605f0d8b351358b08c47ce3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[20]);
            I60b41ade4579462091cc59f1faf9f78f236a3bef12f893facebdf8e6b00096e7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4efab1ca42349d81499a863e52d3fb5877e6d4ddc89ce9f883ee51f06d72fa7f[21]);
            Ib5d526172ae46c2a06c11e15361cb13141d0ba754320f60ce6bcd97a9e495221 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[0]);
            I7def9ddb7ba2e414a44523f17bbff45806f0100ef624a52e91b03022877a7771 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[1]);
            I305dec30cf8323b9af4b0a6d285a31b3f5afb2e79c1a2ea77ce70a4409a7c765 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[2]);
            I8ae4ec097c879009d8316e76b0a2ff9f4228310728d8b4dc196543a3976d26e3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[3]);
            I123e1ea1b1588abf2d5d4ede7027783bfb20d60ce3fdf365b86c9f5c84956a72 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[4]);
            Id9d184571e769ba27b0a5a10807ba8da3e6ba57ed7d66aad1cd984ddf5cbcbd0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[5]);
            I05782c612bec6ce9c2707bd6cb6efd55e1da4d234be502ac88cd02453c61ca60 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[6]);
            I0549cd0fd3abf1658d503a09b0baa63d09b1411eaa524e56fd30b12f8498e549 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[7]);
            I19123fb30bb6e02a13f39e3e96af227e63abb1351e53cbb91b8d9a79be96053f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[8]);
            Ib5d22b614e704f01c688034adcd70603b8e69658cb66c96fe3ea76bdb323c222 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[9]);
            I886fbef883afc3146952de2fc934131aeb38bc2134c096497981d303594f1f37 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[10]);
            Ib897fb3696e7d68b81ff3c1573f5cc234d32e10d066864ec203487a8e56f4ece = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[11]);
            I5bb2c70350634acbcf64debae260225ea2ef5b67ce5d03f38d56d3db9de687f5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[12]);
            If81604260c143a45d248461563d4d94edd94bb71d791a637dcd30c5c0cbbb965 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[13]);
            I0806d1e2ea1771b325ea80b71fe9223f495a3831a560f579401b4e94b6ed172a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[14]);
            I9075819cc111daeabcc2ddedb4a4297b1a42ceac8b93213f7f76d0fe87c8c275 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[15]);
            I317bde7e15c3a4d1456e9653a45d4d574509cca539be5c064af2ea89db634f45 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[16]);
            Ice9dcc5d9ccd6caf90dda22be9ce113c53c7eb492cfd5e0b237da4f92aac2d7f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[17]);
            I54b0290e037c2111cfef49e6b33d9a3fbe3e85f8fa8a5c707832cb5477f5c0f1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[18]);
            I7925970ac367f8374fe02f6e4c8c339c58808928696f0acaf85d96fb3f202f00 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[19]);
            Ib398240cd12e68fb5b3ad4842123a4a16f27cfcae3db8bf1f38de24b82e272aa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[20]);
            I9df56fb9c7b812f3ca5949962100efeb5889d69ff60754cb4eb3e0dd18376d45 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[21]);
            I93f4f945a6dfc45c0a002e0bd9251f56c68570c71e862e222a853f8855fb1165 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a28e9d42189ec8b8fc06092da9a6a167c4c92672de2df8c119ea357bbba8c21[22]);
            Idf3bd173aa5e956e898d5800f3317a1ef71e334901db42b94f9c6aa41c87c2b8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[0]);
            I7b25bf7d9020a7dacab3d15cd039a86780e41ed33520f5272ee788252efd1b9c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[1]);
            Idde70a085816497aa92518899b882b67eb7989897509c445847e24204f5e978d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[2]);
            Ied43949ed7bc9c0c92af912b9e283a3e674d42242e0fe8e3d9132738d512fd23 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[3]);
            I18e4b7dc3295cc6f5968878bde7abe5447cebc77dce83fce47db55be2237efc9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[4]);
            I4a91f2655f96c11b03fce33601bc8f71a0fef4dc1782f7158126cd8cc5a1d690 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[5]);
            I343c495ca033301298c16cbb81a11a7f9d50dfa8b93ea9226caa182c6fae8737 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[6]);
            I451de528c384521cbb78ae32b3d4640b0cb8d507c10e11ff59a74a9caadd2117 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[7]);
            Ieca82bcdc6bd68dc2a28a3b203d8adaa09f89fbf0df6cacd8656b54b141d758a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[8]);
            I876c143c75e838720b2a1ee393f5da5ba08822ea13fa1ff459d68d7b0c0e5cd6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[9]);
            I88e5fe043e16a274d915245b02d2094d05fb7710f6078dd6b33c2a21676200c1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[10]);
            I101eb18f34badddefbdefe0c2448e2a8a243e4803ef3244b25365881bf227145 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[11]);
            Ia249a4e7b5c5f1f4458d969c346e560a28969f33c9b0371c6bb21776d319afcf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[12]);
            Ifd8d2fce7b2a1f0fa487e5be6c007a21b5af1d79da5447d461cd37c189e43561 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[13]);
            I840289556d82218416d7f8652d40586181f7b4ecedd132450594aac1bc47a081 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[14]);
            I98ee0d4994c76a87aaef2967ab6cb88af05ab0a7972d2dedbf115ec19c426fa0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[15]);
            I953a4a4cbd4e6c0ccf4880cec5c947f86d6542f9a7f125d7c8cd71f8665b9ddb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[16]);
            I908d977677aa9b15536027b54cf497ddb8741b339748986180944418fd848448 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[17]);
            Ic0fd25473d5639721dddea090dc037e39e4a0c08776c0a343408dfcfc402fa99 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[18]);
            I46777db6f6f68d76ef34c4a9c585ac04e8a978663fecf72d2dbaea3287dfea2d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[19]);
            I4a4338f7d9bbbf60ef4dc6e821d22619911e41300b49e83d57a0a959218a05ae = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[20]);
            I5cbb1dce1049c737c8e052dd6b84121d353e3ee02202bcb8e5fa27261029c96d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[21]);
            Ib4d2bee91a2ab56208d3d1f484e63f085a162ab9d482690dd3c5891a2a34d808 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89bf7999ff7ed420b16220504f7b91a8e876f1993754225e69b111cc51f08b90[22]);
            Icb9b19c9fb878af708bd3b433b656104d0f1ae64cb5d5a3f8dfbac08da1fdec6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[0]);
            I9989d555a1c808f108dd152608d93b00d7a396de9492733ffd5165700c869840 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[1]);
            Ibc813c005ecf7c077ea48779116cce31bffebb300fab262a78d166c4e270e3b0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[2]);
            I58ea58692cbfa8283ab19d6e609fe472aeb9da51d3f3616a9069eacfb18b0bf7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[3]);
            Ib2fff9999fc00e81b173cdaa0737f3e4f711ccd0034a6611e0e9111acff3893f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[4]);
            Ia441ac067e28123cc7cd9d005d0f5a1628da5628d4473db60d61b85c61e8d9b1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[5]);
            I58aad5a5682b85bf58d67b9b00883f015e4093979fae9138f7dcd813618e26dd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[6]);
            I511b38f7ea620301cc3bfa759ab56a2dac9061fc83fb1281673a6cf276abcabf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[7]);
            I0b2c4982c217189306b4f5d3bace84daaa25f2bcd089f5de092f9a7900106c6c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[8]);
            I3dacdb67f2492ed12375b671dc593349c75562e936401def91b4391c153fa572 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[9]);
            Ibba131ee71ced96650ce76aa4695641a089046f8b8345ba312d6868dfbfb2787 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[10]);
            I82a2a0149ccdf627e13b7d422945e626fa268c22b3c30bbaadd0a8de14ddcf32 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[11]);
            I7efedd1a063df95cac921f7cea9ceea1ddd1afd3a70289c50ea2a4807310518b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[12]);
            Ib91519b86b75cae1ba5b32dc531cae021a01350f4e184d39373bf5553f89a7f8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[13]);
            I58cee4a472b2fa2f17266cd6ab55d475f304bbee835aac31ac7879d77b8a23eb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[14]);
            Ic4e32c1234be0a530c66106794dc1114e4c88611be106ffde42a7ae486560ae5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[15]);
            Id32cba1cfd5a10024378db5089213ad668054033f8614d1ae09b83fd483a25de = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[16]);
            Ib0978aef78ec9b21853831a81aac1d87a2410594c7839432302eb5fa99a4c0ca = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[17]);
            I257c396883faa57c509e7257bed0829f9ca51f30a1004ce730d48e1e5b40c0ff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[18]);
            Idaa2e762bb01a89e36234967b22cc76cf290937df9295939bb4c4ad08cb8413f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[19]);
            I9d7b0f41f5cd73f907351990b23117fcaae4302a36d194e6953b54d40361f8fe = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[20]);
            I8d463b693ea969ef3023c411c0c9a1fbc49f81d348282c031b963bd8ce0527a3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[21]);
            I6822ca486e86051ea654b41b63bfefc12a2218ec87a88d8b5acc3e3c8a604c94 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I53199b89f6c649dcb1f3456cae01b0d115065c6db28de7d89136b2e1b2d36179[22]);
            Ie515c89eac4b602d36f70f52a3fd62fee155da2eafac9c1b14bf1917b62bab44 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[0]);
            I3464299c3a5abaf050c7176e4c0e17ade3cd5d6d86e82addf3e12d662def2b86 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[1]);
            Iefd5db28023cae3483fe3f0f1dcd5e302d642a0b5750cfa9940a9a8d6326cdb8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[2]);
            Ic98b2baa4c4b3d4541ae5e7f9ae0b032d4dee98ebd73901690f561438ecfe5ce = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[3]);
            Ie6d2cd42fa78c1cbf17c7f18dfb4c0cc5f79f1fb0bda02dc92192252f99dd047 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[4]);
            Ibbcaf468c4ded9be4d2d82d059bfad5174f330444c98aadb71831769a32f70c2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[5]);
            I17e36eac60eec64de05cb738d1e6055086891ee6fd7d8fb300df4f98a3405276 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[6]);
            Ib8956dcf80473ed75d04e9fcc74400f54ee0b840fce7500bcd68ea6dac6d4473 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[7]);
            I873ab672a8d92c69b75cd8e627aaec129f1cd371c9f863a6bf88e3965909a6d6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[8]);
            I206a4b82a444ed76c846a17eccf6c9ad62c42263b472949cc97f838f6a416073 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[9]);
            I428333658d20f4417e24a58fe364d5a647332ef76ecb7f15d83dcccf1aeb3d11 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[10]);
            Ifc4886636576352e5307fb1fefefded0d693fd059a3fcdd6b4c9dbab1b908114 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[11]);
            I18886d5e45fe8011ebcf9a20aebf875a01f1b793a54ccefdbe44a896e92cb0db = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[12]);
            Iecd27d9347b5f52e83b7d0fbf7e51de4a3711cbece5ee265b12663b77b58914b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[13]);
            I5246ce1dc41e20a5e4e3312a997e8c5be2d733f0cc95f74caa7e668f9ad2f1d6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[14]);
            I668775bd016b2384bb3d1cb0a1e89a76d2af15b2307cc6a5d2e0d6c699b02544 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[15]);
            Iaad1ab5e7603d5441b228c5e899eea7781b6f486b836a7b662f38ea832c1b8fa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[16]);
            I9d56c14b3465733b5c5fbff528a7a7d85c918a857257ba8e302ae84a0f4734de = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[17]);
            I7ac4d72123feb2b9af1a6c3da5adba445042363194ef471c8761e289178d0253 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[18]);
            I7addf7487638274202ddfd183ba052556f89f82da9e873224c5dddf27d2d5a66 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[19]);
            Ib0de9295b071389ca7b6bd34f7c9371614337b0be04ccd9ab9819a8e39ade463 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[20]);
            Icf6cba7551eee2b4d2b53263af6fc190558f5b29af52c060adf5bc9116d56341 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[21]);
            I01a734e70411ca4d260541915dfb0aa0eccbb88be6043a4a46e412d3b9f1e778 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie87e615bc0857b050469ad82e505ba2dadd16b2cf3d4f91879462984121d1d4e[22]);
            I04257aade4809f3b60c5cd618c5a29008d1b3d7041330bd5c8db7df720da3694 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[0]);
            Ib33ee0ec338d1389ec9010793383d24de32231284e86a9b03fd2902743dc8a00 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[1]);
            Iecf3e0156bbf76dff96948ab7bf67772773b6bd62bd0e0fbc86a6eea8b05d4e1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[2]);
            I80c4eccc6e6be84f8936ed3e9a9457a862eca015298ba2db70745f25a65a6571 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[3]);
            I7355df30b826dd16e0f1fe3be878df80c2ca672dfd1392e2a81ac34fa3df69ab = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[4]);
            I8f671fbd5e9e240cc2f3a9c60c1340fb4bea46c25cda7ea5e42c7ca0c2360bb5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[5]);
            Ie3806d0fc4177d813aade41ad46537a9a335516135161cb2ef18ce822cb301aa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[6]);
            I8e8e17839b8f0cf30290c33a60662c784f062950716903854e36856a58f909b7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[7]);
            Ic46278073f42d4eba79499cd6293cfcb33a74310e7b2ed4bff06f5cc63dc9ebd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[8]);
            Ib1101385e86160606eeb12ff49ee86ca465f227b19c9bcad4811c6a0183c0ddc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45693a666ed22a35f933f7f0593f4c107dade2a6d7168aa2cb2d237e52c6dd6d[9]);
            I4bfb42a957ed14280a129921d4d635017b23dab77b121f51abcc5e738114e446 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[0]);
            Ie11729721562e4a52a189a242aba934be636847d35de867cf00d26690c69abd0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[1]);
            I84cdf374f692a63dab22cd91edd4f71e1aff29b51b06f0bca914f92407bea09d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[2]);
            Ia2aece9bdb39e997b99e491171667091adbee475ea9b1c372ebbec109f9f714f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[3]);
            Iabfa5de761b3413904b919f913ed73bf27f5249b7dc6bf8471a23f06a30431e1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[4]);
            Icf6fe11d7e6948c0bdb9cd50a0135c3b0fac213aef728b8a6555b7601c51cb7e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[5]);
            Idf57b2bf209c68bfc70fe2759595334fabe3d50dcfc4fef8637586c6623c9c29 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[6]);
            I31ea69d26acd05d303178076eb123a7b2bbfeca82c2690c54323889753261f1d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[7]);
            Ia84ec437292f1ad3e702b4fa896a4f545cab7253574d294243af0c1e7de47155 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[8]);
            I52cf6523f0dd5f666334b2646768fe4499c699c8f6b27ec32ae325cc0981a515 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b29c4fc7006e02fbd94a82ad3d166189d6da734c66e3ab53263a5f62129510d[9]);
            I7da5ecb7bb8a413a5c6c51f0aff1921be97bb5df5d56f6648c27ee4196fa93db = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[0]);
            I81c612bc8b32254693a4a0c89fb21865b161dd1673f5610732b31dd5663f160a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[1]);
            I5b143cf694d99dabce0cb40d2d689fd7232531ab3a30888f811171b6aa2e024f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[2]);
            I050437a5474ba60337593b28d17e2bec5c76d26ea8afeac61be93e8ba0ada42a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[3]);
            I0442e99f7519b58fb576a898b41563a174beef69bb6a525712224f5d767a5867 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[4]);
            I4bed271962970c26ab72de275bea4b2fb0565d7e44f15b2a1df631bba9e5d4e2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[5]);
            Iaf95e616f53a061a7bf59bf1128d2cf6a5ef64d24b292671a3124a6e010d964c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[6]);
            I41b85a49eea9c0d773ecce66f0023338d3ee5a94e14a87c867a74960d30211cb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[7]);
            I3390b463514e772ff0afe74698bc4850014fbe363d105ce3d0e8810706977682 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[8]);
            I3e5c11a25b8726c787dd0ffc08e93b671baf84832d9413eb7031a6fc17e8ad76 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I817c5136f126ea0e185c3fbd01633d41751ac90a1a2c2d1f2dcb3c7d0306a765[9]);
            I6b499c648458a2ed0cf0b27d81aeb706a260c5615a8def0ae89a1a44693061c5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[0]);
            Id3bae057e39f6549ce13910da61dbb41693ff87efebfd241bd1410d3da7195ef = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[1]);
            Iecf240e8fe5f620bf43121455ba23a715b23f53e049d2a36f4bf52e2a061a8dc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[2]);
            I7958c747e1ef37e2995c52178d143af6a5f3acdf7c6d1cae518c82653ec18716 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[3]);
            I697a55c4cb2dd56ce91465bb6750d05200607607d7eaa0b27accbf7f20ba97c4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[4]);
            I2785beda1166504e0b7ea979dbf6c2c5574159cfe36c60fced2dc64ebd05a9bb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[5]);
            I0b60295163435ae3d3b31e9613d753e7e41fd66c11fdf2e7248d7864e11d9d84 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[6]);
            Iccacefad631e33ec8e54f8261759ca110fefaa6fd9fad08940205708a7180eb1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[7]);
            If07308cb71758beb15e4a33e3770aba8021bd5572128b9bbc1c8db48e7f807b4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[8]);
            Ic2bb8293812351030940ea0e0a882994714d60a4963e82e2291f6f2d386fce8e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2b1f6e92dce73e19160f1d26bf6739ca3aae17dca6d93a709c0ca72990fc160d[9]);
            I83ded8cd9258de3ae8deb907ae3b813cc228b189df92f42c55a4b0eaf411c106 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[0]);
            I89ca3ef99e4b84441ed3cd9f386109125b6da2d23485fc22513b1d8ded87f894 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[1]);
            Ibf9f290605da4b6295c786c6ebc135cffc80a3352b42e1d841ba5f6fbbf06cc8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[2]);
            I0b2f8e7646b38057090faea20bf55e51f17d23baa4daf0c16d00e75e4c5f0ebb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[3]);
            Id2dbd07db2080c14fd0026396339e31183fb5bb6a476999102300cf81f34b93a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If2b4887a4db3c634279bbaecb72e3bbec2454912bcd7907e12039a38d6f75bb2[4]);
            Iba5fd100311e883873db0c3474169654308059bc4c43d52479a4515fa85e8900 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[0]);
            Ied8c84dd66ab8e8fdeb83c6156b8a6f8cbcbee27c41ccdd8c4d199f70ea67e8a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[1]);
            I1ae7d02f524c03ca060c3dbc879653486c099ecee485690ce40a355fc1ed843a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[2]);
            I43bd10e4f520ec08b30e8474404cf62a6ad869cdd1d280a2d221e0d76f228091 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[3]);
            I7e12dde03af7a5ae0d05cdc9b29f31ef726c7bc51a7f07e374bfbc0846a24f0b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7e87f9075f32a59cb7efeaf794b369432ec9cc0909ae5397293853038542591b[4]);
            I0e7725af7e163a3f4ee8bf63bcb825b6d62f4b9260a7c68d0beeabf35eea9391 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[0]);
            I9a798d59823ac9a032d0daa203a7bb153e483bbe4fc47083c1d7e4a65e400156 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[1]);
            I453d1e19585e0fb4fa66d684f0e6b37f56990cf101cc3942d5d4fc7e2313710a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[2]);
            Ibdfea3d72843376261dc3e06e3f19be4556508098d1b4d37c1c4cf6928860719 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[3]);
            I39249b7f0d22c6116a7dfd0c0748123ebb6a9b7f931a492a534702157ab28c3c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib0b9066af0f6de889b295a7145aa315026d590fac11c49f8ab89a27e76a93e18[4]);
            I1ee3ce036ac0c878003d846cdc3fa9f6b5854855789ea575f0005a9c9937c58a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[0]);
            I91c40ee5121cd738ba7213df9bda6130b101385a28d8a5fef6544c86f6bd1e3d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[1]);
            I465489f86885351586de73a0aed556821e0ce34d1c2cebb67227004b4503eb3b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[2]);
            I37646f9ba79338e88c3d793a27911c88d573dc5c1cceaeaf565606c5b61495b6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[3]);
            I8e95ffa3fdf70dc76c935f7d4dde6f39dfba8eb795f7ccc55510ab3caf678410 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic77a9e7075cd3684473c2d61515f3380ec6428a5d16b3fe8e4314bf54e3aa9bf[4]);
            I592170f431e8a8e15769fe2e5f3bc43a7c514290149bf9b93a8f3d3a748094a3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[0]);
            I2fef37935343317384b1d29a04765327533fd87d4fe82a74f24b8196b3dffc92 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[1]);
            Ie57f94a45eba4db3826b22e3eb6acfcfa04b6d0669e22e5b78dfae4e7659b205 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[2]);
            Id5eaf1d953b17df3896f9a30f37363d1a69fe3a956b97d307c895065ff32674e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[3]);
            Idcb8d71f1ea9d314ae8f26e9f4b9e25ed245bad319b9af2f71b035aca6d8fa6a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6469c3a9f97ec9d2a68c601c692146a7d9206063925890934abc8616a018aeb2[4]);
            If307a1ee8e5164bac03971d07c03c3c0440857c7cc29df11a751b3bef9bb1516 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[0]);
            I3efcac0fab0af81582237cdcd612c8d22eef1a6534816484190db28f3e7f3a96 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[1]);
            I3f5dc950ac82420b73e1bc98c8c412f7e91958fbf455413c6a0ea5b2569e078f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[2]);
            I42ba6c66d951bbe03a57fa7a4926d6323f30784fe87de73cce065cccaa9814b1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[3]);
            Iac102173e8323a836c8f86d266f551fc24ccd14aaf39c7d9ef26c465d38706ac = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic41c580448af189b1132e135b464fb2447c1fed455dbbe461ec09bde73548dca[4]);
            I2976810df2af0dd2879fac8afe975126944b2e40a51dc7dd169051bb5086b3de = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[0]);
            I9c3d0fe7d767050217425eadb8e780e5eeeb31239f2f517ae5d122bee4157180 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[1]);
            Ia7d01a6ab6c0646f75030a0bd04a711a9c50dc4674c921680034012e67a0c3ea = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[2]);
            Ic8108e830a58b12b8e3ef4897cee70758d1539ae6609d73b5455b94b0eee5510 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[3]);
            Ic96ea379edce04b88c524fd17a2b6fb2283e45735640aa3d8ffc7f1bca77c78c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I928da3c238e63d326fa5d7f860b061dfd048bc29dd9fb2ae595881335c7eb225[4]);
            I4c871d8c6a677ef8fa6c955524def78e8df6f9f3fdafb141d43db76d4569104d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[0]);
            I6f7a9d597443df1a96370dbd5e1c1f9cb563fdc4db1d00fa66e8a287fca9bea1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[1]);
            I6ffb18ff0417e140b26d84cece8d23ea507516ebb60dbee4438e9433713c9f81 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[2]);
            Ia187792bad45afcf25df25b18a076d255536e94db8d7bac4df79761df5f16050 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[3]);
            I9c0a341c77ecbc1b3c44afee03ccc5a8f34b1275db9c439eedca9ff61a1a1eac = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7dc7d464b862672ebd31b6b219429a01a6ad790a9b801425f8989c208ca01d8e[4]);
            Id8cd2e026867692af509cd433fda0fe6a8b5ccb8ed91bad6530d14172dbf7375 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[0]);
            I2ad4afbffd2865f5c89feff965381fdaf73ac9ba4bc6e802a39014fe554b09ea = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[1]);
            I31adf91b5f31b4232ee24f82af27e02a7ed1f8535c552409f353690340b64b2c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[2]);
            Ib96bae85b07ff95f5a6716cad97c765010937888a28ad63b16eef3b6ae93b3d2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[3]);
            I91cff501b877ec0153cf2d85abd12870d65d1aa997a6bea7d653bf387813998b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[4]);
            I42295332275fc6fcb94c042fbe6b48d3d03038fc27c535c7e63674f58da60bf0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[5]);
            I445cf6fbf071cc76e6fc981d7f2f201d0e09d3f47c1227feaac47fb57a14e85d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[6]);
            I96ace764b2f8db5049595445104a408a641999152f2a6c63d22bc6946c27322b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[7]);
            I8741cd8af2f9c3a548c5c39709d7a186f0953de5af6d09d88901e0083a539096 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[8]);
            I97a73864c1c919943cec586befbb524fa6d6da6a60e1503bcef8116c646b71a0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[9]);
            I0e4ad715cc833c775ed97e88f28c4196d28bcee4370205307f4266e1fc572cb1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[10]);
            Id1fb56c160d418b26fe2b51dbe78addbbd2743e7a342e0b6bebd2e8d3cb1ce99 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[11]);
            I20a501f960ccd425135a3fcb8e667d68940a5950d939bca37d107d479984c038 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[12]);
            Ie28b77da5cb0eae41811ec7dbc5f86111d64b794121eda9f2f0515324579f844 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4b50cf0377a09e70a4d8fbb3d8cd31f203078ab3467cfb2b9cebf1026fe5c9a7[13]);
            Iefca48dd9d0f3c717b0a3b081894e93ac451ed275f3cfa7aed675f58327a2d02 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[0]);
            If6592aef798f1b26c5c6593d99137d00bab8e8631070e89dbc6a3e11c89b3e92 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[1]);
            Ie14918150ed723163714038f6ffd2c64b07d62079dc03ac8fdeacde45633def9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[2]);
            I5a03d267642091bb2d177a6689d91b995983fde126d703c6474d730b455ab56e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[3]);
            Ib6dfa3959980c5d348630e2edd81fdee8429a3003b0a21369b99343bda03e2a0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[4]);
            I97f8487b89684c5c6952770b0468738f72682d6230be6a5a31a92fe50bfb239d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[5]);
            Ibca42a442c971d363e4f848d203d2782af05ddbaad93e8cbf334328d94a8a499 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[6]);
            I84744085fa951f13f4fef6c44fb0180e543fa6793e89f4dcb14c3da6b27105b0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[7]);
            Ibc54f1c4736e5a4608208441ce8d81831a0b6c7448083d6e6976981f8a38d1c9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[8]);
            I211a150dd66153a3c2c72be4c24145e4c9f0b2f9a3032fee9233985ca9d2c4ae = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[9]);
            Id9a38b1906060dc5739f9446bb2dd1a6b6603924d4b7889c931988fb52cfafff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[10]);
            I8beede7aeefea570e5c65a76dbc5ce1f4eb114e444ea9b4636258bcefd9d5f34 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[11]);
            Iabd5561747d288862c0b289a28572fb5b0159a3fff7f79c59bf60f1612ec1e3f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[12]);
            Ia4205a1d01cb014ebf8e1d539dbe1c7270bf9bfa8eb7920b136417bdfb9f498e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I319dfe12017051baa9b3e6f7545e40751fe8fadb728290b8b60534b29f1a98f8[13]);
            Ic45f0213074aad63c68cf3fe879ad5b0e70a5977f282822ab582ab88ae7236bb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[0]);
            I123d4c26243478ad4cff3406be39503c6b378cdefa50bf60249ec03d3a44270f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[1]);
            I0f75d5771cfa314d28e188de297b4bb53c2cb732724a630e10580ee5fe87cb23 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[2]);
            Ib6f695414c34a124de17de5cee8798a33f0968f7eca5143f21f88c228ffa6345 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[3]);
            Ib43a705a217dd9f2321c3e61ee116d257d8ad59bff5b4f80435f9dd96a8d04fb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[4]);
            I3e014fe75658214d8ffa60f966549b131bff6a16020d7858523ac829b0126838 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[5]);
            I31734ccacbfeb8a5c0c30cfc84934f8d1636ce4ecae14fe7809d6aa8df35a9e8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[6]);
            I701aa61e04d2787a36f529185ddcc94c832834d38ff92b37456b64ce46c69b2e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[7]);
            I4b9dd5299690e88d870ceb4939b7f8fdffc8419431458851a3691de4f78f9f15 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[8]);
            I81b8212f2e15845be4d129b192895f659d31a061a3a033bc3ac9ebecc75f73fe = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[9]);
            I1f070cf569961de917cbd287e7b14a2ad6e04a4474edfb92c095f6e9cea1efdc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[10]);
            Iae16b002804d17ac9e2c9655dda031f3f0ac10d703bc42079ee2a5fd3ede604f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[11]);
            I5aff0a6c62deaff6e9d15280ae8c3cc326ae7f9ea6959dfa41a92c770b592cce = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[12]);
            If6fe8b42d897a8c92c628edac7869deee179622fa52fa779f2d9a0279791afc0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2caf915b3bd168bacd35fd2f40f595e58786d73b55bd518d5471dc002e4fd37d[13]);
            I10a223d797492c10ad8f6aac1cbdae83833e701ae6314ed988ac117debc98c33 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[0]);
            I8cf1c2115398eb404050fcfc654b198694d3c54eaa592d0d725b15e7937d8cd5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[1]);
            I6ec1c8ffb963fef21e978fcfd0268bc24dd283819081437974fa5a06caa64c25 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[2]);
            I781bae0d109036c417f71e00a3df3440df3cecd691fe1f67c147c4d2de217f7e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[3]);
            I10ecf0f58ee2fd15e2b4135dc03cb4053c364660c6d2e2bd03cfc37aa6d6621d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[4]);
            Ibe646b6da0465c3fb411afc4e03d45f553cf91e67cbcd46674a0051ac1092e30 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[5]);
            I8a61ed94b6198131fccf4feb6be7327f59408e9de4def9c4a155167192c5f065 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[6]);
            Ia57f6e4dd9ce4389f90c78df4fca73a681df346f58a85f61a74e842427848347 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[7]);
            I3d284d86f6c46162d3e0f913a5a6b0e1f2e34fc7ced6a0c226d5e78da81a0633 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[8]);
            Ib07af5e0c881985b1aa0698382702f78d3ec7ac69cd0deae7496bc63e519a738 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[9]);
            I332737561309225f302f64e49e8b3e4aa4dc35344858059b21e146e8cb84a466 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[10]);
            I7e3620302652666ddabcd16531a36e7af51722c39bffc4224f256a34ca33109c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[11]);
            I6c8cd97a5a950e00f0b9892a96d99ad1e5bae6c2db215bbb532060b753233aff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[12]);
            Ice95c4df972e8e6a31901269a2d291a70fe4e8dd1d86ea5ded5a16cb1c169890 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3c32fdfaeb2113e4726ace57bfbbc7520fcbc5a37cf38a2de65b9a320f243169[13]);
            Ibdb4937356d2b1cd2091a695635cc7c69b694f775f4c4e8680ea49df1ea6722d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[0]);
            I95e467521db517b858e59156f95992ddc522a7d038ac6bbe691a91b567cd35af = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[1]);
            Ia9160306dcccf07d591c6c85cf86175408905d5e1bdfb36206d9c4bb5b917dc4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[2]);
            I207af234897ed272d784f4a9f8850eaaa2fbf47f583ed1f0564201e33dccfb66 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[3]);
            I0738f605ff9ccae9ae63f8e6fe7a9b537d97e13bf3f23c7b0daa4fc414eb7eb4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[4]);
            I7c10e2245efc27a4e2a96467eb4e3fd9c28be5f26f65c560653ff4742fa5143a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[5]);
            I00e08c73bb2036cde2d53598b9977dd2504934b9ba8b58bfccdd21adc2fd223f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I771a09d1a87e006262791bb9181c8a350f92d14fef6313b3ee7c5474ef49b778[6]);
            Ia718f1fe0157bb564650d817f5ea7960bd0698409dd04d9b31d54c95a3f90318 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[0]);
            I95b908a4845eb4b14e8f933057bab27e44c6a867e4bb02d87417740e3150e018 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[1]);
            I600d6bfc6bdecb80f4f9d6020bdba9b4c04bcb359e66e793a3bd6732173d0b17 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[2]);
            Icc13ce9fe63ee1c11fd5dddbf0a294cf6ab7ae703f742a92150b7a77868a5a16 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[3]);
            I2fbaaffcceb2dc6a4f6d9d34140997b18356dc3803bb0a6c6d5f1b3f980e18da = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[4]);
            I3c91639fa462a2a7e65410080b46408b692ca4639ed17637b1d465f38631734d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[5]);
            I3adad3708bb709ccb06c77ab54c92b6c6629853f740147fd958e6200aeee81bf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0040ccfd97fae3ecb6a47df4203aa6b419c8004e0751629b5068f8d31e0ed092[6]);
            I706a44814e015449aad217d9bd9e0056813b075d8e622aaec4dc08a3518cc0e5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[0]);
            I18e5d7f94022748f9a5645c2b0e385407e0f00d6f9ab28a55982fd36330ce524 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[1]);
            Ia0090ea9b75c69dfca34ac43abee88b20734f7afb9c1d88f95eda3df6aab27db = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[2]);
            I062483fac022c2d74cc4bb84d57c636a3bbb67d68dacf0da453e3b5f71ff8846 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[3]);
            I15ba9fcccc2e3aaba7bb5967d35eeecfc3bfa7ce27f82435be6dee9d0a4af829 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[4]);
            Ic1034fe189ea09f2aa3b69428828a2b7dbfe9389dcf48dbdbe0f15b9157f7c49 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[5]);
            I8a3c94278b7c901702cf1b70e89c1832afee395077555d27badd4e2b6fde0b7a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib64c4ba9b97f1e695d955624c10e97e7a1dd7866a4da7fcbdc940a5aa03d9f7e[6]);
            I23d075a3ac353b3deca0a572e9cbec9b1ae24ffc7f134b36c6f938d949bdcb1e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[0]);
            I3599299f7f89ed3c6b11b31caa26e6b30553b9dcc1d5968283085959f822a4c6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[1]);
            I8954b3335e6848eaec70a960b632233aff75de56bd0bb895e2b4ae49095fe19b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[2]);
            Icb88d7eda8505d92744b075a1c229e3c0f6a9ff062bf5cd35f6f84467b451e9c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[3]);
            I20ac47b3e52f25ce7858fb7952654107faed4cb5cf3abe1ba915710d1af4c933 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[4]);
            I53a66c670d7345059cea712c026fe8c524e74b030af0de054cf6e053bb304248 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[5]);
            I034d52d03f918c91bfc6236c72b0d40b688e2bd353f9ca1f03f4c61449bf128d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I352169a0053c41f2b24e1b8eeffa8bfeb3d8a8441d33049ddce36e9e566524ed[6]);
            I727007bc323c90e0c264e5b8688898c0df1bb72c976fbc3513439c14f15b5733 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[0]);
            I0011eafd50b7df59be2a4f143443c0ca8ea87f9a93586d07292ba02fdc2b9b4e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[1]);
            I7f3447e248449854eb030c79bc32b602d376441a193e25bfcf9b8a0eda83b57a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[2]);
            I288ddea916663f74bb339e7a94ac9c86412f39671ca69dc7ec1da05a1800092b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[3]);
            If023ae056e9b4b370bc83a2d5604602f45a01a005bc19a769c874536faf4abbb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[4]);
            I48ffe541268d63545fa48263d8df3c288af7b2646b4dca546a4dc521aa247651 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[5]);
            Ia81ab6d41925460c11303075dea72c7fb3fe533d88450c32414823fc5b10bfaa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[6]);
            Ia7a158b91a24000cb6211d129d65e781a4e28b8333f897bb401042fbe17c37a1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[7]);
            I698aa30e42ad4f250363d29dfc5117677b19f2da0afa75a013718ac5b9731d6e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[8]);
            I144fae9c9898630fa027b3237ed3434c76965eef2eb015effa7c8677b19c91a3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[9]);
            Ic595c984782ebc89b61fa2a64e994aa66eb4979ab1e30e890886355dc247a67f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[10]);
            Ife11a6b34a661bffcf9f0147459d2f5a23d6c5460c59142668ee0f0506755225 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[11]);
            Id73bbd3c91f1e5fe13f11e8849f77aad2ddaa35d1399140ceb5e133da8e11227 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iccfcfd062e5bb23410c6bf82b107b3d0ce0d89d527288ed6a40d057eb1e1d3e2[12]);
            I2d89506b7ec0311db709c4aba53b749ec1b531bf4bc7867f3866c39a73aada38 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[0]);
            I390750ab5fb20d9be34ce0e294c95ca61ab6e511578b636301037a34f9bd9c07 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[1]);
            Ief01c27ce040b3f50c19615a8f5d9bc8b467c0f88a778888fe186887b19fd580 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[2]);
            Icd850fa1e932d19313713c2d376413e7b81faea883442278fbc700a2238f6779 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[3]);
            I5fa215eca11a15c7ad85760cc87a0f8e883d02472c7af460b13cbe214a596c62 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[4]);
            Ic336cf50b44edc74db080d1127ba09a4313c0972702200ac5207aae8ce6b1062 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[5]);
            I19b5f6ad3c2f2551b49883fbab077c8e3d76392fa42a5030b1f832917bc2641b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[6]);
            Iee901b35683b34719c33d63d90b8ae11fbc338a170164aac943fb0b495c92b97 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[7]);
            I4d316d60bd6537dcf09dd9b7eecd93c86af11ddecc1ee65e4b9d65c136527e0d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[8]);
            Ica10d27b8c94c1e740a2287ef28e5d3fedab4221b391b0a3a1da3a472f094039 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[9]);
            Iac3e25273f8b972112775f3aa57274eabadbc2da5eea147328f85a941b959bfd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[10]);
            Ifc38f7d8250994e5e62716048122eabe81722a32478caab729cfb06aacfc09c2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[11]);
            I47b18bf83ed7f7e8a2c69814aafa41a66b6838a5a997d036c634f488f1c584f1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib04b8478a07dc3d3c189726aacdb0df6916ce4a77c4bd1dce00b3d3d2d40c54a[12]);
            Ia9f80db3bd889aa11f43f6aa371715d6aadc7d3aeac0e9519f79b787da6e545c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[0]);
            Ic4c53101c741f07c928018af5696d83f45a29d0e5a9f766bd2f1f1404f3eb59e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[1]);
            I4b15e4ecd6a6f2139463d94eb4061a410569136410e469abc38dbf8cc03948a2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[2]);
            If377629f88304a78a44bdac612907792b54c49caf9dbaf85b3061be5baa2f5e6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[3]);
            Ibb72bc519d54383d213250311085f6368ead1c943881ccc23f944e652f934063 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[4]);
            I91e90d84eae561663a2e9e59f79782a78095807b98187add5501500b8c1cb126 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[5]);
            I7af411084739689195bff036e9d5e9a950a7691f7d771d4d406aba4c32d95116 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[6]);
            I06414f803df7c8e59f01524020e09627cb11f3809c3456a9a64655062b110885 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[7]);
            I4eb359966514f007fea3e135207ab27fc596987f985b8a3ec6bf51dde2ff9e38 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[8]);
            I60f3a2c7d8e3935c04abc8aa09b0a2ef540f13bc98beefc600fd70aa25421191 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[9]);
            I698accb14122caa36f489e7fc522e39188ee03651ef0c6670eecd60162cf2f0d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[10]);
            I49a96e94f51c41ba36bb7a8d466771682602e2dbd6f65e13d7e858a60b554f3b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[11]);
            I79d13cc47977ecb1fb0ca304be8c225a427063b4328cea4c4a227521a1f26018 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idf7f4aa4535f55a76d32bff341d36b5188df8ce756a79bb3a22fd7b8e523b008[12]);
            Idcc1ce57eae666070b5b9984cf69d5d2409ea92b36718906218185325b5611b2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[0]);
            I54feba5563ca84d4a04e3ff7ff5ecf689d26961daf0ce27f0be8988087296fc6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[1]);
            Id60b48bbf346bf95a242f425de7f456aaba5b3ed35cf16a07ac541ca8f480319 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[2]);
            I8e89f3937a947ff09fef0df8085edc1dc09a36d7bbb39027d358384d54088060 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[3]);
            I800a86b8eeb247f39df85aba37dbaa93060858c235c6ac6b0912fca85af95477 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[4]);
            If4b0b6bcc29aecf6816eab93edb0cb358730913253ae72d15db63ae06b19c52a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[5]);
            I63132df742cc353a39f27a7a5a00e0990e9e9e023f5c2a8bd571fcd6dd2d760a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[6]);
            I0734166e34887037bf713bdf1df0f7219241551cec455ed45881734727f90032 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[7]);
            I9f08c1a4053ac65909c96d240c83e15017c81fa41f351b0a707fb7882e49f4c7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[8]);
            I3af491b2352720f2bd378052706f4ce571453d59b0fc78b3cb0bce2d51ce5700 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[9]);
            Idb883f1d90a389f89c3e04f54dac20f205951bba3fd0a00e9432498c4def1131 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[10]);
            I4e556f27c558f3d1f76d2ed4a3f0b1a68d74e5c0ce6370b9eec599e7f76f8bbf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[11]);
            I02962ee90b42f9b95262049bd2dcb7da2f43333787a578d5f5721681773db287 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I45150a7792333cfb9e2a54809077b74025da043fb37bb73abcf52598234e71e5[12]);
            I739fb2ce1dc1a27f40af1c53d575108539718f9d60f83de60531d7bb201685ff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[0]);
            I1a6ae2cf67f356fae1ec533488e09c6696277823378b06751db7ec97115d9c00 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[1]);
            I931537d878467c473ac81aec8f9a7d79f286024e62ada1e5f363b93d6887070a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[2]);
            I61e7244c25e176443b24d592ff4299482d572c1705c3e0a6b44698b5366ea3ff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[3]);
            I3b3f53fca961a376010d1a5b0c49f91d58b351d0306b8433ac22a70f5a1f1673 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[4]);
            Ica809c2eeaf6926552d9f811bf16c30146853674185c2315876fb5b2ea6d0769 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I321a7a2723625e553d5f3b7f161644f16fda67857d69397e856ea39b00bb558d[5]);
            Ie3e85438dc476813cea40910227c7d63eb275948fbd481f56cc51656c1bc8b34 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[0]);
            I877734e2edefa267510037759c9490dae213d2e046beccfe87e16c1aeb5583c4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[1]);
            I8b5d8146640c84b84d0d6bcb2362fd5bc7e7462e1905b32b998b1f00f2da3645 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[2]);
            I57ae0fac4bc1fada55e48ef9952dd7b81a55414196fc22fb27a20b723832aa84 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[3]);
            Ia2343365eee39c9305def2bd744d3e44bf20b5bab8a48c6a2d95908f74f3cd18 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[4]);
            Iadaa0bd11c77d7ea8c8cfc4b0c805c5afe6b75f597b03729ef2cb704dfe48286 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icffd9793c13e01d998b52323008a613f8811c2e073ece0f291c24eb0c1900a8a[5]);
            I0543957798ccd8923b2a5b736175c6888eb71c1466a1e9cc7d7635701e103823 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[0]);
            I87c64e9e81da569414617b07e39a7f67b0b76c71643cf7257b7374feb6fc9750 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[1]);
            I481cb000cdc7a32db6aa5a6b0da57b76f53f5bec6ef93d4ee25557e1b12064f8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[2]);
            I23f5e95dbae4b1223d603061df9b75b9a9ae8409c6bc4ad1fe23d3f5c7a68bb1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[3]);
            I16778a093510ae433495baf9d2b7a74ad4c5315403d0e8aa39eb09cf508dc201 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[4]);
            If2cfdc638b3cfc13d31615533cea59a4bf8123299239956479d3f1d702ef54d7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4dc683cd869884a2169ec5238c2e6550e5fa5b1f3971c9cf959b41bc8819b28b[5]);
            I114dd7172ac111bca494cc4230447a2dc167f12f198288d34cb5311c279a73b8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[0]);
            Ie72b5524b212840dd1e69f4fa41b4955ca028c1ea7fd2f3440843cc2ef6d4be2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[1]);
            I8b151ef6b3125cf983140726d775d948a253c13f020d3d1e75b585afb979bc8a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[2]);
            I72329ad9fd98258074b92a7e88a88c68f8db57e7d6460e9c29ec7f3cc251de29 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[3]);
            Icdad18f8878b4e9645b4f2d2434f913a6e0f732a20a6a750e25c2398a086ac2d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[4]);
            Iaf14e804e3bb7cda8e67e39af906be2c966fbab4a6e73b8d60ee7ac5733669e4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I09ac577d9e4c28035c6f78b2ee9170195f64c2e0207fed3e3976f5175ce39b8c[5]);
            I238b01744b520f8759a7e466290a15b15b96fc95b4b8a14afacbedb1657f7069 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[0]);
            Id29a54af13b6045a8a43f741c229ff88d4aeeffef29065cb29cffbd861479f7d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[1]);
            I9ccd1f3aa9f849bfe7dd9ff5f9de6fff64a444bc5286321a1f0e73e990d6a996 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[2]);
            I02ff320cae73fe5cc67804e552bffba75496861f085869eabab140094a18fe90 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[3]);
            I6eba99f7e39a1779ace2db8cd1806d099e7cf0678ec385baba570209f784b5eb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[4]);
            Id4182b8f05992677e12502bcc058d967481d0dc2c9c4731b657f04696a5b5bbb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[5]);
            If4927b8f31777ef2940c413336113e906e0e3556c31b9b3233107b88b1d71999 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[6]);
            Ibf57f9e63049a49e05739966f1ec2fe4520b2959db6fee3a18ead9ca03aac230 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I14fd7aa04c6b2aa32d5d7897a0eede3b12244cd38980578dac0e5d03b02014e5[7]);
            If0025a7dfd37802d1a1fb43d82ff871c2867504735093f0ffaa8b0d85fcd4d1e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[0]);
            I24dbfd322139e6a1964e587f89b06274c35617e961a5f61f90c67ee3b20ff208 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[1]);
            I8bddc257a28da31b71dac60701bade264fbf14f8377b1f504ef874c72e0d45a1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[2]);
            I225da3a8a67ccba14e13c78ca2ffd83b37ac9a961371f1aa617f5752b1bb337e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[3]);
            Ib9855ec95d5c99f93ad4c5565e622dc1c2d1c4a3b5d0937219172d97ac290756 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[4]);
            I598f53ba5c7ffa41f21af94375843b0b7a911670719edc80705508ae32ac0ddc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[5]);
            I18eefcf5075eee79120ffa0e5875cbe7632d1db84b1c498107413f14b72820f1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[6]);
            I7cd31013bf73ff7f7aafbf06eba3fe8110dc5490a280c2d79ce53c77896f564f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7f43e980f3c42c2641cc52696f4d777ba7e0d4f792f8529a5aa511d4c69ffc5c[7]);
            I804112f16593c6ce81f6459599203b07642485939c898d78e113353659a62a68 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[0]);
            Id8a5ef9ce42d57c3feb442ca091604f1fc51e648a89794ea3fbe4b30537fd286 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[1]);
            I6ec3df474c20bfab5d99aca971523dec8454a5ad4536765f4f9bcb0c31978cd4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[2]);
            I862b7b7769e1ce1579c40d6363e23230c9253630d97fe8abe72b80e8a8b5440e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[3]);
            I1ca12951f309a25752defa88fa366a90a13ce83b7fb40610c01a8c11a3c2e59d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[4]);
            I786cf639910ac9a90b1abf55f9e3b66d87c4bb98a2c8e38142969ee5aefcf6d4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[5]);
            Id059fc689baea934a9f278b1066a92d6aff850608c0797dd7257693cbfa40102 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[6]);
            Ic6d228f83da7a1c9a71d8fe70d5adbbab8856e5fd3640d805c4076f5f7d53553 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82490f05bd078a3b8dea1d11209ffe17439a638997ccf6e20f67359fb656f08a[7]);
            Ia61e8ceb90369d4ed8ed86b9cdf7d4e89056cf4fca5c7e223bdd7b2c5656ac9d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[0]);
            I30a86fd347fff855a807034e13d6e751b35d4330df8436470af7bb42af947668 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[1]);
            Ic3d44900d87d02e6912d962514abecacc6e1f20fb71c052d58a896c5524e1703 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[2]);
            Ibdb62dc1ed705231a9d0a9e819d824f81e62746fd6d9877557622a8293c7cc3e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[3]);
            I1fd78c97c2a03a51b8d2a3dce2a553514aaeffdc051bfd3820d409da4b8189a0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[4]);
            Ide94701dd8ad54a630c6eadc44221ee5786180f247fcaec8a7787f25c4070968 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[5]);
            I4c5882b979d1f315e20e4a8fc06c794c0217b97de2613e193cb7a213c2119c97 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[6]);
            I5b480e9176a1bb70ebc65f73af78889d266a8efa7414cb97cc5255a5ca5f01ec = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0947044253d3a0486e360a7d81192e3ec15c760d362a91f78fc99bc48f49f2d5[7]);
            I35ddc6b67ba559d53bf4b297c2cfd82bcc814a88095ccdf7d6f22fb59113ae98 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[0]);
            I9fc15e538a85dde7207e48d484f796d96ac712463c802b6995b216e71fb74d93 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[1]);
            I8029c5b828acc50a3a785cab42ada7d51c82647934a9dac7f4a738920f1a332c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[2]);
            I1d5563063ac8386b450a3a36bb3d0a3586cfd6d11471071685e3f7f897d8eff2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[3]);
            I99c4a78ad7af699907cae52326915f18ac1a2a6f9d99b2aa71c34d10fa78fbce = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[4]);
            I1de9fe186e9fdadc6c62a9c6645dccfd3709778f3243d2a4155bdfa20d27a544 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[5]);
            I4b18b20124a63f85e812047188401b685693ae009c87ae337b840a7a3e03f140 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[6]);
            I73c8c2e52e23d992ea9758a361fb9550f0ac7f08bb93b6b26c6fab3b234720a6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[7]);
            I289b4317d3472843dd49dc75a39395f8c39b9fc0c70000205510d08404d824a3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I105491ed20b4b0c24c455617d46df21c8209717604526581da77f2394020a7fc[8]);
            I95b68240d25deb08902e18ba5fc3ed7af68c0a6ae8e629edcf59930ed55c22ce = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[0]);
            Ie6ccfd08b7627ae7cdfd608c7054781099d7df5a0f133672db189134161f76bb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[1]);
            I96ba46d5aa5ea6b2cc6a43df70554584d43f49a6bb171722373d28a2b0f1caa8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[2]);
            I1a54a485e54cb6d528feed952641c7e5350f3d386ceb62ddd2778ad179aef345 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[3]);
            I072f20811fc3b3515b7794a416e5ba39cca6a9579de36442fb39771729dffa8a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[4]);
            I7f1329fd762cf679c07aced91992aea071fe128bc24f06ce88bf49e876578a9c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[5]);
            I26c556de81da143a85c36f6ba98648e110114ab97302046b7aec581a62689a3d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[6]);
            Iedb10f981e08498950a50589d8c2fd5dbff191f233da39d5819ddf2dc5172651 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[7]);
            I2e063205340c315025edf32a4ba91e5f7cd39f37fc5800906a3862780cdf7d9a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5dc456906427bdeb2e39c9a1d79aaee5fb2d61113d155d9d68c6f5b88356fd9d[8]);
            I7bbabd42e7ee42c653f61b4bbd72ed2b076dec2c89baaec2b4589bd55b92fa6a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[0]);
            I90a0e50a5730714abafa98a7ad70e64903062bfe6f8deeb528bdd7008958bd11 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[1]);
            Iff82ae02f527d0eff3c9f8bb9d8fc818cf9bb7e3fac1a127849eea6ba27a62d6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[2]);
            I4df045f8dab91c2eee20a03bcbea586a003659b77d8a6e941bd2b2ead3006d04 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[3]);
            I9e8877d4beab63d4bf103c07e1cd9330daccde2cdd266b2942f56b2a8e8a926c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[4]);
            Iaf763109fb82e88c7ec019f7b9b668f88f84a5d4f760592d2dc9172c75be0aab = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[5]);
            I5059641c5d09a0369f6237643b75899865bff068e9aa8779d0befdbd53a6b754 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[6]);
            Ic24e91afb654a0ee04d27daccc66b42d5e001a5962acd08aa73c3e962e1f2c88 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[7]);
            Ide8930fe855e6fb7dd5b689395a121a16f491421d448454c9c021f62753732c0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie66acb6b881350c655797124edd3d17ca6730eda92c453ff91a5e96df484624f[8]);
            I4909110fd7213171cbddcd3545ba2a0d3a135e723189edadc7c64599fd2f1f53 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[0]);
            Iea55b5544c098ecff239cee665c2642cce17d3b546df6ea3d0c832a118c535bd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[1]);
            Ide09a550a1cc61dd543f2dd7a6e38af908474f7c815ab70318871dece429d0bd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[2]);
            I1edf83d193e0825c58f470cb0d4ccd85e3df4652ab68fe3a701a6ee0e8a0658a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[3]);
            I3f3cf1014fe01e02bb46b2e8a19716cfaecfec0e44fcc344107589dc409044b1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[4]);
            I3724769b2a595469f910cfcf1f002009d9fc27808df7e59ce728af9a923726d5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[5]);
            Ibfb48072643b2cdc460b7a667940129aa243be78b6d57abbd483d5551fa36eba = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[6]);
            I6efd033a5e005d772ae427cab43bfeacb72354d6905822aaf8d484125615d0f5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[7]);
            I44445d003eed631dd6933d4ade176469fe9a4ef0b21b0ee20067b5aae73704d8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id4faf966876a8ffac8e331654199e1260b964ab591261e923f006ab6fe6b6895[8]);
            I8be8cfdcda8c42fc83b767d9cdd6af256d434d307b8e324bd533b5b016383bfc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[0]);
            I31ef992f17daed0e1947c4d26611e7377d8b3049bb8ae2ffb3d56f3db5f85916 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[1]);
            I6483bb2ee2f7c35aa35adc7fcb6cf8cd426e048f4aff95cb9f4f732f97adaabb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[2]);
            If550dcd8751a8725d597ff3b723c6b5cff949b2e3087c71d36782ea291f7bd3e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[3]);
            Ia810fbec78dcd5215c217347900257a8f892a4805dc2365ea79eaff74af7e64b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[4]);
            I5e14fc93aa39853d74e7844854278275828d0f5428f2af96c00c8b0ab141c868 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[5]);
            I8a5d6a4832abe68ab6e9ae33b1b6026805c5db0d186df37fe623a2d9931b2534 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[6]);
            I00c96393d166280a0d866d1999d4306a650507c7bc407202924f6684f61e219e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[7]);
            I2cd11587dc2659cd92fb2c4f894bbd9d252affb93f75c3c691dbb02225b4e887 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[8]);
            I6aaddd1a59b6e96dd8cdd4a57d8fc03132dde1c5b0bd06dd6f0a240c2a04f947 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[9]);
            Ibee0b890887202cb33c8fb07639c7bc536951ce8e661d561d7e7a7355db5f9e1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[10]);
            I0a22f1dc32c83db6603459232e78078eac21f865aabe0b9a03923e63cea874ff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[11]);
            Ib5e2defed9b5fe67a6a551e253cf68006aca5e13092f7e9b53f8186c76a156dc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[12]);
            I102751a9d577151cf6f780ced3299363623ab308737d8483ccbe02118244d2bf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[13]);
            I5c29250eb53f0eefc2332419b6c8e82f97741659657c08af97f8443954a5385f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[14]);
            I4a55baee8cbea583890824bd3ab4c4391b9d44203332575c030077c6e0e9f862 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia72e1164d6bad8b556b6e42d6d779868f93892cdf7029ed11ac48ecb13332092[15]);
            Iaae1f131bd6bb3b2fd8e363e97f6f9e680c7ed035a086cdf2bef5cb7e023c6d5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[0]);
            Ic1711dd767cbb72abed2584c5bc27d5422882cb4299da3914c684696eded290d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[1]);
            I1f749b245e6db4722494bb36009a7da73ca94f408d8a0ca7829b6d5258f78e4d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[2]);
            I4dcd8811ecf9d39f66ab4cf1e07e739c7972e9cf2ef9ff6c0a948336e22dcc90 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[3]);
            I48c76be33e4d7a127ef1f7eb5f4952f81439eced5be914ff90aac6d963267659 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[4]);
            I1a1149d160ca76d7b9db443f5095737e563a7b75de7375f9c148f4f4dbe7e7f0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[5]);
            I67e66b155579d855e0c14e91d2ce1fc6fe1d2f869e4f56b37de5f700d84073fe = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[6]);
            I67a45b7ce414632252362c1556be0e627757c871c136d8570d4300fa316205d3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[7]);
            I51abe903b403df434eba534a1102cabe0a0e976c047fc5cc97a6c8e73263c531 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[8]);
            I0c851ecaa50ea3e1769828a7f51da7a8c3b0c0a11eb9002b108693f09e60667f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[9]);
            I31d4c202b8434aacebdaf5a60c34d7bf3864a5a7c4707efbd1cc3dd82a9ba59e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[10]);
            Ia28734d68fd59a227094e3d5643b87d918753610e867c1d047d8878bd9a46be3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[11]);
            I735ec7a402f471520335d15ee3415e874f56381a2c0cab5c3a5b21f7d6f71474 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[12]);
            Id9db55519cb1208a2555678410c950b6fb31e5fb04a0ae12d6b0a9de4d750b43 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[13]);
            I4e6e6be5d9a7a85cc07a42c3a252e38fad4229a40bd68bec6728e7efa85984be = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[14]);
            Iab63efeaac16bfc91c71a1a0819747c4576111221b2e355300a6e02adddb1aad = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ide72146d090c80f30a5454acb79169de03af6e887270b9828129dba70f0c4186[15]);
            I0e9e95de14abaad3f4dee2c74242d09121b496fc60f22dd3513b90860e7d03ab = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[0]);
            I67874ca15a0723ab01392f527151dd5a60a71a0dd16cbbd572fc50a343c684de = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[1]);
            If434186e818b5a899ad4add63d67ba1dbed823165df4559ee78b39d8c758c727 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[2]);
            I843cc48bafe9c4d2e4647f2909064999da8c2f4d8dcfeaf533fcd12c32c37ce0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[3]);
            Ia6ddd4cda9a70e95a6ff1a9369bb2851b90588337f2cdad6ab43fdd6c6e32fdb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[4]);
            I0cc63aa921326ebb19427e9e06862cc0a42b375a328061bc7f6580bf3f1d3b12 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[5]);
            I0c92cee9eb9e3c8300210834a106174a25005d9a468a481e0f594a960b5995ab = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[6]);
            I3e73f999bb1a0c087c2d4023920d56b1525bcb43f9d1bbc1b49b57d6c9c55127 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[7]);
            Ibfb1cfcf89fe21ebca17ed6bd834fb8567cef4ccfb8f03fd5edaf59000ba0cae = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[8]);
            I4878199f761be0332cf7d653cf1e73cd52f938bf9ca0f32724d499765f313d46 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[9]);
            I9dd21c6b63d36e7dde6f3133ab04263a47559b648e8717de7065e7f140911d3d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[10]);
            I3db60bf522be36d36bdcc35d1d5da9cff2db6e8f89b179726fabca1a7c67b255 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[11]);
            Ic5921b5017385aa779a2016014d381a982c32c64d1643e79631a8ac842d5b584 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[12]);
            I29e9674dcb3b06489c5f9017b95878c6a75503e1dc4e2ba4c9c6a7a7cd74d885 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[13]);
            I6853348c8635a69100a45e6b2b255d6111daca84f2eb28629edd64f8c36f014c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[14]);
            I0bafe9c7cb10e6696f6b6dafb74a2113145f7ef1cb70496d068a61ba1de1bea1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib07f28daa8dda3e4ebfea42be6064012196605fc2769107d157cfbd1992b76d4[15]);
            I929870fcfce11dff715cf2210ad4a4c30db9af500a8d380153f38f0ea2b7c2b3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[0]);
            Id56cc1c8a7f6213208fea3ab1298a107ea854d908609dbe2358ba954989e1784 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[1]);
            If7454cbad692d8d1ed806663944dde3d846b241d1f69736da66374c5e54b8de5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[2]);
            I9d23867d2eb5d9dbcc21e9242aa71e141a2ecad61f5ad2bb69d798b2fdd1873c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[3]);
            Id4f16cdf2e148fb2732fdbe215ff0edd44d29c41dff8c5b307ffcb8305832972 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[4]);
            I32a7df875889c28b6d8f86a42071ad142efd5a66d6328669bcdf1901a225079f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[5]);
            Ideafcce97c26d412480370ab40d8261f37e8bf0ba68bf7d04f4099a517195dfa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[6]);
            Ie3cada5731ce9e6c51353952cfb87527bca19aa77436766bdcc843dd92f1cc60 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[7]);
            Ic56053af1a36bedb5e1670282ac0a93d782faf76d25a25edab3dadb09a302de1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[8]);
            If4f8191d57bfd0311981d36c3836f8da526830c6fe2dae5933650b290075ef17 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[9]);
            Icc14287e817338eea415b9f8dae2527d6e71853a49869ea829d1b51aa7013dab = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[10]);
            I42336bb9a452e51859fbc836c4294468aced58a32a221057096f5119d459edc9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[11]);
            I424c57a79fc220d56d1e499af6318dd2a2f4a4ebab1c83cc7762658b8c34479e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[12]);
            I89b44baf278e7cf024304d7bc6cfa759a735e5da0cf25a96a83e29fa83d12bd8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[13]);
            Idd51d2eb571b7a35413e786a8a9437a5ef34a13b84d269e29c3319a4bb7531de = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[14]);
            I5b2b2323ba78f198e4c86b284772fed82ae708af1da14bfdf215a7b34f811204 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I02e84fe40c4a440d5c7dc0b919caa02f2b4f479a00708766bd3bf4fda9ab5bc9[15]);
            If51ca9faad7b057d5a086daeaf1118808bbaf90b484e38571530cc3bb497dee9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[0]);
            I3c03db46b6474bbd284be2e345d2fae9939f0925a62da2ff9b1e2f3632740b0c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[1]);
            Ibc35679e4c52c119bb0ab5c5a485b11a4bd43ceba90f9998d9704d08ca3285f9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[2]);
            I9244711e562e8ea7e5e0de1921bdbbc5b64363d51d121922f441d8f36e949c69 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[3]);
            Idfb0ecafd00955b66bbc43f1585659b2fd82fa239ab0274450da985354bc4c14 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[4]);
            I6a5f07e66bbd7e05ab9c5adc7bdc99f269386519a6212431d5793e766239e862 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[5]);
            Ib423f5e14b109a601cf9e9d403a7b5c0ca0de8d665d065d8f317760c5705071d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[6]);
            I0dfd7663ac138a56ce3fe38c03c10675da9e417e38f56ea0fa4f9f1902d725b3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[7]);
            Ic3f066b6b8dc09e89e9796c2b739b37e64af709758029ee21800f9fdf02c533d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id5b951c7a2de350a71995dd258eeb274a112c3fc359cc7a93f44ad93a65e91ee[8]);
            I8e6aa1d0b76cee0ce4862aa5d01ee91caa123335ab19a2150e8c4315c7d958c6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[0]);
            Ia261f7672256403997417633102f8c1332ae17195bc38faf0fb85c4e4dd14da7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[1]);
            I4d6d60296569a9b2a811f8064057743f13fdc60379669472d28df97061ccedb0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[2]);
            I81c33c11a5d878aea61749e54e68c024fda21f27f7f4fcf45e5b042e8ca4c3fa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[3]);
            Ia50c90193d9c7ee51018451884df0da92f138710bf95fc32e439b39bea3f3b01 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[4]);
            Ie81fcb1c1ed576d911918860ec73a2b7823bb2d435a0477ef407393052729326 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[5]);
            I2d2817ad47b56d0a7ff72c326eabc6e2ffb1819a2748ffe3a4a42d3794cf2fc2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[6]);
            I80c7df909269b691013f9d178bc3e8c896d4d06ef4cc4b0ac42858888ae8b92a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[7]);
            Ib36374f40465c181d1b8d65f23001a10ffaa250f0fd89077848e6a49a19c56dd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib199706a13db6b68e376532de4c1488dc95bbbe3b30440e60513074b391eb7fb[8]);
            I2a9f642cd74521fb661e381a3f57eaf539ca18ff62ee2130aa94da51cd13d4c0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[0]);
            I2edaebf9e3781f53167708c4854b01219957ff020915c8d2fa7b68e50ede1d66 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[1]);
            I2f928325d150ab718f3b764d3fc4e15d88af5567b4554ef8bbd02f4c3984f544 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[2]);
            Ibf0c6b2fd7ba6e86f7cea34ea8434ec5353399651fae6f00cae29cfd32174563 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[3]);
            I157157e9b85b39f2f22c57c4beae22472512ec83319dd9ac30075b4266761031 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[4]);
            I0162ff342347e70b1361d5f3ea70c6f872d9b95ede7f80a0a18a69c84b5ebc8a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[5]);
            I1f9214a0b2b730fd678664ec457d15dcc243ba1d68ea198ef2792ac2440608ee = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[6]);
            I581a3a40f892233a7bd0dda3bb84e2e46095c27e45d53ed32ef5226f9d25ce43 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[7]);
            I8a3b07f660ad94b304ffecabf47d3378d3ea73b1deccd771fd1982cec9f23e39 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8ea359a607f7bd970935f9025e187a62a31f2a7b021331c359b764985bd543ea[8]);
            Ib1e8234d991235274c74ac026c33d868403b3d03a18a0c674e07dc4f94d614ff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[0]);
            I730afd6404f505477b32f86185baccd692e9e64865f66f048a93e33d1cac8df6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[1]);
            I30b6c3fe760f221d2861a5b6061034f6dee7320a04cbd7de2a3c728427f927fa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[2]);
            Ia7c03e6396e5145d0027d0963c1f8b7068636ee262fe31aa442a5512e0d4e99d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[3]);
            I7fed914efeb5727bba8c1dd0a5cab385a750a2cd9215923b596d1ae914639761 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[4]);
            I0cdb70836bdb3237ff43b23b1676a274cc0dfcffb214799b78ea02c2b59049fd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[5]);
            I5502a12455fae3619e0c2297d5e4a8062415aa3ddd8f0bbf67a73233bb6df733 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[6]);
            I7a52610226b8a85bdc6a0b49cd74cc644d2fad0e8f98ee24c46ccd3664d0af24 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[7]);
            I55d6bfb606269d9d01dc348f732caf9cfdc7042c845744b7a25c0a74d0afefbe = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2814f5d35d7636dbbead87d87d202103a9030e0c355aaadaaa38ac9f1390112[8]);
            I7ba56fb0b187c50e86b74d8dfa7d7b3a1e2bc341cfb56a6343de1e7bb60742ac = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[0]);
            I95d408de4742f651f694ccc8f61d215af1e9b9be2b3860dca46c143e03b3ffec = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[1]);
            I446e1574b1d7bd427fed19be1920c5c29a3276d9ec816ebe1e4465cbb762b1fb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[2]);
            If2f521cf64a5e19b1f744d41d929a37a37689534d0e564224b128866d853b043 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[3]);
            I58d3b6391c1720bf6ac7458ce499fe3b0573e8f7f324db1a796d1126e42e57a6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[4]);
            Ia3690db3bb1809f3df1fcc3a2dd5f807a0ef26c4cf61810b0f9bb590951f8e36 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[5]);
            I0583863d43273e6464e5e65a8714be627f867a0320302382d94ef661b21f73d0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[6]);
            I47d2361b09dd6690b6b0a7827348e9e420d8b97c4b620a4e4928c8cbd84c321b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[7]);
            I6f71faa84bc155810576a85be759d7c06d84dd53b5e2dbc74ab0175e5d64d3fa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[8]);
            I403d7b440509677065b38ca8634080a8edc4c8eae54a9923c50885861866a7d8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[9]);
            I3a8f6218aa06df768133a9b95140db0cdd600a5d1a04a2004479693cecd87571 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[10]);
            I7c843a280d8a673e3c59a22f8bfbd5860c3284b189ffa281759aa44233eee225 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7946354be04c293b27c4734269bca163027de898436544f05d95a634f70d1769[11]);
            I7f31f363b408908ca5cc070f150594db404279b7c5326f5da9abe8f60138bd51 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[0]);
            Iff8bdf9ea44924628e777925357dcbe728f0ef4be0a3574965c811485fb57689 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[1]);
            I0d58818dc0f3ed67f1e3a10ddc7cd0592bfcb8cb3db1c329edea24dfb0ffde5d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[2]);
            I16863fd89fef9bef09bbfec8d23ba6d42f4de7902a5928e9b43546b4078fbb0c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[3]);
            I1d5510ca99815d74f26804206bac7f1e7eec3727fa89d91b014becb49a815abc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[4]);
            I241e6ca6efe96759bbb20d710c448c9c322aa3345fcdbedf625e297070af52e4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[5]);
            If8ea1abf5aef298950b84058c5e76029f717309fa685556f09c32b72959f648a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[6]);
            I4eb03f5790e18ea72980b8c37b602469d6dba5f850ca3721f49279b4e14cb7c1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[7]);
            If4c7abf17850a5fcd64bb4ebaef1dc806938542a3bb2b9eee643fdfcfeec23b8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[8]);
            If15171a1904299c55ffc5b4c9059900188c1c87caca3f4807c4498abe038becb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[9]);
            Icf3a16773d04781aa96eb511825cc59c609fc887b464a86c7839c57ddbba37db = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[10]);
            I5eef24c8de2049e0e8bdd49346b6be22708a135d56c096907e50ecfbf3affdea = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e0407fef05495bbacc60a763aa8e7bedaaa8ed4285a441a84ddecc88515344[11]);
            If0d87a6c6a4dd34bcb5411a845e6e7bc7fbeb0e6a34933f64283c880ca5d3d8e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[0]);
            If8c51307ae2c537425caa18b7c3dbbf0530e94ada2a2a600262f57f93bf60d24 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[1]);
            Ifdcd4016757d0cef222265289850476e0e2a6547732f999ca0cd8449f7134bbd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[2]);
            I27737e1ab6f67dba3964412127cf6c91c7a58f6ba77e5b6a9808e2775069ad4f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[3]);
            I72e85032ae85773b79f3a3dab895c9667cd32c6aeb44c000096ddcbc0f7be0d5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[4]);
            Ic7abe3b0fe121e025ad7f7802b7800f4097111a1108ad088e869e81e5374c42c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[5]);
            Iccb7ca5c2ab8a9a4e3776ef42997d1d645c5542c25ed35b161702ce450f90fd7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[6]);
            Icd7ce463860bc6f62da8d62b71970658ed2c5d5872a56b8429d9223197ef0ad5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[7]);
            I8952c026089661f4ddd0720f6ab16e46334fc934e6775e7163aad8cf5dec6b68 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[8]);
            I9efd4f4bd4d8dfa270cb1c5a2e3f5c6cbfc3c5b672540ca268e0765170e6c748 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[9]);
            I4408d142165f7f5bcee86e820e4ce79b4ecfe2134d8e50809080e0c27e4e2df9 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[10]);
            I29141cb56b9f52d74c42d689b180cfcfe7daf23ce573c1f4eaf21525370e5376 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5a1850c40c5d046f87839d8688d1336475d1c6f15829bb9ba5cc592b1df0bd02[11]);
            I567366a85ce4a20ac4125a297426463bc2f2c71511a97bfe2f4a01f6e8da6403 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[0]);
            Ia71d81a2779b6eb5f39fad80ee4e7bbcf394b97657cb094aec163180224939e3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[1]);
            I9beeb3f92470748db1e059cd6c5a929d1eee2a3ecd0ac097032c74f4134a22be = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[2]);
            I387ea75c114fd752ced502cc147dc9ad385dbf69607c04edf81ab74b6867f2bb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[3]);
            I8d10cf5dcbbd1a765ece13156db0ad4651b41cc5ee286720226649a707accd16 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[4]);
            I55d5daa0c4cb89aac08ecbaaaec1d6afa2379b277051281d3c15abaa6af05edc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[5]);
            I5460bdaa1d2a7c1cb2e75baa2c211593afac76ce5160a620b385393217b4185a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[6]);
            Iba39b0599ed448a7fdb07f6042ef972612b54c7251b256373b30788f64f616e6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[7]);
            I58db55229ca30218227b598184e85d57a0e3a8b61308f8114cd709232573e566 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[8]);
            I94ba926e07e8b3cbc5429ff6bf73020e95dda7b7c0059dc10ef646b2980bd80a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[9]);
            Ia6058d7a3749f21a827ae6a0f4e792d6cd62ab37d668d607861bdf3985489d97 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[10]);
            I405b2f517ad52ec3c94eb9d1d695f6fb9700fbd32fb49fca23588911b5dd0ef5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I501041d56f5195310a81b93f732abcba9732d90d5b494e651ee823e95f146c53[11]);
            I0217d8dc004467c4c431dbe27dc564c042c33d06a5be72a29ceab927708c4de5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9aea0703810e5cd52352d3b0ede17aa0ccb943f1e0507585e4cccd0d0c427e98[0]);
            I14102f52e9c6fa58677dbf1260a5049a6c2807b245f123cecfc3f1a413badded = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I42c6c1d7cfb81335f01807b1d1c6b77c109482d338e81eda1ed174f739a6bf1b[0]);
            Id71b753d1cf473f4f4bb7718f412471692e08afc0ae9d25e617c2360df79ceda = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I839de42c6f3369ef5c6200c12baee8c9e698b3108fd6dcd58a71351d9bedae54[0]);
            I443558f78c6ebb16bcd49ca586ea62d2ba12ed3bade0e54ae9bb60f83d2598de = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0a1e88a592eeec68c060dd84ca2d75809b8fd80dd97a01a8d12cd9869bf94532[0]);
            If5c2310896ae5dfd3f83de1affe79fad0f0b6b2b673efbceb7d296b33a6900e7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9114e17d37b4346674c23a6ef3a2aee35426292fbf73d7f30c895090bb749034[0]);
            I7d078740e07b48774c64f6dfd7bb0f56821dd685e014f0b9d4e3b7da45383e34 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ife5225eb20e50e3cc959d9080f6faa318b4977bc9d04a67414a6cdf16c98e295[0]);
            Ib3562b77830a64f31728e11cc54a6d19b55344891eb82355e3fb4491086e8808 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I28dfde2c443cd84194231fc87b8a1c6382ff3c2ff9b6d43e31e3a7116be41169[0]);
            If7d42431922752de30d5506e1d501f65453a4754d7cab03976695cdee9c0c9a4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I55da00c15261d3abb33c69ecc3f2090fb2bb3c29a3653fd999f6232982cf31ac[0]);
            I269a90aa42086a30a9b03141bf37e3abea46a1f1c06710baf2d052a5bb404248 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I05ca033870ef7adc8ce911a962bbd120591a1fe3b3044782b7e569e2b94ac629[0]);
            Id88de8b0cefd527c486f8239ff6f61d6ff86085e420d2be56ce58f4d82d78a7a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4ef4ed6e15f48f289815b7e00b2454a26e076b8dc9b8903e118507c9688e905d[0]);
            I107db18dddc718b9fe7354d0f352f72df94ad4653ab0712d5765a495ec29242d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I25e57b538f9a08a355a5ff8d26d94f81bbf2ebd0039881e74aec76ffb1dd48aa[0]);
            I642c0e5f0768f835a6ca3ee6f65875346121b502770acb1ce833e9aed46d4ddc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I070ee6bd21603d58d3243ac556db2ca3c0476c64fde6d32aff54e0577b0472f0[0]);
            Ib699efc076bd227e0138482c43c5fc8cf0d0d87078e063262fc4b537f554697f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id2ede5f3d3ce0652bc9ceeadf1de91fb99234718893eea8cc1779cf900284e88[0]);
            I8e0d77d4d38cb3b1e5ece19e010043e9a4f0802819f3e70f0ecc9440f65eff4b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie251294e2cb883a913e91485cecfa90bbd107955ceb6d60d4a9b1808aaadb2d4[0]);
            I3eaa094e28f19bdbec184b0ba0f3792f90e67c77bd8dff9af6042c5002735505 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I983e8c64c323025590663edf53b0666d93d838f15879b5e3df245a8e9ac6fb80[0]);
            I62b9322a1d5ff38480981e00d8469983588d084289f2f927f3339250b5c35985 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46e5ca785f6f4304dbc4fbbf3816d83106047f0eceea77717a1ad5c41a9ca441[0]);
            I2af0f38cbf134ae07c76f06d4aafee537bcdfe91b1c4aff1ae27898e18da5113 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ibefeb67be2754ad6b9a6cda09c66529a7ca51536f5c6ca6b05e6ac1de34ae514[0]);
            Iec6be5ba578c849ae0e4fee9c059ff88c36cfa7c14cfe218cad7f7f1d6744024 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0dd45b65c82498edff9ac44b5b07ed30818dc1ea2af48e5c1394466865f36adf[0]);
            Id18c335cef6d5d988e55f6fda5a09a24ee80f4d4755f797a11ee94141b69b97d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ica92be8c7303e09b9f549ec558e655816c1d23a39b8d5324060f64a391984c1b[0]);
            Ie85ad3f88a177d67b69eb3a03e4a9d92f7431af9de9ccd06f2caa01f9d144f33 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I726b6a7ed2ab76b049762263a08d5121a597f30ce25a6880b51d6b01aff801d7[0]);
            I53e788aafc97015db67a8363c91d81d369d80c4d24542fa45faf7833fa4189c1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I89362accf0644c192f06b113020d2071f1389e8ddd8d4fee492205db15b25b66[0]);
            I8f74cd611f5df70ef183e9d4a86b5ac23349be8cb99cd470c596fcaa6ec95248 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4473c0cfd2d569bc671ba814a524058946271eb49a04fc384e9373185e1f4a6b[0]);
            Ief3910aa326e0d9782566c81ab1cbd09faf46d3552f78d7ef5fc9de1d9c245d6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2ba73f603d9cb767572f2b2f2a9732e2ebc066392aa85888df87da4dd8b84113[0]);
            Idddd98e139a087c7aef3922ea2542dd364c9d30f70665754f751ed88dfbd3701 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I82f10eef14d4ad82b1f7f8c5d056c398386a6cf790095113a615a8bb6cfba233[0]);
            I474f7c67e6159d041be6d6f4f96fe58f9b7086757936ebbc86340bcd9cd9962c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2fd5dd69a5f551c26d9970d09ab0e26ac5183a0022af58e2bec1dd1efefb139c[0]);
            I2a1c16f7d4c3261619c325f4b5cfe98993d5957a2ff466bae11c9cec6006cac6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2fd258374a5bda5c58c1fdc6e305789a598fbe70657d6dc18e8878b6c2b0441a[0]);
            I881a2d7025d422202455bdff165dd982c2f4953b361f29688e75ccdf9e04d476 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I76942d3b012aef2097112a1c1adfa2bf986414df19a633b87d2f3c2a61d27351[0]);
            I8245c1ad016aa3d7290e1097eb966b09c8a38fa5bf62bcb7ef179f448104f47d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ida428d199205588ecd8cc963ceb39e24bf6f2d004b675f3cb883960e0f089842[0]);
            I10206e80304f6e623a256b6042ceca13c691a34ef5b6d67667ab4bb11f0b0087 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I91f0247d07693c53d716345c810ffa0ee8d3f4b793ca8831763f5465db649c89[0]);
            I50f15058dc2e50a994089de4a0487158352c882d4639449d9db322a05ddcba3f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I754c4c2dda64bb938ac60db8cd469c6f3ee0831a3a6b6b98e902c1b72663ff28[0]);
            I0604d25b233f4206fb580d729452e9694d4b795553a4a788f993c992bc433b0b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I567c2801d5598a057d5773ea5045f594de038bab88d554ad2c713cf56ef632b4[0]);
            I5b2860f88d7cbdbc92264ca1bd0f97c610e7b1cf340e2b65832553a1762fc865 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic9f57a4a1184139b219a3a5e3c554705469b79d3ab175ddc74512ccbfd5898b0[0]);
            I62f27f0dc53be101d8fc7f026a673fd33a5397534153859f45c113e6820e9c26 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2dc38e534505cf47f391eb9f4b090e16136d12619b4fe91cc8029bb5a050689d[0]);
            I92cfa50424ddf1ada795366ac6c7b31cbb1b1330486911824b881a1fda443c25 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib83aabc196c7633dfb4a9bcb4b8d06959130620de297f9dff77b1454a8f2f96d[0]);
            I1d996fec699e93fc4ce63060990c6347d998a81f0b3aefd88339d5d620fd152d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia23743e423f143b75923bc7b1a4363323d46ace080c8ee9d15ff687afd4bef65[0]);
            I33546fedf41dca9168afd7d6916823e8c24aa3c4a855b93820215c68c807a56e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id49eabe82a09acf1b3a3aa3be9bfbc0ff958b96b44ada842e892c587fbddb8fc[0]);
            I8617f958a4de5cf233240840c770360befaafe599fbec1e351b24baf301ecdbb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I93584fe5ab7128b24b2372bfeea00f7a2bf09d50b1fb535d01cc141c6d6fc377[0]);
            Id824ed4e68ef3624b9a4d6c5924b08a7b727df62fc9135c973c5f79768c627fb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I44142c70d3ba4660f5b85d895710afc623ed3470ba85eab3dee5e49a59e1b124[0]);
            I3d71ea5bb4c4be8ea80abe59367519a071132c913eaa5c6538baa8c3faf243d4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id8b538e6a6c4a147c7000388923f1d89a193f8ec53ef214556e005218d2c240e[0]);
            I6adbf5489cbaa65213fe0804e7494a2b8be9db9132a6ab7058764a1a53480999 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I658f9399a929745b4ba467a1e019fdbe214acd543dd4f5f51a95292420281401[0]);
            Ib4e392b7b8f87358dd5cdefe7c272531bc6bb1f27bf1411c1a2f4331809a83c5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id1ba70174cf019078c719d1d50a82a61fbfdeea2a13e21a1247e567b9266365f[0]);
            I6b528ad76bac25170636a86ebaf7efd14ee7159ea2c83500021e39e968786428 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I797dfd66b521bd680024b6e46455d624aa58b4271f5e6ca19fc7abf520f26222[0]);
            I294be7c0765f0d4209d4442136d706edb2080883d5c78a3c71d66b5946116bef = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I74f49d84817f2467b8ccdf03acbd7372c58f1a4fddcce45cb882431b2be20b39[0]);
            Id834a34ad825df7c595e3754b5a5638badf560cfb68ec8de2903e73e88b1a113 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib756dd9d8d9a5233fcd368ffa91f5d7d9c8825b01bc26140e5a717d3ce263e64[0]);
            I09e3897931014e7bd9540023eb8fe1097e36eb5c51db24357b492a132c3a8805 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I1bb2be29dd44258b24a36ad9b1625ead1cf965856f1d9695c62ae80de142169d[0]);
            I674ac3fcd5872491a3c412a02e367a9c29e4dac14a8ffe8b6382c60a29fde8aa = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icbff209e6c8353c58f46c0688f06da0cdf71a95defd8937f2d52d63d387d74b5[0]);
            I9ac796f1901c19aeab344ea2c785af3ce41bd23dffe88b1b5216f8f8c0b16e40 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia628bc749f04b3d12509effbd4e0bc5ac0fadf48a2cd5663e4c2094593870a42[0]);
            I0d186e0127f200b704a4585b2fc43ff1a9ab19833a90ac881abde94b2da89376 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5ac2c7b61022af9bd2550f824b8e129ca1c336b1ff900b0af785d86e33cf3358[0]);
            Iae8191d31be3785db5d8e5d328fb2d96b0b5d5ecc7f9d14f0bdd3f61a9bb6781 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie511320217185f90f1e4a23ab51ae9686801b09657c714a5bdd9c4e26f070bff[0]);
            I4694c593512d9d84542af4ca5b0f3022f9b1433d7d6435ffd4b1e53093bf4a58 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I032b833c683eaf0c1c4c60ad831278ab0ed11ed856361be3be59dae656141fb0[0]);
            I78c5059e528b7671e27f847d6042b3fa707258c664749d857004679c6ff96a73 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib41d86b318a3004b648c9a1b0ad00bbb144511fd63b1c7648cf3ccfb996686d3[0]);
            Ic83ed3610853814d7c9d6932b644f9c924fec7d67e303160a3c5b99c625634c0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icc4bebb1db4145f9cce0fd4c250f7501f300b6cde1f31327d80b844adeeca1c7[0]);
            Ie33f8884c8fca47e2055b28f4398f3207f7ea20f8d0858d2a0699ef2da5a8f03 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idead9dbad4283dce602c05f81e98610ab7f65f9911342174ceff7c95dfa9ddb0[0]);
            Id140833a04f0b4b903ad4e99046b17f76d4c405703fba227d36342b6f1fdbd08 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If7060467d2fac9aee8d69c5ebdc24d515a657bedea3da55d13ed6ed4e3c8e79b[0]);
            I90d7a3c4ac0a18444eceec2569cae3d5dcb3d33d2e46c329068b0d35ad063971 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6aefe769159bdc69fee8e09e46357993c13dd8ec9f059cd51d43944ecd7ce3ff[0]);
            I5c7c7df860c87ada06c17210746ef84d27aabaa26e9cad20397822629716d4a6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icac3a5cc88034cf8211c158a1bee2a04c228afd4eace1b50c7460ad5331ae02d[0]);
            Ieef9e0d39f2e213f365af4a6a34d0d2c7d50155e8052e9b1944473641922e9eb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ifa5d23491b028cbdcfd79fdea2e0784f068c1fd381dda7ebfb5d457800e510cd[0]);
            I4771e59053fbd3e261c49e0be7e742e7cf9c5bdad030b67f1b955e13e9bcf083 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic27b23bf87ceb2ec2d6460321286d798980f966c89d0f8ea42a79a0549b2128e[0]);
            Ic8c13812ba09457021ec6f39406b1106dc025551c62da4259930c361f19c3a2d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I01500dbf2528609729acf26a24c11bab0adf8cdbc0633527f21644816cfa0dc0[0]);
            Ic7aae8edebf83f3971440fd0e86e7700ac4cc0c087c9996d55cfecea8c489fa5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6db96717b6fe00f1f87347adf69ce2d4b4464faa472ca989bb272b36454e868b[0]);
            I091bf548253a3b22f92aca6479b70ccb74a5f9eda8bd80e6bc1e059021f04b9f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia8cd57b3b123e08e2bc00f82da941eb4431cc816928254135dd13ef52eb9c03a[0]);
            I5c1c30033bd61b271c765ba00b033a58c6389d4bd353ce68d1b193bc7138baf4 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4fa8db615d84b02196afb2ad926769bcbfffb7c81170387b4d460c7403f0dfab[0]);
            Ia4370635785f2b904fb6ab3b8cdb86fba5445230a9d3d02cd908e04d92726f3c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie81813a1836449254acfcf7674552545d2cbc852ee2bd2f37378345ccdfc61b4[0]);
            Ie73ab4d16ef614a27522cdfd47f670a38ab58f89bc10c74975cf0b30400e198f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id9fde3ad430d66c92a5aa6797b76ce147e39e4245ea761e36d81214e7a02b4d8[0]);
            I76b8cfe5d3985f3c0f249680ed81aa3b21cd7af725925846e8875ef9e98a550e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8f2cae5483691fdf6ea64a4ccb2372967aa676835ffd4f562269bac888840d17[0]);
            I58919d58783467b7ad0108f86d6260f3c551692d00e6639260a68a7a512d8689 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icd8572ba29de1a399bc077f53730492f4e89deb95b9136608da0d029ba60ddd1[0]);
            I0d276f9604ec2b8621a86706ad1772058a29e94902e8eece60e3d07948e24cee = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6eab6bb656dc82d656eea6da9dea574b230f56c6ab898a7f80973183896d8347[0]);
            I5463c05b1b55c142012470d627accadd8e34924e77ef6d139b3fbe1db1cb91e8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Id802e388c3b33f7d0a0960e0e51da02e7128da423d518a916f761a16b73c17d7[0]);
            Ifca2987d8c7f1ca30013ddfcdb82a888ebbd7bc3dc421f7e3d6806f5f3a9aa2d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I47507e717446a9ca85cec7e5fa382cfe435affddcbf5b25d4e74f23a143b02b0[0]);
            I5ff269ab544d2b74059a73d0ffe0492473b214d392d8c2ee760847e6c07a361a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0d76ba051f3db8c1efd9a8f0bd0ca77cb28c7dfd68cf4c290ab00edfedb15237[0]);
            I26a6366fb57427f6a0d87d4cff8a293a0752887e71b829e747c27980a1a3dbbf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I39dc59000bb2e3fcdebec08ddd22a460fad0c09e8b68adc7e72a6e4c3025da49[0]);
            Ieb5560e3a4f6a9c4543d941ac57bd3805afa7fa17624e5739e8e639e8d0d0c5f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6db1df05e1ea3d8011bbd6e08c9d50d91e672a20aa2448167343b839e8f6f888[0]);
            Id1b9b5118024dfae0e058f5418c9e988e0a5a598ef7553947de6f92cd7399201 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I0d11d2b76d26d33ebe0c7577f5d7bc68ab8f4840deb765b17f4f7fde0a4b2fae[0]);
            I50e1a6fdaffcdf8fa99074f4480dcc21971ba8f5747b24a33232f9152b07af1f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ifbbf33f600185eab85dd2c0dc5ab2f5e0e2cce52373cc2acf5e466a2e27ded58[0]);
            Ieb31a59d63544ea160d3934f0e38e6333f8571e77352bdbfd338d68c437f02b5 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia38b628fe0740039fd44aa0a75c751e1a9e176bfc305a978377c1fc9525c00e4[0]);
            I81e45b654bee6c74edb5e034c89bed7151c60a69b554a35710d1b173fe45ea22 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Iaeb5b860946e41cde629a762ab6e6ea4a0f177083c9ac84d90ca99fcb90e7c9a[0]);
            I5144a2cef7d82b7a91f9d83ff8fdea356bb01db215bc167f0c498d55d1faa622 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ibc0b2c21012904530a727f0c5643b5187d7bb8706a308bdd0de67a80147db974[0]);
            I67484837f2e585fbb85de404cad8f08ba58bd1faa81b9931f88473d7f4a9a06e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I008d6180d4774d2472158544239ee654e73570389873b54b695946cb78ddb7e8[0]);
            I4404bf7e923ee1bc0230835c00684d298572238aa8b9602dc48e177464224a53 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idaea720265ed96d87e8852c36eebd63e2be5b9768c7803f13fe85e7532b75ea2[0]);
            Ied796eff44d61681c5d5de05933e785d387a97b2430fee26d96b0b24a1a54c12 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia7bf8296bff6d2322977b0a31ba519bca04a1d6c6f6c0cb5a47e3408bdfac573[0]);
            Icd8838ebb43dad19fa96e741b32851dbaf5c469e0591a1231898a7aeb6ecc788 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2a69131c92e4454ec846c7528679731db69a2aa63420f0f22289d5c0be743be9[0]);
            Ic6d60bc06b0eb51b5ff4b8cc0d0ccf55fd8e5c53aab23b3994ca8d094920d619 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia5fc094477d9d66d7fab491b73a00f50abec21827f63372fc1b7e0bd31ccf375[0]);
            Ia0feb2870e46760bd3c58e5af56a40a73fcc6c9611766c77c4784f88c35f440e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I41d88c1cdef0448f878686d88600bd254e722761979a244cb1d00724fc1d35d8[0]);
            I60b4f2cd3f513ded6891a6506d0ec74357660440c94e62f4f7e2f886c1233204 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I85e825a905ae7dd292f400406048736ce90fa7d47b6dc5507254283662fc7564[0]);
            I90b9d06240e2a49693ac4ebe37203439a157a38d068e630c45341d7d677b816a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I80cf17357df8073b050d80de366bbb919c5f6c8983ca87f6606a84df1b92c549[0]);
            Icc84144f0fef09379e456de5410487e7882d373874a686f1b61db92511a91e2a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I68a074e808119d0f33d54d3863c907dd5d761b3f6b144b9283e67f956d5932ef[0]);
            Ib5ba52b9ecafcedb064e66c38273f7833d0b6d0239a7fff9ef3a0e30d0f77dc8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4aab61ec97ec8dfc8da6d2ab5898bcdfdaebb0f024fea498a6ecbf0bd15fd1c5[0]);
            I38a6e64d23e0dc1a449445bf10e786777e978aeab68b3a99dc5335b93c67da45 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I26395ccf79a44d582b559acac5845eae4a01464019f7739b7d52d8c8a4c11154[0]);
            I83b2a186b150fb7290623bd1cbab9d044e9b5c760ed36ae218fb775354e46fd2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie9c493e499f4b2aa598c54d5a5afdf39447612225daf7f9f5b3c2a23b5ee0ff0[0]);
            I507512179a289ecb7d9ddf5e853bb42798df8129655c06e568e0a4a1d880ef71 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4368873c6f3e3d6ba5e7e83747fb90120e80de634655a9d2a97bbee88a9d8501[0]);
            I6182a01d42a30ec5e8883e7d4f5d8f1d657f78052fa4c8ca2c160aecffda456c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I082b315a51a6a180909ea4f576a9a3c8b0550e64aa222610c2e6906ca78aebad[0]);
            Id645d98c8a2ba63ba9060280b1810d0ab7120f007f3f174e1a501a1f487190a0 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I23872b1af6db7e455f25a7ddcc050167bb10de0afd16973c0a90804349210372[0]);
            I6822880688515ff8108fe78fadc5d22b953ce5face9928836f824aad9355a713 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9796589e7a8535d47d56f792d80838aa402e3c235035b517765096d2a6843215[0]);
            I694ec7b5bec025b308c4cb56eefedc2be0842202dfb047b5a94dc749c757bdde = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46d39260d96216c08b7940ea3bfe542bdbd0966f5e798321bc90a2a00f64360f[0]);
            I99a4bc7f129030d12eeef0507cf52503af3df70717d1ba9c38b5dd3a5ffcb616 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I1033817563ce88e3b26188a88303cc6703f47afdaae4d5457fab8b73bade5274[0]);
            I668aff5da6360f719a2467c5189f3e53e8eeb310f4c4e26f55f8c39e9dcc4be7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I343bc73eaaf00a82b2674c8cdfbbc5c6ea52d10fbb9e9453cf4fcf2421b97e47[0]);
            I4583579034ed3bcee2ef0ea2b32a4adf0467f78a2770a84da9948e8d366c1f4f = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I1af6f4d00567aa1e302e7d8830d761e7a9a616f5e4e958b264701c476216de4f[0]);
            I86729a880fe730068d538da490087a1ab6789327f964722c9c14bd9b1c2af35b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I1682f44d820722e2566b0d6c02fbf3dc72547221d519ed071e7c7d77728ba21e[0]);
            I0f8046b4f96acee2bfb4719bbff91b4b1b81c78ac36ec6e95008a3d9cb5ea6ff = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If0095cd5e911c91331d2ef6ab3866101080b3cabe8d1ba9104b6b5ae5d18c713[0]);
            If08c85e70828c39162bc16d65747d3d3d0a6176e8db106b262bbadd651f745b7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If7f60dea1e83c3f86ff8ce3adda8214324b2064d06d69ca68477288522ad9de0[0]);
            Ia0ee127b17b441cc11d664edf15d370368494e31b52c4865c97a065ef8bc43b8 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I3b1abc53d350b3b39e60c3a5725e5a21632e7f0275988b98c1fdaeed5342f9c0[0]);
            I8c494bcba3ff73ff29d9d388708fa34caa73b883730349aef6c2648a2f5a1409 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7943272afdae80761f8b673788c92e4461bf3de3229f7addec1e54743b11beca[0]);
            I7ea6f607967e7d251d71b4c4b3dd545a4a9ae8298c3ee2356bbc16ebef06cb2e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I8417f8f367de885ebb86571786bd964d4a81d6712a88c3a8071c08d13cc7cf58[0]);
            I215148c89dc37a59b3eaf2f38679554281379dc6c8e57718e1c22c091f4d76cf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I653822ee3643c81b817be0d9c3f682d0c806ae17dedb0cae5b1aa0ca914e6857[0]);
            Ief3b5e8fee2d099a90990de9303f34d600235d989d25a30b5a7e2654c18b5c3c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ieb917f5db48f3d352eb252f6ce309bd972cab47f09ba1c140f66192b260f3925[0]);
            Ia2233f4704a9724ec75efe5e31af6807f8f1529f641ec05d053d6a12308f485b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I313a01d9fe403e838310c49dc37a50b738025400e99faefbd9b8cbd426edcfaa[0]);
            I6754b9c9cc470509e67ba88c2669e1f70666489af9ca14de9fd4e4328d18e245 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I1b81a8a827bd2222ea6820d80d13e537868e0157970625d628f0c062733ec3d4[0]);
            I133d5432ba2f64f1ad612b2505fb95ce91962b6ac761dcd0e92f75d1b663d7b6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5615438871373f7ad838fb5e8c24b9517fb94ecf6627c803e66a78f778fe9c42[0]);
            Ifb664074b1a8bb954cb940a11ae4e7de1278edf3614b861ccd83dfaef95319c2 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I07f9ecb15d2696b2cacc35c935b497b2f8cedc55e2a661fa57f2d0783e6a1001[0]);
            I76ca3c17438c05fc53f6f7075ff7404c0838f62472ffebd41a61afb1f3ea5dbe = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7fbeac90b85dfc78e20281021fc1d7cc90f9deacb2091ab55ed07f51fbdbcc11[0]);
            I27ed900fc3d84c4ab4570c3bb88b5e9a7077389e5fa169cc4e1d606f09c9c755 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I46dfb75396740f84b7758552420a7ba8693bb1ca5259a67530c588585de1c337[0]);
            I3ef4c55a4a3281a468daa3233ccdbe660c46a930220b5c9bd3caf6041008bdad = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I60e36bd866a477c35110e2688e7fbb13b0303d210e014c9e151b313d130101a8[0]);
            I9d323aa17bffd7ea7a66ef99d4d004ce664a0e7e5388ed24a4d45c69a4d9b396 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ibb36dcaba8439f48b18ad2dc8399df26b940f7cd815996635da092d41ee5b106[0]);
            I8e6a3df905c8c5778e1fd6e75b091c545389651762d9cb3e0d21b20d8dcee6ae = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I387a4fa48a52a029d2bb0c8e5163f15c4cd55d570db8d89e5f73d7bd6e21ae5b[0]);
            Ic935d033e29fa4baba415347d379eeb1645c65388d3c7c9858ae48f5a098e2bd = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie2ad7096c10eafa6e451ff7793b2dda562b6623b1eaeed56bbad4019662851ac[0]);
            I1f212ee134daea9d568f52fcdce6452048326c2dc243c60d25ee71b95ffea50d = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9de97cb2569312c40a541c0038e02c03024581050590e5677dcde888f4c6c3ac[0]);
            I3a25f0d4a6f0fa33f493d9aec6fc7a318a826b3885a3cccf04e9b1a85bec345e = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7a55e4af3d00a3684ba08ac52c3dc7dd0188efbb684b859ecf017f783fce247a[0]);
            Ifbee83b3613941d8ba27021c2fd37d0990a8af8fa3e0399f0f1f8a92ae18d273 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib1644713e1c2c63d093c8af3a2be146dabd70cfe25a1a6ac062174576477b113[0]);
            Ia1c056993094512262fa3f3d38a2a46cd43eb08114e1af8c48ce2f6705d7297b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie907506d9949011db3e41c72b9581fb832dfb29f82249768fd9893a3de358b35[0]);
            I61e29bdef580f4f1057d7b4ffb5bbf37c67d3b8107d7979c2fce643282c7d861 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I678204e14a0213dfa7135814f07e5f6c4d12452a503ed555ca2c20c10f047d5d[0]);
            Ib07a3587e3bfa70ff5dcb296b8595c5d15cb8a94efb13c3e5cc92cd3be3605ac = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ice68b876a3b3943637914d8d12aec7fd37cb867f7a7c20be11a66dd85803827d[0]);
            I8c443a2690956ee9d0171ca05534d698f75563cd74ec9f4de33c7e8dabe8105a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I35e112474e97e65f8e8aa9a4dcce274c7ffda9cdef901ba31801b4daa68888fe[0]);
            I5dcbde9462714577263040534f0560b0c126ba001e959add92d0529cbc94bd9b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I84992c3714fef30f928dc3330821045f20e176826278d42a9606f2dfadfcb9c8[0]);
            I3872eb448ad521cf99b3a9d07ecde078320dcaaac45bd387137deaf5dec956b3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I011fbcda61a4f528c38920d0077565c4592c5f6d1a2f5a1a7dcb6a4a734e0c83[0]);
            I144443166f296f7fdfd616492bb4b1fe44e0353fa6b0fc822b3aec0c1ea0c894 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6d2154a30adb0faf296cf58ca9229eb1a298767fccc4a1214092a2b977f7442f[0]);
            I5445f1e35f9039ef623a77ce395c2a888153749fe8226e9b844b271c1c69d760 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie500f9b1405b49a263908c145ee4a337f2ba4cd2d4d784a2acb77068d09d1662[0]);
            I5d9ebd6a6829c49b0e41f700d29bf8acf06a5dd87192846e5ca204ea8bf563eb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I26997f7f737ba99dcbde55d67661cf9e4efecf397b1ab3ec59e0cc5d8654a75c[0]);
            I7e26d67803410d5079a43dbf6053aee09ff9b0242133282679c3beffd05aae02 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(If6181a32c0ba3cb93e47ed1f1279bd4e739882c2905d6d64d0149f26d052f0d0[0]);
            I685960b47e49f3ff64eca0e1f26387605e48d325d533550beca6bd6d0f3abbd3 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Idb4bd19284288df2a5b701cedcd57347e4f7c37947ec1588daedf3c9ede0a12e[0]);
            Icf75218ad23cd1505d2d69d09c0305642a8be48b8a3b7aca4aa4d01a564ddebf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I4be880e4f25fc41932b9ab9295794ffa2f334ee5338ef0d59894d18918d3e0be[0]);
            Ic9adc8e66938cafc1f6974ab9e2fd71a29bcd6520e6fca93ce7bab4815494ed6 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2dacf26260c042fa148fa6c4e97bf878ad2e89e221acc0616141e1841b0c320f[0]);
            I4f8e5bee14ab1e584593fc15140a36cf071f2949f1bc86fc3fb7dbfdeea7343c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6cc3662b07a43d62f870bc24d55a9e5675a0e50d923f3b293d7004c2c62ad31b[0]);
            Idbadcb95f603dca2fe62a931973c10429cefef4d6cad0b8e46cf34b2f7c7907b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I670beb5586ec69af20e65eeaa49be81826908f01db21d27643e2561621962b87[0]);
            I9f94e32610a6e83f5ca5d8eb0ad81277c7226ae8ffa7f1e734959a614bf1edd1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I88ba583883fb596ad6cc6716008143d6b643816e8e694ea5f32ba95f3cfffe48[0]);
            Ie023df7145a8643ec413fd62bad9e4dafc719f7c882ae969eaccbce255ca7748 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia8545410ad46518007f6812cf6132f4f4482933818a0fe103dae14b1530518d7[0]);
            I3a210f2cb408bb61efba033b0ea8f1cda9a3341500248e1443840c24dfe04cea = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7018895fda9af57bf39b18e9edc144f8854067ef25800ef8eabe76015fc207b5[0]);
            Ifd9d392bdf654a9146eebb9a670b75f4d74807786708350ceef7c79d54805ccc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ib57f995d569a522f5562976385f777cd6cc39ed15491d0ad8f88cc0e908c326a[0]);
            I3cf51d0ae95d4e3f7d0809785f84c5d25153742e5dd0d370235828d4f9c0d1cf = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I35636bd5c56cd95d41880b5c936108a3ab7c1517a8e09f76731b2154d39c87f8[0]);
            I4fc7c4344699ed94536cb79d86f697e9da22498a2938b10360763aa9bad9da33 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I84280195e0f72492aadcce8eda907d5de2e05dc16b9c5ba1fc2f345192ade355[0]);
            If7b4cbde972a67fae839c5bc9ddfd64dc244041f6dd60f95c5329105ae08e460 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6532aae67414dd9e03b874fd4b6a321437892a7d89bab17ec2d5a684aa9ad55d[0]);
            Icf608ba43019dffad0c708d49076088f2a4b5e126e76b3b2fefa5a0f1edeac7b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I7032c41ce2651dbb03999e2120193d71ed608e40ac2d51329837f3abc0a976b9[0]);
            I0a5867bf6971ed11db3a6dc9af8cb356352990bbc3032878e82b6cb2ca8c402b = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I9a800fae8c9498d12065155e7e781ba817ee2b03ea6540813400bbe438f4691c[0]);
            I56253c88487a75fb5f830a66c0dd3172ff25795a2509eaf5367fe045f9e12b61 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I1dca7dc76f83994b077209eb2742069045e743b6eb763805cbddf87e6a8fcc34[0]);
            I199abcfe7a0dfbaa58ab1dbbb16223bd434b4ce5ed3a65633d506d668aa76f8c = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic16409f8fa42d6ac05643c3943352c03f19cfee0c3068e96d6ca3630b8f2cacf[0]);
            I2ff52a8e46c22b626ca488ae87c88360d413ad08dfaa6701fe7b237d42c2cbe7 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ic66f776d5d728142606f048e3cf27e927f094082fe1dd31f90e757beebd5b5e9[0]);
            Ide088b881c7dabf6e2fab61eb4e5db3ea3750d7b72eb26cb79877bc23429efbe = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Icfe7c47d401f26676f3f8f13e34894792fff7a3881d754de5b4ac1130cfad989[0]);
            I5df56a6a00d4d8ca1c6b1a79e5f0e674482cb9541d86dd49c2ac361d86dcea1a = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ia6852c630d3d698cbe47da7b990ed04d4e0b995b3d765ff6a8146da11e42dea9[0]);
            I16b3b3cdfef91e9cd5ab763bbcbe2188e61f45183118f5c735eff60965fe4138 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I5e5d78a5f1d49833052eb3e84c516dea9f05d6d49879c593f5e0b9745f84fde7[0]);
            I78e49a2727c2f25a14e0f8937e6241f54246c8f42a643dc569f0249384909fb1 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I6454add174b2968c545e831c5bacd6b95b351b7d68448b3fa9c2e5476a8cca35[0]);
            I6563fc7a6bd595720441778baa975487126f50343c92ccba99218e274cf40336 = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(Ie062df11427db764a0e09705579e134d08f4ed2a027e913a43495db5d5fb9051[0]);
            Idc94a4d308c2e301c3d3524f1e20817f9b666827f340874b5adc763970f2efdc = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I2a2245385398379002074dfa174bde148f97bb3bd83073505b550c0c0bbd1e65[0]);
            I3167835472a3c4db7f1b7fbc1895c44e547122e9ad273066e6bdd43bccde11cb = I1dce4d69e7e04f3253de313dcea6b0eb6035abebd2eccf8ed1db45c6548b80af(I862f2564a9e7f99bc8370fe12c1a5e57612d564f1606a21f6a468d558c23fc5b[0]);
end


   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 <=  1'b0;
            I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 <=  1'b0;
            Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 <=  1'b0;
            Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca <=  1'b0;
            I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 <=  1'b0;
            I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 <=  1'b0;
            I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 <=  1'b0;
            I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e <=  1'b0;
            I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f <=  1'b0;
            Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 <=  1'b0;
            I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 <=  1'b0;
            I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e <= {MAX_SUM_WDTH_LONG{1'b0}};
            I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 <=  1'b0;
            Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a <=  1'b0;
            I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd <=  1'b0;
            I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e <=  1'b0;
            I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 <=  1'b0;
            Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c <=  1'b0;
            Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a <=  1'b0;
            I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df <=  1'b0;
            Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a <=  1'b0;
            Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 <=  1'b0;
            I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc <=  1'b0;
            Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 <=  1'b0;
            I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 <=  1'b0;
            I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af <= {MAX_SUM_WDTH_LONG{1'b0}};
            If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 <=  1'b0;
            I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 <=  1'b0;
            I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 <=  1'b0;
            Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d <=  1'b0;
            Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 <=  1'b0;
            If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d <=  1'b0;
            I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 <=  1'b0;
            Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa <= {MAX_SUM_WDTH_LONG{1'b0}};
            I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 <=  1'b0;
            I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2 <=  1'b0;
            I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a <=  1'b0;
            Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de <=  1'b0;
            I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb <=  1'b0;
            If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 <=  1'b0;
            Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 <=  1'b0;
            Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 <=  1'b0;
            I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 <=  1'b0;
            I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b <= {MAX_SUM_WDTH_LONG{1'b0}};
            I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 <=  1'b0;
            Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 <=  1'b0;
            Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a <=  1'b0;
            Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 <=  1'b0;
            Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 <=  1'b0;
            Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 <=  1'b0;
            I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 <=  1'b0;
            Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa <=  1'b0;
            I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec <=  1'b0;
            I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd <= {MAX_SUM_WDTH_LONG{1'b0}};
            I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef <=  1'b0;
            I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d <=  1'b0;
            Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00 <=  1'b0;
            I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b <=  1'b0;
            I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be <= {MAX_SUM_WDTH_LONG{1'b0}};
            I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 <=  1'b0;
            I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac <= {MAX_SUM_WDTH_LONG{1'b0}};
            I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 <=  1'b0;
            I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 <=  1'b0;
            I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba <=  1'b0;
            I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 <=  1'b0;
            If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee <= {MAX_SUM_WDTH_LONG{1'b0}};
            I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb <=  1'b0;
            Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 <=  1'b0;
            I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681 <=  1'b0;
            I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1 <=  1'b0;
            Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851 <=  1'b0;
            Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104 <=  1'b0;
            Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f <=  1'b0;
            I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd <=  1'b0;
            Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 <=  1'b0;
            Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 <=  1'b0;
            I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa <=  1'b0;
            I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe <=  1'b0;
            I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c <= {MAX_SUM_WDTH_LONG{1'b0}};
            I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 <=  1'b0;
            Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 <=  1'b0;
            I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995 <=  1'b0;
            I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2 <=  1'b0;
            Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218 <=  1'b0;
            I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a <=  1'b0;
            Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e <=  1'b0;
            I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c <=  1'b0;
            I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a <= {MAX_SUM_WDTH_LONG{1'b0}};
            I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636 <=  1'b0;
            I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05 <=  1'b0;
            If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0 <=  1'b0;
            I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f <=  1'b0;
            I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea <= {MAX_SUM_WDTH_LONG{1'b0}};
            I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474 <=  1'b0;
            I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987 <=  1'b0;
            I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e <=  1'b0;
            Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229 <=  1'b0;
            I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96 <=  1'b0;
            Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5 <=  1'b0;
            I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icf75206b75ca695f888c3d924d2f1822806f452b5d29a0d6084dbd1c00a15790 <=  1'b0;
            I8d320b2d799e480d78887d5a1483ff7fe5f1a986d75e808863a9085bfc3634fd <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4a1896458491f2613d2c7274b81fbb7a9d405272b871b504455b388a3695acae <=  1'b0;
            I2de3b409715599c65489338e9218150f6c33cd987ece5fdd9c7b2ba5c06d3d60 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If122210c8dc39e7ab2fecb27dac5c167b39ccd9e8e4cd076b2b3b92632357248 <=  1'b0;
            I56c293e90676ea7b55934e3064087e3a4ea95a1c6ee3bd4d606afabce05357af <= {MAX_SUM_WDTH_LONG{1'b0}};
            Iea6e52ee89805cbf2f2a65f695323d8dd7669c23df341897eff049fbcbd1db98 <=  1'b0;
            If32e43e89968b9f008cb77759dc7047519d200c512cb11c105b74c404603fc79 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa <=  1'b0;
            I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2 <=  1'b0;
            Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236 <=  1'b0;
            I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915 <=  1'b0;
            Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e <= {MAX_SUM_WDTH_LONG{1'b0}};
            I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204 <=  1'b0;
            Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460 <=  1'b0;
            I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3 <=  1'b0;
            I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253 <=  1'b0;
            I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idc77bba153be5873f87a4cf88c6ddc6a89bf8aa3ffcd29702126b01053f012f2 <=  1'b0;
            I1ee241dd9ec346bf09b25ccd2f1669be719a1411914d367372a46c8d60cb0f44 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I8674756fbdb78fab124727c8154adc4dcfd4674e3a4d9977d2fff619cbc42e5a <=  1'b0;
            Ia34cf7cdac966a47b902c17ef799ca34f3c17e4f5a410b97d7f07933b977db3d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4a3c7a36a82811aff327ec55776f5077aec859d5557df45568abcbcbb0fc5d5a <=  1'b0;
            If017b6342521fac4000803837465d5793375e9f4b8c2d9fda18843ec7b9e0752 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I931f943f5db8edf3580ebe67b3da2a0cc9a1b68ac6485930d6d9dc792bd36eb3 <=  1'b0;
            I8bc9b50c83facba8db598d0c5c71cf811e181fd16038a08f5aa04f00ff2bed87 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 <=  1'b0;
            I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 <=  1'b0;
            If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 <=  1'b0;
            If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 <=  1'b0;
            If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7b3ff601c78f414f5f48cde79235444d13872a0527c054356b3af150315b0949 <=  1'b0;
            If15a6d2660b407d89dda6c113578519092d37491671c47feae8a7a68565a9184 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I434491ac49be9939ffdcf469991bc3d23ef217b8414c677d78ec9a062e74ba07 <=  1'b0;
            Ibc0fdfece0d7aab4a85b2874a047e1bd390aa826df0d979166e8721339410c39 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icd717b9b3dc725b8579e62b042051399a3b21cc10076de8e0bae480fcd24d607 <=  1'b0;
            I09301323ed69c3f202b9693f2db743880d6e7618dd91405aaef90c34e61d1caf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0c556fb5fa4a1297825cab8dc64089faa86f1cbe67bf106748d927849e16e007 <=  1'b0;
            Icb4397b9bafcf2461e592a0050cf42f2832d3497c940f82fbe98e855a1153129 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e <=  1'b0;
            I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae <= {MAX_SUM_WDTH_LONG{1'b0}};
            I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec <=  1'b0;
            I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b <=  1'b0;
            I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e <=  1'b0;
            I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id3bfe7fc5e0a1ea258f912127a3c77f7cc5ad791dc6166266f64c574b8ed0e81 <=  1'b0;
            If999edef9d50e83e5c53e4715e8f0ae2699c9ad1960e7e16ec5049a8ce0068e8 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I370bb7df3320249e804ee9d3d371b1e82809433e4f7e00f74ea0ab59252f4176 <=  1'b0;
            I17d1cca0614280eb976be22c9779a9238712e3fd3d27b84bc092911227433180 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3d17552542ca2452e4f458fbd0aacb1a5b62ebee4be942ac561b87376658c9d8 <=  1'b0;
            I20665258f942651538aba58d63ca7f531a375ce0ad65c83a1aad4cda0815b334 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5ae887c145ca6af35eef2229e55c297f4b6ffe0a2cc47e55e6dbf09e1f11a9e7 <=  1'b0;
            I5337e70d66d8fb81df05813fd3a172c8337b5d2ca39976efd9dcaeda77844be7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 <=  1'b0;
            I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 <=  1'b0;
            Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 <=  1'b0;
            I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 <=  1'b0;
            I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I00fca56df853315156adf3a6a5cdecaf6256b108f16f65b1e93272f0c7796e9c <=  1'b0;
            I7214b0ea3f1135ee6e703c8e873696254a514ff1e88c32d42757c8ed40a5b907 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia6934e7e07061fec0575e9ceb1910150463d7c530d30091ee48fcc50bc2d0cf8 <=  1'b0;
            Ib9f05dc23ded7e25eec5344da5ea617060c2cb525c22aff7dfc41f86026b864c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic8358c4f85a5a177702d111cdd3e705172bedf92a6d01f2c5d25b5e33c75538d <=  1'b0;
            I4d36f91f636848b5418807d5da024cbeb73a4b63a9b55c2b9bf48f22f2196857 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I2e37b13b583174f0ca14a3fff3bbdd50d584c2a917a020de586b559bb7df4c45 <=  1'b0;
            I55699a1c81182c259ac531c5587702742eb60c998c424e33a62849441a5a94fe <= {MAX_SUM_WDTH_LONG{1'b0}};
            If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8 <=  1'b0;
            I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601 <=  1'b0;
            I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f <=  1'b0;
            I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6 <=  1'b0;
            Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b <= {MAX_SUM_WDTH_LONG{1'b0}};
            Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9 <=  1'b0;
            Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb <= {MAX_SUM_WDTH_LONG{1'b0}};
            Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26 <=  1'b0;
            Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67 <=  1'b0;
            I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d <=  1'b0;
            Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab <= {MAX_SUM_WDTH_LONG{1'b0}};
            I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d <=  1'b0;
            Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70 <=  1'b0;
            I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d <=  1'b0;
            I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf <=  1'b0;
            I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb <=  1'b0;
            Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02 <=  1'b0;
            If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8 <=  1'b0;
            Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436 <=  1'b0;
            If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd <= {MAX_SUM_WDTH_LONG{1'b0}};
            I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2 <=  1'b0;
            I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431 <=  1'b0;
            I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5 <=  1'b0;
            Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f <=  1'b0;
            I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I99fb6dd2fc4414a231a70d23f26ed6b852ea4a563b41d3d8aa364e16d953eeb3 <=  1'b0;
            Id6e462224a7c7f18670d48e3a7c6d35465875f9638395e7dd87b3c494985d418 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If0e6db2779536df3835ac1e3c316bb7d9cf2e88aa7cb70f5b05563886cb4f3bb <=  1'b0;
            I2c0782e7324e49c90f18114dc327f50948f9bf80b906f202a50b101832a88baf <= {MAX_SUM_WDTH_LONG{1'b0}};
            I32eb2fcd88eff04a6295199db748b576fc1d585c2ae058acbf3150711574dd5d <=  1'b0;
            I3d8ccc88024eed4b5d118a6c3b8c06553fcfc8645a8569278e7e7e8d3b41597a <= {MAX_SUM_WDTH_LONG{1'b0}};
            I244e0f2c03df982bd121a8a0240f862b4e0212ab54dbec0984f987577faebeb2 <=  1'b0;
            Ice2f6ae40746fa0bd1c5b2db1aa0bac608899f3ec311d6e8459e126e446f7947 <= {MAX_SUM_WDTH_LONG{1'b0}};
            If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027 <=  1'b0;
            I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec <= {MAX_SUM_WDTH_LONG{1'b0}};
            I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f <=  1'b0;
            I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66 <=  1'b0;
            Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a <=  1'b0;
            I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e <= {MAX_SUM_WDTH_LONG{1'b0}};
            I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228 <=  1'b0;
            Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40 <=  1'b0;
            I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b <=  1'b0;
            I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6 <=  1'b0;
            Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50 <=  1'b0;
            I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f <=  1'b0;
            Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d <= {MAX_SUM_WDTH_LONG{1'b0}};
            I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5 <=  1'b0;
            I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a <= {MAX_SUM_WDTH_LONG{1'b0}};
            I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18 <=  1'b0;
            I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df <= {MAX_SUM_WDTH_LONG{1'b0}};
            I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728 <=  1'b0;
            Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6 <=  1'b0;
            I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0 <= {MAX_SUM_WDTH_LONG{1'b0}};
            I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205 <=  1'b0;
            I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219 <= {MAX_SUM_WDTH_LONG{1'b0}};
            Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d <=  1'b0;
            Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884 <= {MAX_SUM_WDTH_LONG{1'b0}};
       end else begin
          I6ee21517ce790f9f0c0df756f3ffb81e8f92b473aa3a832f200b123f92b8f782 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[0] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[0] ^
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[0] ^
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[0] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[0] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[0] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[0] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[0] ^
            exp_syn[0];
          I8f4ba7628db060b8f44380670c5cf582ed6d7c45c9e8563007505ef6b0d68f13 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[0] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[0] ^
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[0] ^
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[0] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[0] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[0] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[0] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[0] ^
            exp_syn[1];
          Ibd878e938a6444bdbaec2e6ffbe10d2026d17adcb953c1a57250fc3c37cbe299 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[0] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[0] ^
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[0] ^
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[0] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[0] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[0] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[0] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[0] ^
            exp_syn[2];
          I01007020629aa19960e7a943697256ab337edc7b6f5a5557d8699ff724fa81ca <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[0] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[0] ^
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[0] ^
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[0] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[0] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[0] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[0] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[0] ^
            exp_syn[3];
          Id0eb597f7706ccdbdfaede9ac1c6fc24baf34822ac13b31ab45985954ac8e3d3 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[1] ^
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[1] ^
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[0] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[0] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[1] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[0] ^
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[0] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[1] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[1] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[0] ^
            exp_syn[4];
          I43e2980f6c2201e05c9f5b0bac67485fa16e4a35b317a16c96c476da446c5252 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[1] ^
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[1] ^
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[0] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[0] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[1] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[0] ^
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[0] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[1] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[1] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[0] ^
            exp_syn[5];
          I20ddf203cc5258f44ae8ab9eca4a5fcc8828150b1020f9fcd6d4a461e585c8a1 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[1] ^
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[1] ^
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[0] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[0] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[1] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[0] ^
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[0] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[1] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[1] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[0] ^
            exp_syn[6];
          I92afe9a4944fe9569c99a57f089eaf5c6a8916238d085b117ca4b91ce246624e <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[1] ^
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[1] ^
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[0] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[0] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[1] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[0] ^
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[0] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[1] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[1] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[0] ^
            exp_syn[7];
          Ibb0a8078dcaf9a59f2a082e52b2046fd41fffeffc562e2b63d6a511cb549073f <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[2] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[1] ^
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[2] ^
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[1] ^
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[1] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[1] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[1] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[0] ^
            exp_syn[8];
          Ib45d4a2da16f3e153ef2d7f0f00976f1c04ff74e4be02d91347e5948e500e8c1 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[2] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[1] ^
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[2] ^
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[1] ^
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[1] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[1] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[1] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[0] ^
            exp_syn[9];
          I078213d64077ccb9c9d2ab54056912085290b9991570cdf8ee9c993911c030f6 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[2] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[1] ^
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[2] ^
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[1] ^
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[1] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[1] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[1] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[0] ^
            exp_syn[10];
          I30bcbdc869c8ff6580c51d6e19c0075686b84789339117bb505a94883b2421f7 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[2] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[1] ^
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[2] ^
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[1] ^
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[1] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[1] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[1] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[0] ^
            exp_syn[11];
          I41f8ecb76f361e6ba95c167daa463c26ca322e1003fe4cd81a883c203ba32c2a <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[2] ^
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[1] ^
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[2] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[1] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[2] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[1] ^
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[2] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[2] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[2] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[1] ^
            exp_syn[12];
          Ia72a5387982eeb074987759a03534f381a7686a3a0dd37ee976e9d24b35181cd <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[2] ^
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[1] ^
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[2] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[1] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[2] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[1] ^
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[2] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[2] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[2] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[1] ^
            exp_syn[13];
          I5a06e76abd371e4c41d5a3e8c114cd2f00fd83d0e4034a50337a069a11fc342e <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[2] ^
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[1] ^
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[2] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[1] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[2] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[1] ^
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[2] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[2] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[2] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[1] ^
            exp_syn[14];
          Icef503053b3935af23f4fd15a4153c10087004244deecba16de08755d47c22b0 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[2] ^
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[1] ^
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[2] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[1] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[2] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[1] ^
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[2] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[2] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[2] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[1] ^
            exp_syn[15];
          Ifa579c9a4100b0deffd10b8e7117dee8e314e3d5fdc0901374733071b654226c <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[3] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[3] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[2] ^
            Iea53e5522afe762dd4185f0262512abbb94b905893974c13e954df5553942b1d[0] ^
            exp_syn[16];
          I9c8783fc0fb914087ba39c03d5af75540509a4ab6843daab77eb3655933dbb1a <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[3] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[3] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[2] ^
            If481e9fd41cf8181d432f397381b8376d9da7ddfba17b52e65e301e74c3b9b0d[0] ^
            exp_syn[17];
          I73dc56690ada4fe5416b75f9e676fd034467304bb80bc3339d9b2ffc19d235df <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[3] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[3] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[2] ^
            If2e4ac195be838db9dd7b062319aba299887896862f1a340013226fa025b18fc[0] ^
            exp_syn[18];
          I2c9ed4999c6abbae39c66c8c732e89c5a83159e42c7496d601357dbf09aa738a <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[3] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[3] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[2] ^
            I40914301545dfe0b6673f76e0dc0d1ab3968ca3b18fe8f4ff63d5623c31bafa7[0] ^
            exp_syn[19];
          Ia3849a09fdef32ee3bf8f8bbf0b263cb4df93c636a58b6b3c6a4b1f6bbbdd2e0 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[4] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[4] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[2] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[2] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[3] ^
            Idf30e1a70a723113d32f621f0375dd85270da2f7386cff5ef4ff88cfca78b848[0] ^
            exp_syn[20];
          Iadda860d5c46d86f9f258ff2ef03d2fda2a8895f98e777d871cae6ecf682c5fc <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[4] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[4] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[2] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[2] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[3] ^
            Ic246bc24fb918b7c4a32727a332df57bfb205adc05150ae8d944a77cbdc62822[0] ^
            exp_syn[21];
          Iff0b3fe32115773a66986305d4d85789258512650b28cc7f376b72bd69e29592 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[4] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[4] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[2] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[2] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[3] ^
            I6cac9957a16e7cfa8a125b40d8ce42cb7f502078a791b177d9bbe9589b612426[0] ^
            exp_syn[22];
          Ib4fa3c40c0db93bfe166367856df3e9d33f540784a1bd21ce64f5445cc417985 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[4] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[4] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[2] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[2] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[3] ^
            Iee4ad1e7709a56d53cd8b97f587f1f791fb88bf278fcfef32a29fa05247ca13d[0] ^
            exp_syn[23];
          If3bcc5f70b827c253d5c5fc9eacafe53d378c56ceca4255672752ba22b1fd115 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[5] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[3] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[3] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[3] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[4] ^
            I16a4499c48e5c24fd8a6d49ec3bf63c20c85f440c0c897cdb840e9f28fa2e68a[0] ^
            exp_syn[24];
          I24ea303a0372be74d9e3651f637ca159f23e1d597c648c8e79739f512eb52aa3 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[5] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[3] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[3] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[3] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[4] ^
            Ibed209db0bc502e3fceb4ab86ac20a2ebf87c43391a546d592e5aa32709aa8bd[0] ^
            exp_syn[25];
          Ic36af5996eb453d0d437f6593f6887666ce71709175372df5a61a92af56486a2 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[5] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[3] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[3] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[3] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[4] ^
            I05dc9e8db597a2123632b2934d864ae64cab5192401d8f66ebebd95618590ba2[0] ^
            exp_syn[26];
          Ib00d19f730ebbcac6b8caafbbee3f9a90ea8d779035970d9e81eab829b24649d <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[5] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[3] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[3] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[3] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[4] ^
            Ib309786164a7d646c17533008b3aaf0fd86eda3c5ee167efc2080ef5b26a9ddf[0] ^
            exp_syn[27];
          Ic713b604d3860b1075827665601eb7beee6f865b2ff8d21b526827cc9cf0cc99 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[5] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[4] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[4] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[5] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[2] ^
            Id9bbd0f5c16ba0ffae6a0e5304e1726b97df06f06feaccbb1bbcaf0e01be3823[0] ^
            exp_syn[28];
          Idab8ddf0545b142b17b765bd223c184c14a2359d62d0d80f81dbdc0ccb47676d <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[5] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[4] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[4] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[5] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[2] ^
            I4294b001f220e009c2a65fbf8b36ce1d8961c317ae8ded31cbe5aa288191e009[0] ^
            exp_syn[29];
          Ieb27f787cb12da2f99d0a2cd05bde9cb14ad9cbf09fc28f353ab3aa95cb271a0 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[5] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[4] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[4] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[5] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[2] ^
            Id1fe66d1340965020f513e73a4f77d18f4703c194c3954d40a7f1bc37fc1342b[0] ^
            exp_syn[30];
          I82ca84f5350eb6a25c6bd19fd69c2e77591b7ce1527915d2e163f2faaeacda25 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[5] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[4] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[4] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[5] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[2] ^
            Ie95c9af987f352eca30c8546d306af7cdada8d2a8037200d303e6afbd5a4f448[0] ^
            exp_syn[31];
          I23b9b0e15031b325365ce3eb3fbb3f477eab0176485c78ac75c182abe62e1fa2 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[6] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[6] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[2] ^
            Id34d005cdd89bf304f95101c6fbfdd40d6c0b1742b5f3bee3bf043bf88c3d063[0] ^
            exp_syn[32];
          Idabd335be59111567e4c3f9cd0c8de42985f8a7ffde2b839275e16363d47888a <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[6] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[6] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[2] ^
            I79d61ad4114817a49b1dc8e9314d9e3be9758d861974ead362ff0ac862d1d77f[0] ^
            exp_syn[33];
          Ibc1b7b9562dde9182b76ba3eff2b99eada4ecc209a724d1f7f4d58e45dab48de <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[6] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[6] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[2] ^
            Icfe1fffea36cf64044389903be9550fe283d4dbb7f1b47aff2005e70765a6045[0] ^
            exp_syn[34];
          I78a73a0e17f8098bf6efc416f1f53a7b06d530fc5312715d2f1459cca79bd0fb <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[6] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[6] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[2] ^
            Ib08cf17b2065d04f587d1a8231ec1e4bbb6b2b15819de8a7efe18b477515ccf8[0] ^
            exp_syn[35];
          I18d1df6ca8b63b773cc5bf167f3d1e5478b87e8196496b194a671dba78027114 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[7] ^
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[3] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[3] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[6] ^
            I21832b7270210e1bb6a23930ad9ced36d3da201d80310263e26eb96bebd23612[0] ^
            exp_syn[36];
          Ib636386b424212a4d33916a582156d5f25f4bac707dbede4024742a53fb994d7 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[7] ^
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[3] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[3] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[6] ^
            I5dcc76c47f3c9129431152fa6f7047be203fc556198b45db15a9991647bb8c85[0] ^
            exp_syn[37];
          I90401740df191294d9164bd7888f8dbac7c43b4b15e8321a6fe9721e019645b5 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[7] ^
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[3] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[3] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[6] ^
            I450f5b0f5d2b96636ae010048040ebd744fc4ca164cd764bb33615741ecaa62f[0] ^
            exp_syn[38];
          I4b3449b045a8a8ecf4b5b1d79ef7c1ea7cc504ec443d5fc51e4e3d6a8608d7e2 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[7] ^
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[3] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[3] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[6] ^
            I35d64df6881fde0d4836aa408258db7cc1bfb2f066abf8c9345670b78c466b9e[0] ^
            exp_syn[39];
          I8d6d77db07f73b8497be0a4b44f3167e9164f5e9713314c8c1d3a10bcbe8f482 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[7] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[8] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[3] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[5] ^
            I11944fb91fa1b1d5f076cc36db77f0f8434f0edbb1236c7a9bcb45f79432ea9f[0] ^
            exp_syn[40];
          Iff84c319baf90d7da7f57283cd971b357f671571e6f8a5423ec7913ea6408c08 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[7] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[8] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[3] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[5] ^
            I49642204473312df5a3bcab2692aa7558f44f21416226675a4ec10b0543cc5e9[0] ^
            exp_syn[41];
          I640309e9c94a5e5bfefc2737e37b7d3e0b980a25b16690150d4b6f70489ec03a <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[7] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[8] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[3] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[5] ^
            I24e0d361a2679430549932a968d7cc25f980275fea5554e3453ed0a652d31caa[0] ^
            exp_syn[42];
          I3e829bf4096e393a222d88e37ddc6d577aeccbd4fda1eef4728d69be2acb38c8 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[7] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[8] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[3] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[5] ^
            I386015f8daacd2ac9cfed376d3418b56ac13f075a43dde939e4056c29565a926[0] ^
            exp_syn[43];
          I85bd6dbb2cea9bfbd7eb6cc1826103f428a95ff58aea3f414fbf8b7cbca47de3 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[8] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[6] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[4] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[3] ^
            I32832b039ae7e6f4b1e38cfdf680e5044e383b921a76189054511ebe5b8c0d7c[0] ^
            exp_syn[44];
          I0a85734265840c5b5ef728cb3e81d8bb18f56608a097555b6b27877077b70557 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[8] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[6] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[4] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[3] ^
            I09fff9b84a38f3d19685f9627d01a7183cf65d72110802f11e8da0e01194bf88[0] ^
            exp_syn[45];
          I4689705a155aac79c9f72e3ef3879b1ca92391021210f1054be51cde00e344d3 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[8] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[6] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[4] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[3] ^
            Ib82c65f09934744abbba984b6e375bd69ce7231a5085bb00ba4e673cfd3aba38[0] ^
            exp_syn[46];
          Ia31dd2b8cb0d6a1f5c8b3517a6da3a845850777c59db154074a8e58ce9ab38aa <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[8] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[6] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[4] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[3] ^
            I8ec5727130bf67c04580aa1b5b46cdf964db65750f2fc9ce55025b1c117b2bef[0] ^
            exp_syn[47];
          I9723a6bbdfc231db541d0ae1c3800f980cd4de117e1b7de89736279039674dec <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[9] ^
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[3] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[7] ^
            I862dddc300df692e8bbf4ca45a24d840e51ac1e975631cf4ebb8337ceefc2eb1[0] ^
            exp_syn[48];
          I56dcf6fed1db254cc17a64bff391cfb0a959071b0b7ee8cd8c727f26dcb69fef <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[9] ^
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[3] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[7] ^
            Id08a37df0c5095196e2d760938c4d0b7e8716c25b55d9a9656d86c2c473f9c2f[0] ^
            exp_syn[49];
          I27a84e81c6cf875715ddc8a589f7d5f7426ffa55bb9d0472d931d6396eed024d <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[9] ^
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[3] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[7] ^
            I40204cd18eb803f82fc3ef933553c6ec41331f6d4a15538c287b8f57adebb89e[0] ^
            exp_syn[50];
          I8a79eaae8d2b04cbda6a7cc18c5fd0c1b5514a8ce22f65c9c8719485ed38cf00 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[9] ^
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[3] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[7] ^
            I677f733f4e801d99dc2fd1987683a7ac6c8609d84da6c95b8a7056ce07845665[0] ^
            exp_syn[51];
          I7b1b82b93dfd54281caf7fc41c41f48508e6435859f467c564a835c8550fbe1b <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[9] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[10] ^
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[4] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[4] ^
            Ifeb10787a88bae5943b616e3bf751faff5e7eea80e45e24d60a760f4d6b0154c[0] ^
            exp_syn[52];
          I45f134dd80c1ff780d4ca1baa0ae88fa5d24c1b83c07a8dfb951a1b602dcec10 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[9] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[10] ^
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[4] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[4] ^
            Iecc97eedc286cd1c3d301e35036e81a10d164d59da9252a92ca5f355a828367b[0] ^
            exp_syn[53];
          I63a558b4ee8e45aa77032388e162cc308e5515884cadba34a9763c655e566528 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[9] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[10] ^
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[4] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[4] ^
            Ia9a21e6f22a6cc828e041980ab142b418938a92bf8e868216402a46b8c614a19[0] ^
            exp_syn[54];
          Id827df6a528de116efcdc6a2886c61f0275a34c68943ca31f08ac689d6c7e7c1 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[9] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[10] ^
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[4] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[4] ^
            I355f4f82732333ae56692d1c7ee89b368d938d9ce1d5f806be7e46482c10e19c[0] ^
            exp_syn[55];
          I771d38aeac495f434ec620f504f84dbcf29157c8eeeac8e9843e27cece5069ba <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[11] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[4] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[8] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[5] ^
            I9b2ce64b97ca55921bacb9b6aa4cdc8da5c1e33db4215a2470b7cfab3693576c[0] ^
            exp_syn[56];
          I0ebe8ac9c29e84c809995823a7432e48950eebefb58e493c1fd4c754d1ef1c56 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[11] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[4] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[8] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[5] ^
            I2d78ac4a4125ec25a02df6484c0ae640a37f915383b72f33b91e87cdf376fdf7[0] ^
            exp_syn[57];
          I75a1978d2861be3b079857bc35373c4c74f5670643a1d5dbc21af88a729ff4eb <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[11] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[4] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[8] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[5] ^
            Id727bdc545af53e8f89be0ac5627d0c0c0f0bd7d75030bcb41f198a4fe9c7d64[0] ^
            exp_syn[58];
          Id1ca10ffee67658ad7ab86e7449b18d0f56cdfc5b1a412a57b952f09a4334930 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[11] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[4] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[8] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[5] ^
            I7661c17a1c73dbca82a6d3bfba2ab85ebb0131c1e513f093e1b0aec54907595d[0] ^
            exp_syn[59];
          Ie62a87320a380a68cb58d498ff82ef4c4f7af32cd26de51987223902ad1f2681 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[10] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[4] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[9] ^
            I553a83634252c50164bdde3576d7e1552a147490d02eac6dfd1140a46b813d08[0] ^
            exp_syn[60];
          I394c2d3dd82bd2343efc9db0df11053484227d7f333072886ce86fbb9c4b8bc1 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[10] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[4] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[9] ^
            Ib450c1ee41d04516060a410bbdfb605f0ce13cd8781596ce5218928ed207de8a[0] ^
            exp_syn[61];
          I04a1da40c42992376de93a54424364de3ec8e973972d703bd5dea2ef6cb84851 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[10] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[4] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[9] ^
            Ica745abd4de790f1cd3e2a5a32a9d0b5edf1b64e85759c49f3b4e51779443709[0] ^
            exp_syn[62];
          I68dd22d008fee3d9e66e9c1e49b040d5cc9346c72bc5f85ddf6cc5acfb7e2104 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[10] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[4] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[9] ^
            I6399b29558311ea40cda1388848ce13bb7593bfed01ca2a10fa5d8ed6700df56[0] ^
            exp_syn[63];
          I002db99720c4560402ff200a83370414346082834bb760833a432a007d35575f <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[12] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[5] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[10] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[3] ^
            I6f529a4dd77f75d9af4350baf53ba61c1e9c5ea6227c26690987d244dfe71528[0] ^
            exp_syn[64];
          I6962e6d857d6953aea6e3c1427e286406f1ec7fc2e7daded155dd966123937bd <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[12] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[5] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[10] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[3] ^
            I7a94e46f1351801c2edf76bf3b70e3b5100b8e6108d60d9341591aa59f4e95d1[0] ^
            exp_syn[65];
          Ieed9c2276f920cbc4c89a9d480e5aec6da11a6d338e7773d16b6bef39eb11713 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[12] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[5] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[10] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[3] ^
            I0b761d71a88d70e6228dcf7325206f840d9da85892ba151c317e06079291fc2e[0] ^
            exp_syn[66];
          I77e5541055e9d48028160913b75de655b90948f684d9b9ceeb11f611fcffadc9 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[12] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[5] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[10] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[3] ^
            Ic2ae521a3a6fef956f28a89da365b0838d535c9f7801a405cf60cc776ba0af2a[0] ^
            exp_syn[67];
          I72aaca7519608a15749334da9efcd7933b42c1a518af152e258057b547fec8aa <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[13] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[5] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[11] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[4] ^
            I01d9f8a8900be1981c601c0ccb45c1f39a0fdc16179245d80fbb2ad6d7060899[0] ^
            exp_syn[68];
          I95b9eb8bef3f6b9982fd2a61853e3d4b18c6cf7b0257c4b09f98aa15fd9abfbe <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[13] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[5] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[11] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[4] ^
            Icdfc2f0ce24f01af7df8a99b58de3a74e1dda0eea5b41ff2c342106cb226abdc[0] ^
            exp_syn[69];
          I63e669d33b348ee1b40df315c4489376a1b691d7dc57e058341155eb583e6238 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[13] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[5] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[11] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[4] ^
            I929ef5474f10c76c4686fb044b2833b6ba1571f2e1c82b6d92cfaadfa44946e6[0] ^
            exp_syn[70];
          I23047f37783376dcc5232f29f2f841d6bd9228d4dec0c9db45e10cfc3f9ee402 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[13] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[5] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[11] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[4] ^
            I55312932ff9d69c8ffa1e42efdb5e775ccb21a8f9e8791b080b67654462e537a[0] ^
            exp_syn[71];
          I08bf8248972f349f1107037e9a1df754ae0981bc9835565acb312b6b620ba995 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[11] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[5] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[7] ^
            Icbdbaf4eb2f30bb78db34a582e06dc91689b9eab2f8fdfe4fbfb41a8cce93ca5[0] ^
            exp_syn[72];
          I1b1b6c2669c041a68c0b0f1db4d1f44e6e684bee9c31a8081d8e632b0f1aa5f2 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[11] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[5] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[7] ^
            Ifa4cbbd5c3ab5e47a7d5135e4dbaf365e79c4c6a806bfae88c9c0e1c9ffe2fa5[0] ^
            exp_syn[73];
          I37d95c5a96c5eb89fde0d74bf754c82b7767f473e1a72b9354d901eeda8e6218 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[11] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[5] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[7] ^
            I2341907334935e19ef0e392216e39bb35c215730c464a85c0e1b804b364b492c[0] ^
            exp_syn[74];
          Ibb76917f15c13b60592d825ab57784cade5ed9d2fcc73570087c24577c8b965a <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[11] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[5] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[7] ^
            Ic0bbaf8314688690b5a15a5613ab149f604a8bfb92a2b9ed014e7ce2757d0743[0] ^
            exp_syn[75];
          I7ecf3d9150397837b07ac1147ea6c0a93a4437ac2f4af7c694dcb64396e8166e <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[12] ^
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[14] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[5] ^
            I19ff0bebf62a994a2b5814ea41289f72cd62a38d2f37dc0027beb0f488926d4f[0] ^
            exp_syn[76];
          I7b242943c0e5f5b5bf86b8e4df7fa60145071bb62621d6f3ed0d1fe58241de4c <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[12] ^
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[14] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[5] ^
            I4f9435bbcce379d6d591547481382ab188003b97877c0f32462ef9e33aa8bc1a[0] ^
            exp_syn[77];
          I66d4d7d027fb853b3892957ce08f8643d986fbcdcb07643a0067714a52c52636 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[12] ^
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[14] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[5] ^
            I9e497e3ee797c274b82ecca58218c47f9b663bcac21b1431b45c17d5e54e5a4a[0] ^
            exp_syn[78];
          I65b7e46668333ad0e83cf9e4ea9755004ce4dc4b9fa64810359c15513cb9fb05 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[12] ^
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[14] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[5] ^
            Ib929181cef39d751d2726a054cd0478d309e58350ecd11d3363ecba8bd4cb7fa[0] ^
            exp_syn[79];
          Id46c0b7f54cbad7f16743a2b2a3e6d9633ad145f14c5fec385ef993a23cad6c0 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[15] ^
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[3] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[12] ^
            I64fa7f4fa09b7909840d8edb83f29f6a2379419e65b80f592b37d8ea00e59475[0] ^
            exp_syn[80];
          I0f68a80a623a4ec3bcc979bc0f041426497a33b0d2c572d5f63ae909e901e27f <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[15] ^
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[3] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[12] ^
            I35beac843abd6268c39acb691d3105a5c386f05461bca8c63b951ce1c2ed07bc[0] ^
            exp_syn[81];
          I26120ecf137675200083e575ac94ab77905163eccb2081b575259f7acb729474 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[15] ^
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[3] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[12] ^
            I9d8fbde44d35c50f5f24ceae6f2e16ca2f280573caeb8a3021b6f69dec3d04b4[0] ^
            exp_syn[82];
          If050aa312bfe6e49f93d40ff3bf25b55bc3bb55120aaf0810fd6a9d02041a987 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[15] ^
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[3] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[12] ^
            I507d851a78a765c18af6d529292384fb4cbb06cfec0e22d516adc79b8ea13c7f[0] ^
            exp_syn[83];
          I7563504da937c8587a7d900c67d3bff551ac013e2bc9b9f59124a94dc318cf6e <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[13] ^
            I26a8fba8171078ca1fc053c98583785cbb1f372207836bbf59bc3dd3a47cd546[5] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[6] ^
            I80fb8d450dd144ffade989cc2cec363cf6bbcdc267f5372163fde38313387499[0] ^
            exp_syn[84];
          I411a087e83c12e95c02d0948c353c2bba94ed5667078d99612373f2d1df55229 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[13] ^
            I08da1ef5ba49c1e8bd92ad043536907eeef52820296fff2713c49c16da973290[5] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[6] ^
            I7844074cddcce1b95a010729a9e4ce2bfc4f7e1962b84af0e0a3cbb2c2c08206[0] ^
            exp_syn[85];
          I70803211043977c58b694cb493a9d0c36e61de5e1b99a39a55f8f6dd31cf1b96 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[13] ^
            I5a740cae2e1c2dd5f3ce362674a9628e450169869b9368f51e409c95965ca6c0[5] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[6] ^
            I88be0c0499713ce396832a79853e9918ecdfed2519fba6fd7c0bae51450478e7[0] ^
            exp_syn[86];
          I2d29552a2cc0e9cf62c62e47f5d62895b8247aa3fe3090d6d5412ba9bfa3fea5 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[13] ^
            I2a5cb52fcb770ea32660a0300222304c341b53622f6ab018487d6add9656401a[5] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[6] ^
            Ib585733bf4c3eb59a772866965420fc7397b01272410cdb701f289daf9549fc9[0] ^
            exp_syn[87];
          Icf75206b75ca695f888c3d924d2f1822806f452b5d29a0d6084dbd1c00a15790 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[16] ^
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[2] ^
            Ida673298c761bab46fb26d4e73caa99f5b3ade7f924d99fcedae4e47c70b5b67[0] ^
            exp_syn[88];
          I4a1896458491f2613d2c7274b81fbb7a9d405272b871b504455b388a3695acae <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[16] ^
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[2] ^
            I60bb81cc7cd9a6212f7b4261a21655accd6cd09e7aaf5f78f7f1f4dec0e8489b[0] ^
            exp_syn[89];
          If122210c8dc39e7ab2fecb27dac5c167b39ccd9e8e4cd076b2b3b92632357248 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[16] ^
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[2] ^
            I85d3c885ce504524ab43daed7bbcb599cd7e5d6d3635cf46e278345134e97e22[0] ^
            exp_syn[90];
          Iea6e52ee89805cbf2f2a65f695323d8dd7669c23df341897eff049fbcbd1db98 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[16] ^
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[2] ^
            Iaa08a49e0ca4f92f38c7f4d115ae1b275e45c42dfa6fd4b6a2ff40536b7f5f15[0] ^
            exp_syn[91];
          I4cd4c48f741aef73ce7cfcea67b5d0d86f1a1d84758985b8403dc2c3f1a27caa <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[14] ^
            I0f5524aac3a86098abf732fe64930469ee7e55af9e1c3be5a50f833b54111c1a[4] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[6] ^
            I197b3231cb1da107c5001075809e9fa75e4089871d473490981a8b44d3ff5e4c[0] ^
            exp_syn[92];
          If177137333d26dad87a8b5ee41a4205216335f82eb4d49ff21d9e1dbf15742f2 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[14] ^
            I5718908cc8693d723dc81a8b7152b3ba9c006fe7e4119a92e372e2ca84c1ca34[4] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[6] ^
            I384c04b75344f97c691f70965d7e08266ab9cd8862e04ba73b502a0f36ac5ea7[0] ^
            exp_syn[93];
          Ib9db7c1bb2d23d3889404f153b56866edffd9faba2b97fb2f134574ff5192236 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[14] ^
            Idbc0c4a1cc951a261d1b4b84a73e63d056381404d40c97d6685e533582bb582d[4] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[6] ^
            Ibf95afb3941a2272d76cd7256d0789f11fb35a3020c3ccca5b099d335d4a2330[0] ^
            exp_syn[94];
          I07d0819a5155f9b5e32c97f318d288db24503fae0b9c8d62ede275c053cf7915 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[14] ^
            Ia1c9a4ae72bfba2ac774f44d7d126aef7540d7b4ff83981351c5b1c272e40b35[4] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[6] ^
            I885622bb1c7371f4afa3e9966f870d2bf7750c2d2280a2a993a5bd9854187994[0] ^
            exp_syn[95];
          I61eb796cb03595cf7b0eb4a5b27eeb04e3fa5fbed30bd6257023e334c748a204 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[17] ^
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[3] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[6] ^
            I719a3e78d6a298f7db920bf7e355f6fca2c46135abb8ccd1cc3ea470912d05c1[0] ^
            exp_syn[96];
          Ied6f12581ce81037303a23d409e752437dc5aee5b4ef55b216b31c315300b460 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[17] ^
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[3] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[6] ^
            I1729b841d155c32b617727459f01aa9a9a6af56de5f464e20e900e3a4da30dba[0] ^
            exp_syn[97];
          Ice6b5524fd074cb7141d8ba75de45a8704371fc2ed9c262e61b65c79dce891c3 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[17] ^
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[3] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[6] ^
            I96affe6d042e09b07278ae45744977fd3719a31fa5d578adaa2b3a66b2c3ebd0[0] ^
            exp_syn[98];
          Ic88e3e9f8a3ef2dd0db0244877e0eafba8a08899da157a97eba6d4452bbce253 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[17] ^
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[3] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[6] ^
            I12e1e01b28d2d443785fac1d0314b477b221b17b715f1153c5379a85b4b5e3aa[0] ^
            exp_syn[99];
          Idc77bba153be5873f87a4cf88c6ddc6a89bf8aa3ffcd29702126b01053f012f2 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[15] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[7] ^
            Ie244ea5cb57e0b4c14c0c8c22592347d1389a6b0f53b821335b821ca5130ad6e[0] ^
            exp_syn[100];
          I8674756fbdb78fab124727c8154adc4dcfd4674e3a4d9977d2fff619cbc42e5a <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[15] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[7] ^
            I5a07f349b1fd7d668d35583c50dfa3ceda070e5dc241bff1ecdddace6624bd57[0] ^
            exp_syn[101];
          I4a3c7a36a82811aff327ec55776f5077aec859d5557df45568abcbcbb0fc5d5a <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[15] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[7] ^
            I6e5f194e3acb27a7fdd060e05aff00bb9fcd0904b3f920d7db0fee84c1534558[0] ^
            exp_syn[102];
          I931f943f5db8edf3580ebe67b3da2a0cc9a1b68ac6485930d6d9dc792bd36eb3 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[15] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[7] ^
            I09780397509ca78f4b4aed5b08cf22d8eae797d1d1864cdba4a951ac8d583c91[0] ^
            exp_syn[103];
          I40b1832b56853e74839a36f0408fddd25acb01f4718784442483b5c96d268bb1 <=
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[4] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[8] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[5] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[7] ^
            Iefcb9b5b2f238005d0f37bc519349bbbc130e3e072814ec48b4edf9c853a6913[0] ^
            exp_syn[104];
          Ic1872549a4bcfecf7bf62d38a0738559c46e0e0f6ba85e8594f4f35caddfd7d6 <=
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[4] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[8] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[5] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[7] ^
            I9835f6f38580d8765566723f5a9adbfb4935af8bf719b3e4918e1b746cf12241[0] ^
            exp_syn[105];
          Ia125f16dc4a04100715dc64f5826e9c8408d966258c5044994acaaf85176cd70 <=
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[4] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[8] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[5] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[7] ^
            I2266ca44e019a30bb553f955a158a5b075035c4b20a0b3fca6a3675ec79b9997[0] ^
            exp_syn[106];
          Idbd0026454a7d04876616102a79fdd8672ed3eb6c3eaaf4645b5cec2d559ab48 <=
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[4] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[8] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[5] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[7] ^
            I684ec077e37638f022f10b5eb31403e6f9117a83a606f2a5013c2c33b8d1a8ab[0] ^
            exp_syn[107];
          I7b3ff601c78f414f5f48cde79235444d13872a0527c054356b3af150315b0949 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[16] ^
            I799cea0d73d1bf1f2ff9fca84cea71f496b77e5e4e14ce5fadbdce5e2e2f5562[6] ^
            I9331428911b817ea45d1b5ae75eb3ee6e05c189785c995e5d2625f12ce4e0846[0] ^
            exp_syn[108];
          I434491ac49be9939ffdcf469991bc3d23ef217b8414c677d78ec9a062e74ba07 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[16] ^
            I8ac76c0af59f4be06d8b28e62de49db77e7f34806dd57faa0ac52a4a90830857[6] ^
            I7769e8ceb72790c37b351c32983860280aef172974d19a2e99348607863a97d4[0] ^
            exp_syn[109];
          Icd717b9b3dc725b8579e62b042051399a3b21cc10076de8e0bae480fcd24d607 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[16] ^
            I67e38e46bf20d0d8c1181b4878fdc69d352bf0e7812c4d69b9e29532c9ce4aca[6] ^
            If09c36408407b246848b29df63e789fd1041815243beb4f27db0e774e853f1cd[0] ^
            exp_syn[110];
          I0c556fb5fa4a1297825cab8dc64089faa86f1cbe67bf106748d927849e16e007 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[16] ^
            I495ea5f19d2de69b2ea53e5733fa163c602ee7042acbdcae4316ae7e2bbccb1c[6] ^
            I533b63eedc528cb36abc0a469b66b144a6ae5122c038eef85d8d0557c3dff3ea[0] ^
            exp_syn[111];
          I48a1b14c1983ebc25d5c14c5e5b72d67d66880fa94534a3755b3382acb5af62e <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[18] ^
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[5] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[8] ^
            I051e3b709db2e7861d31165ec1e5ee679f1e6dffa5a951072831ce479c16f27f[0] ^
            exp_syn[112];
          I41d616edcf5e6c5aea994c4af9ae5befade7d086df4784c48b34f82f3136cdec <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[18] ^
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[5] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[8] ^
            I2fa018ce903921d0a174a63dbbb29eea8d5700b376335b2ba9bd448e8782018a[0] ^
            exp_syn[113];
          I9a8455d3fa03c690c058428cb884d0361efe94d8b64d38cf1f34d72874bb247b <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[18] ^
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[5] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[8] ^
            I36e06c1d77080ff75778f3dfa4ed60e66f9a3bedc39b214e3fdb5b6c21f1cd3e[0] ^
            exp_syn[114];
          Icb2f6a49f67b09c4aaf933f54a7eb2cdcc361a7275c56fac7da9bec3b4be4b3e <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[18] ^
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[5] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[8] ^
            Id647e3bd88fdc7a3642092d071f66f74657c8364937caf63c723f1e027c157bc[0] ^
            exp_syn[115];
          Id3bfe7fc5e0a1ea258f912127a3c77f7cc5ad791dc6166266f64c574b8ed0e81 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[17] ^
            Iaeb151ea1017a9bf7fc9c15ac1a6060295ec9f9c909f973c9f6c641ffa239379[4] ^
            I015b73e7e4bc4c2a3073a304e58d24f5c8c32e90299f004bc0f75eb9e18e6d41[0] ^
            exp_syn[116];
          I370bb7df3320249e804ee9d3d371b1e82809433e4f7e00f74ea0ab59252f4176 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[17] ^
            Ia3182304eb67400ca76d996f150e688ec4ca57d4c571908d08a1e597246246a5[4] ^
            I7c211cef6a581c5a6871d4c9a2b7ba29a9d05d36b0a758106e006caebfc592e5[0] ^
            exp_syn[117];
          I3d17552542ca2452e4f458fbd0aacb1a5b62ebee4be942ac561b87376658c9d8 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[17] ^
            I41a12e5b292f6dd25298b534ebaa166ad2a116a4d483da24d8a78281fe2f1729[4] ^
            I3f2014435aac47a3c807e9ad3f0829179f9285582b7ff2e3bae250a25e800aee[0] ^
            exp_syn[118];
          I5ae887c145ca6af35eef2229e55c297f4b6ffe0a2cc47e55e6dbf09e1f11a9e7 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[17] ^
            I68b2e0390232509539f6920641a75875a9dfeda72fe287283bf7a8bddb85f063[4] ^
            Ib27fb4891a6edd486a99f23a750057de12a5a3e3fc6a5fad7976aa7e961e0c54[0] ^
            exp_syn[119];
          I5621853f87e8f91593763c53ce6cf90dd157c210391d427c5035fd8bc2b8d238 <=
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[6] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[9] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[9] ^
            I6431e46a646bce25e1c4819e64daf3e828c13b59fb43128b507e50e9afa0157a[7] ^
            Ib58cd067e009a5f4b72af8cfb1e5c49c18f51a2ad8880f65aee683bf8ecd40ad[0] ^
            exp_syn[120];
          I106ee8679d74ed324236708bbbbe2cf265bef53c401f440d474cf58825024415 <=
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[6] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[9] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[9] ^
            I201ecc1efb416aab61694ff3ada827a182d4f582fb56c33874bbd610b43123cc[7] ^
            I7e40bd6625b1d7deff82f67d46817c7af70f1da57561ab528b553b3d244b3f1d[0] ^
            exp_syn[121];
          I22325abbe8a13617d40f316e1d098a27762ec900ed8d90794e447f4930b9f4d9 <=
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[6] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[9] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[9] ^
            I59af681bd1c3330e1c4ce73e36a1c8f0225bf85f1bea73ac08cf0de1e671e16b[7] ^
            I01949f24f74578cb63dd095e8ce639ce0d273c14da81e75d00097535e391aa4c[0] ^
            exp_syn[122];
          Id59ce261d8e6b8a9bfad0db8c1376be178b8e5670bae402ac83134005b73a466 <=
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[6] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[9] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[9] ^
            I5b72d3619d5f7dd82681bc6815561bcca9b404c1733bc447ca22f0567cef7c3f[7] ^
            Id8f2a0d3524b27621ca5a576bf16e15789e6257060225da04da2a5fcc8cf751e[0] ^
            exp_syn[123];
          I00fca56df853315156adf3a6a5cdecaf6256b108f16f65b1e93272f0c7796e9c <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[19] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[8] ^
            I6020dcffd9e047c03740cffcdfe790eaf614ea1036a50fefcec9e13e5b5ac4bc[0] ^
            exp_syn[124];
          Ia6934e7e07061fec0575e9ceb1910150463d7c530d30091ee48fcc50bc2d0cf8 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[19] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[8] ^
            I815f772d86db329f78fa75c3326c129ccf0f6c5f383b42ef18033e48d11525d2[0] ^
            exp_syn[125];
          Ic8358c4f85a5a177702d111cdd3e705172bedf92a6d01f2c5d25b5e33c75538d <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[19] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[8] ^
            I2c8a33831a21c4c21dd58a300467abcc82d52e7636a73a12a003a4144d43e0dc[0] ^
            exp_syn[126];
          I2e37b13b583174f0ca14a3fff3bbdd50d584c2a917a020de586b559bb7df4c45 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[19] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[8] ^
            I8c7b9ead4ab28ae2c2aa5185a0746c9cfe9fd90bdd68f2ba05291045a296d566[0] ^
            exp_syn[127];
          If6b00f77d32e998f853ea835083e8e2b86e4309a998d6abad1df9c7af0c7d1f8 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[18] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[10] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[6] ^
            I32ed4ecd4363760151c1accda085c9afa3efe63daf7a312feefc00b804401c27[0] ^
            exp_syn[128];
          Ic8ebb66e8493594b474ced873c423d77da932a2c083cfb4a33d7e9c6a89f8601 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[18] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[10] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[6] ^
            I6aa6d6c6213348ea0cc3e8b207bca2c1db81499441e4ed721ca0ee01ae831291[0] ^
            exp_syn[129];
          Ie3c4b54cbaa7eb2b809fdfd7625bb142935c0aadf04efb0faf3ee5e169adc54f <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[18] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[10] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[6] ^
            Ib4f23d2e5f8c73110ae24212c4ec0e7ef29c09c8178ec3850f061a5b0386feca[0] ^
            exp_syn[130];
          I4e049e88bdd8dd1b5cca1731919505f814fd6944b80b1f4d87098f9f0f95bbf6 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[18] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[10] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[6] ^
            If2be986b27ce8aa2117f87e9a144015a10acf0a07847f83acec2804b9e987e8b[0] ^
            exp_syn[131];
          Idfc2c9ac2b78c70f60f9f434810cb65b59ae840c0b7362e3f2be02f0efe73aa9 <=
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[7] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[10] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[6] ^
            I9f17331c6a9858b60705d889b5b77078042cffe9e956de20eb067ad7e70626b7[0] ^
            exp_syn[132];
          Id30dc6a5499c9df5e9dc33f0a1f3e9cfc0afaf20ea7091c72e1267f237b4ac26 <=
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[7] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[10] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[6] ^
            I2b70416e96231188e62b7bcf0300c4a5b2d2139449150d31414b92ae075aa0e7[0] ^
            exp_syn[133];
          I3b5436d5dae88a759148c649aa25a4e92e51ac64ca855946d09cceb59cc45e67 <=
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[7] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[10] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[6] ^
            I29599a1dac362c87f4780a94478787a718f63401d2051ccbfe543b44e49b35bb[0] ^
            exp_syn[134];
          Ib291dcc993cc84b1e85473f22b911066ee2c287358dc6d55874b0182d4db7a4d <=
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[7] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[10] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[6] ^
            I5ff7defb023005e77164f9f3b852fa60ce897922c6b814015d3436fe1d1b4a44[0] ^
            exp_syn[135];
          I4bf5fdd6e5ad2775331a904855cd1c53f4d2ae153d394b78a81672c30736fe6d <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[19] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[7] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[9] ^
            Ie132a24e667376de85b8fff9a639698df164043422122a8058c968bb7996d3a7[0] ^
            exp_syn[136];
          If5378be1742837fcb2f8df69abf523cf1fdc1c2f93cf79a4196181e52ec1ae70 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[19] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[7] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[9] ^
            Ie8d5dfc9a77dc01055a551c5f37416d0b13ef83428bf751fb9f95c7d10442697[0] ^
            exp_syn[137];
          Ie7f92e3b79bc40605b3a0fcc9789a89b53faade539cb7496844f05e1eacc626d <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[19] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[7] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[9] ^
            Ic94f2b10208cb23bb5f5b1a46c11c3bbae038308b385373cfaad9a18e09ccb90[0] ^
            exp_syn[138];
          I0bea911517dfd41cca876b6850ad21c17d3ffe83e538063923c222a12e627dcf <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[19] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[7] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[9] ^
            I3b79a6c69be124aeea9d1444f9f985201b55ad0d7a4767a01f612eee12a6ad73[0] ^
            exp_syn[139];
          Ibfb5420c0c0672f5f7e436bc49ee2ea64326350f48ce55305d7552da87a39fbb <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[20] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[11] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[13] ^
            Id3ac4bf805d3981ac1eb1b396b3da5c0dbc68754d89668f0a4cf7c6f2a44ddfa[0] ^
            exp_syn[140];
          Ie623e35b03f7d8c8a528e455024539c6f15ef6bb3add5769649f3c4ab15e4d02 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[20] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[11] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[13] ^
            Id77fd99c6146776bfc20804c67ae41b88cb0441eecba4f40b87828956b7158b6[0] ^
            exp_syn[141];
          Ia46ed08fd0edc8f5a85b52d495ae06a5a9c114c4899495b4911b9873e8d890d8 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[20] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[11] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[13] ^
            I650a7220fd4eb743f652c6c1f9431191621f9fb1a5b5d64bb9649b43bad5b8bf[0] ^
            exp_syn[142];
          Icc20dc8421b747d9b250ddef21ad29eb0fd9ee116222ec79513a467f391f2436 <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[20] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[11] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[13] ^
            Ib7417e90e9dc35367f110c364878657dbbf66b1a714d5807e6347095b833c62d[0] ^
            exp_syn[143];
          I00a3c3ed80bdca0720d8bd3d96715651914bd24002637367f2cc7589b124c0c2 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[20] ^
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[8] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[11] ^
            Ie59a4afbd0d65de2149e8c60229bce12b77f8f1b2b232a11fb9714371eced2b9[0] ^
            exp_syn[144];
          I6bbf54966e14a65f2f30dc25bbef2574d93d81ca0f63b01ce942b55f7a230431 <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[20] ^
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[8] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[11] ^
            Iad3f7ae48f752d3ee71320875a2d1d170e879dd5ff51cdfd662241e6a30fca6d[0] ^
            exp_syn[145];
          Ifced21a37808e62ef684530300b9ac7438ca8dcac747ad252e0e81524ca747e5 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[20] ^
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[8] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[11] ^
            I4e9c85ad6975994daf65df213a2d2fa5a6a2abd91e66d9c9a6f540caf4c2afe2[0] ^
            exp_syn[146];
          I5a9b5af651f053ff5d5c925f7ef2bec1ce82e84f056253cc91bd563a51604a4f <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[20] ^
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[8] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[11] ^
            Ic8f9966a2711f4810086d09b86e16ccf0d31339d146ad5c38d34c973c757947d[0] ^
            exp_syn[147];
          I99fb6dd2fc4414a231a70d23f26ed6b852ea4a563b41d3d8aa364e16d953eeb3 <=
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[7] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[10] ^
            Ic1385b7aee4e3b643e13733b56157e3e92e638da28cd1234e275fc9263709f04[0] ^
            exp_syn[148];
          If0e6db2779536df3835ac1e3c316bb7d9cf2e88aa7cb70f5b05563886cb4f3bb <=
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[7] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[10] ^
            I3a173e6b224a6415ad442ae28a0af62756975427859bbcfc0af6c8e5effd62a6[0] ^
            exp_syn[149];
          I32eb2fcd88eff04a6295199db748b576fc1d585c2ae058acbf3150711574dd5d <=
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[7] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[10] ^
            Ia5580120af4590da8aed890f81ca17929e4c998617df957686c095e891649c83[0] ^
            exp_syn[150];
          I244e0f2c03df982bd121a8a0240f862b4e0212ab54dbec0984f987577faebeb2 <=
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[7] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[10] ^
            I58a3910d475757bccbde2da0e6b5dd5723cbe44e1f4d3e71ac2973fd2a03b3a8[0] ^
            exp_syn[151];
          If81e1446aaf4d89bbe8f4df139e2f8b2dcccd5bc4064a9dd2563f8f7cb978027 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[21] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[12] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[14] ^
            I1b76b0f61e714e21a844e429806d641f6a24f0eb19c23a3c2fcfb76baaf3e72a[0] ^
            exp_syn[152];
          I1fa21cef4f98f43dd1729760aabe5bdd99d18d6c1bdd9d7c94a52b31e480e10f <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[21] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[12] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[14] ^
            If0211848e6cda136970069df5b6156d4ac213717491c68ed49ab39d2cffe9999[0] ^
            exp_syn[153];
          I00d10acadda0e23f5b1a465dfa7819d0e468a0e6bd040087be83e6b658429f66 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[21] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[12] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[14] ^
            Id23ae21f713f4f452abcb1c1839b5524c452bb8bb0b6c35683f9bde212bc5f96[0] ^
            exp_syn[154];
          I9ad44282fb2d860dd098372ef20977b875d663be8fd6a829b91fed2e8f410a3a <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[21] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[12] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[14] ^
            Id5bdb0f5a920710b1af7cc3abade245196df9d1ab4b7f26277fd93e1bbee5556[0] ^
            exp_syn[155];
          I6af06ce0a4a38fc28f086ab0c06646ecc8dc0003594bba91a42ef31a8db61228 <=
            Ifaeebbe4060ba1a9c6dc5491a84c59a693b678098b6d0d44a9b89be60a61b678[21] ^
            I1ca9a79fb26bef43750f8144dd9c0abe6d458f66b977f9b3ad3f5d1e241e5960[12] ^
            I0e0b5f415832bf679922ab9cd21f5bf822d96012e88c87ecd764f01c5c4a8a42[8] ^
            Ic72616171e7fb8489fa12cc29be1f74602ff8e4bd28ea085e938da615238a0fa[0] ^
            exp_syn[156];
          Ib3f898b3907dce900bbf00caab13c7ea1ab6165fa3afdf1d6789bc7fdb765e40 <=
            Icdf5c6901dd15ce395dbf3d466634ee1f8c8311c76a9f604a5026c0439ee9626[21] ^
            I71fc01a6fa081380b5aabf5202099e4c6fb2e09cbc4f0bcefae2a98d809449af[12] ^
            I309a898be24c9a7f39df6bfbf4f71af56796fe2ee0171cb4cc28efa118e8383d[8] ^
            Ia09db6bd7cba6c6e15cac4c6ad0d4c98235a7437beeabca1388fb1b4dece5d67[0] ^
            exp_syn[157];
          I0b68932677e37d2db5c6704679015c4783367622955d449e3699315a3c547b7b <=
            I97e644676e20616386f46777a53405899b681dac58b2fe33b8c6e277a9843b56[21] ^
            Icce85bc0469c071a70002660c182c8244e6fa3296877ee8cb25912677f785f0e[12] ^
            I8ea0f084484660e0d2f0fd76e95e9d339c4666926242ece6d7713922cfa1baa2[8] ^
            I15ab76f6e4824af9b3b4f5062e8dd3c426e1ff0c5f68e4733828c710eb7bca54[0] ^
            exp_syn[158];
          I77830c4c901b9552bbe045ec6657868d3a7dcb05e676b2d9b8fbea7860b194e6 <=
            I93b88671e47b887b9cde5820e2625f52ffcf60a71ef190b3bb4fb7f948498135[21] ^
            I1e176de0e36b5a880960755aa26f0d66537fa0631d1c1dc70eace5bda32a248c[12] ^
            I02502cddc81e406eaa2e914f797aca18163cc1579bd2fed2bf17cccc75f99ea3[8] ^
            I12b276cd6b0aa86ca2e28dbb1f4008ab140668e16e4ef96604a6d1741c7f2f95[0] ^
            exp_syn[159];
          I7376a11af3ef04ae4fc2ccf522b3021a7a0911b0113b962fdc9cb92df16a6d50 <=
            I425e824daf703d39d5688f676ba1d11bf573ab0308f1b3fa294b6a7c2c81a02f[9] ^
            I8b810b9b983dda9dd98763d7974cd85bdb7ac4b122f7722747de0fc16eb92c0e[8] ^
            Ia6cb3ab27f7e08f41b22d411918cace07ba49f4159713ee608a47d183024e1f1[11] ^
            I01577c8c0e65ca47449450a8b2455ee84cf5c48bb26a0799b5523258a039ae40[0] ^
            exp_syn[160];
          I3ae29581faffa9a03a77c0aa4e41defde1bf2b3b41d77df706a89427dcf3e11f <=
            Ie0db2b75b39b02f1d15ec93cc5d18ede36e54de5e43fc881df4f513ddaef95bb[9] ^
            Ieaca075b8e83351dd1502d536fac3e43a93029221645835ff9b9ed5022ae756d[8] ^
            I4c35fcfc93d6d7b294e6fb4f974e52152e57f7c88f1f35b15fdb1e5f71b9cee4[11] ^
            I63ba87cd2daa7c3c625d3ff5bdaca7f2115fc2d65e13972a22b2c2ae5b746d4a[0] ^
            exp_syn[161];
          I729e35453588cff0a3e593de8c56f4fd896ae5a667dce5da5e2612b0becc13d5 <=
            I0d8eaffbb780a352a325ef9744d4aab9f387971c879b7a1c89ba486299b31d7b[9] ^
            Id76b9a6257c2c433e187ad259573ecde35765c2f36d037df7a393082b6d4d2bf[8] ^
            I22f2ba65bcf560979fe1ebcf8cb5f7847d2656e04af27f301c12f9f30dbdae3b[11] ^
            I576afeb6020cc0a8e35837b4b96968ed04cd444999558626adac849848fe7c6c[0] ^
            exp_syn[162];
          I6cc425f04fe83abdffa6966dcc37d641a52a856b3a529fbae80581581f580d18 <=
            I16ba9b1e1ebaabff27a138f06408122fefc981f28ed6ea33d6d67e8ca7f5145d[9] ^
            I1e8f8c5b1cf9fbe08826f2b91cc9774633992b6f05f41dc1638a4b45b6578ad4[8] ^
            Iaf4545d6a73a8771635e55a787a716283fef959316b26036c81317109b86b021[11] ^
            I3b8769ce28405c0bb978c458bd6272f10cea5338af4170ce4e93a8932ae8dcaf[0] ^
            exp_syn[163];
          I5e089ded4efa853364abde2f4129e9af2312bf78df4fdcba389dcc74e1756728 <=
            Id08ab516f98a936bab3a6b0034024bd300aa222e1cdf672ab7d787488d9d60e2[22] ^
            Ic5200a467757cc51baebfab422cfaa7587eaac016e02a21eadb8a30604fa361f[13] ^
            If609369445b8b6abe0391dad7636c727ee1da738b47e731d10ef71ecc162b9ad[15] ^
            Ib4638612fcabc0a2c2f2bba5a2b9eb71cdea23575641b3f81fb6220fcaf284f4[0] ^
            exp_syn[164];
          Ib5f5aa8ed397a623c0669f557aba5be4b2a83b629848f9ded73e4d01da06d5a6 <=
            I688d388fa89509f70042a8afac0b9449c34eb72e0209dcf7e93e01b9df1ec129[22] ^
            Icc02fe735d92b91bf791b60d7102ee0f6a91a6308a1d84785c87d79cfb43d810[13] ^
            Ia7c0e82691d34cca9442ed86daec1e54727edff65043ed10ff441d0bc3c3aa5c[15] ^
            I16ea389c88e4591f7686eae3f1988dd5361bf893895697c0ade8627986a9fc5e[0] ^
            exp_syn[165];
          I3d6354eaa36a8b9050fe8f02633cf0ed6da1cdead2507521f18bc2dd4bb07205 <=
            I63eaf65980b11a76bf8b4bc5bb90d0b350665ee5cfe25686cfbdc53a2bfdd856[22] ^
            I64cd982ffe4ff7e84bff41ad4f74272e33e6e4ec8c09f146a2c440ebba8cf4b4[13] ^
            Idaee65de7fa7e042778069b3648e83923dda4edcafd1b4770fee53c67b706cfe[15] ^
            Ia17edf214ab782c25bbab97f6bb4e04b2fc46d41f9a97fcf617418d54ab76a7e[0] ^
            exp_syn[166];
          Ie2fecd103258f8e7459fec436f8bd34851d6255bd68ead4895348058b62e063d <=
            I87147fe3179cb51d7f3d7edb164b35335f6b4d7d90ce589041d3e2fe0046b777[22] ^
            I7f366fcdb65f3a0abd2630961fb80a331052dc1896ba6c6156c4513fd4addf15[13] ^
            I42eaeb8b47d76234958018b4f06b6df1bf53b0821fc2644de55b3e1bbeb7da35[15] ^
            Ibcfba9f1fb81d976955a1fa7101f0b0db16c344c82cc5ce81f50dd3aa2928d37[0] ^
            exp_syn[167];



          I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 <=
            I435bc44b4b8aac5fe9ba3c30a74d51a42250154c16d5750e075057d1743ffd69 +
            Idf3bd173aa5e956e898d5800f3317a1ef71e334901db42b94f9c6aa41c87c2b8 +
            I04257aade4809f3b60c5cd618c5a29008d1b3d7041330bd5c8db7df720da3694 +
            I0e7725af7e163a3f4ee8bf63bcb825b6d62f4b9260a7c68d0beeabf35eea9391 +
            Ia718f1fe0157bb564650d817f5ea7960bd0698409dd04d9b31d54c95a3f90318 +
            If0025a7dfd37802d1a1fb43d82ff871c2867504735093f0ffaa8b0d85fcd4d1e +
            I35ddc6b67ba559d53bf4b297c2cfd82bcc814a88095ccdf7d6f22fb59113ae98 +
            I8be8cfdcda8c42fc83b767d9cdd6af256d434d307b8e324bd533b5b016383bfc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e <=
            Id60b432b19836d2e0919dc2e0201d162d7446434080aff7165fb949aba097f7b +
            Icb9b19c9fb878af708bd3b433b656104d0f1ae64cb5d5a3f8dfbac08da1fdec6 +
            I4bfb42a957ed14280a129921d4d635017b23dab77b121f51abcc5e738114e446 +
            I1ee3ce036ac0c878003d846cdc3fa9f6b5854855789ea575f0005a9c9937c58a +
            I706a44814e015449aad217d9bd9e0056813b075d8e622aaec4dc08a3518cc0e5 +
            I804112f16593c6ce81f6459599203b07642485939c898d78e113353659a62a68 +
            I95b68240d25deb08902e18ba5fc3ed7af68c0a6ae8e629edcf59930ed55c22ce +
            Iaae1f131bd6bb3b2fd8e363e97f6f9e680c7ed035a086cdf2bef5cb7e023c6d5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 <=
            I2e17b8ef0d25ba5beb474e7007ce1fe5f99f6f7cbf24e5241761880a551f3c12 +
            Ie515c89eac4b602d36f70f52a3fd62fee155da2eafac9c1b14bf1917b62bab44 +
            I7da5ecb7bb8a413a5c6c51f0aff1921be97bb5df5d56f6648c27ee4196fa93db +
            I83ded8cd9258de3ae8deb907ae3b813cc228b189df92f42c55a4b0eaf411c106 +
            I23d075a3ac353b3deca0a572e9cbec9b1ae24ffc7f134b36c6f938d949bdcb1e +
            Ia61e8ceb90369d4ed8ed86b9cdf7d4e89056cf4fca5c7e223bdd7b2c5656ac9d +
            I7bbabd42e7ee42c653f61b4bbd72ed2b076dec2c89baaec2b4589bd55b92fa6a +
            I0e9e95de14abaad3f4dee2c74242d09121b496fc60f22dd3513b90860e7d03ab +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc <=
            I7bd679f7d7da9dc0742c725247978f1c14611083c7de896c4c2de108c6766fb9 +
            Ib5d526172ae46c2a06c11e15361cb13141d0ba754320f60ce6bcd97a9e495221 +
            I6b499c648458a2ed0cf0b27d81aeb706a260c5615a8def0ae89a1a44693061c5 +
            Iba5fd100311e883873db0c3474169654308059bc4c43d52479a4515fa85e8900 +
            Ibdb4937356d2b1cd2091a695635cc7c69b694f775f4c4e8680ea49df1ea6722d +
            I238b01744b520f8759a7e466290a15b15b96fc95b4b8a14afacbedb1657f7069 +
            I4909110fd7213171cbddcd3545ba2a0d3a135e723189edadc7c64599fd2f1f53 +
            I929870fcfce11dff715cf2210ad4a4c30db9af500a8d380153f38f0ea2b7c2b3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 <=
            I7cc2cdc76a638cf4fabcdbd60142d7e4fa11f11486c85b7add7d4f9ba16042c5 +
            I9a798d59823ac9a032d0daa203a7bb153e483bbe4fc47083c1d7e4a65e400156 +
            If307a1ee8e5164bac03971d07c03c3c0440857c7cc29df11a751b3bef9bb1516 +
            Iefca48dd9d0f3c717b0a3b081894e93ac451ed275f3cfa7aed675f58327a2d02 +
            I18e5d7f94022748f9a5645c2b0e385407e0f00d6f9ab28a55982fd36330ce524 +
            I727007bc323c90e0c264e5b8688898c0df1bb72c976fbc3513439c14f15b5733 +
            I739fb2ce1dc1a27f40af1c53d575108539718f9d60f83de60531d7bb201685ff +
            Id29a54af13b6045a8a43f741c229ff88d4aeeffef29065cb29cffbd861479f7d +
            I31ef992f17daed0e1947c4d26611e7377d8b3049bb8ae2ffb3d56f3db5f85916 +
            If51ca9faad7b057d5a086daeaf1118808bbaf90b484e38571530cc3bb497dee9 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 <=
            I11abd59187e2db0058526cb1ea58af9061d439139fa151aaa74184499fcfd24d +
            I91c40ee5121cd738ba7213df9bda6130b101385a28d8a5fef6544c86f6bd1e3d +
            I2976810df2af0dd2879fac8afe975126944b2e40a51dc7dd169051bb5086b3de +
            Ic45f0213074aad63c68cf3fe879ad5b0e70a5977f282822ab582ab88ae7236bb +
            I3599299f7f89ed3c6b11b31caa26e6b30553b9dcc1d5968283085959f822a4c6 +
            I2d89506b7ec0311db709c4aba53b749ec1b531bf4bc7867f3866c39a73aada38 +
            Ie3e85438dc476813cea40910227c7d63eb275948fbd481f56cc51656c1bc8b34 +
            I24dbfd322139e6a1964e587f89b06274c35617e961a5f61f90c67ee3b20ff208 +
            Ic1711dd767cbb72abed2584c5bc27d5422882cb4299da3914c684696eded290d +
            I8e6aa1d0b76cee0ce4862aa5d01ee91caa123335ab19a2150e8c4315c7d958c6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c <=
            Ifc131936849b96a3bcc7bed4c38ebe94d51c56feb4e96d25dfbbcc3670568a16 +
            I89ca3ef99e4b84441ed3cd9f386109125b6da2d23485fc22513b1d8ded87f894 +
            I4c871d8c6a677ef8fa6c955524def78e8df6f9f3fdafb141d43db76d4569104d +
            I10a223d797492c10ad8f6aac1cbdae83833e701ae6314ed988ac117debc98c33 +
            I95e467521db517b858e59156f95992ddc522a7d038ac6bbe691a91b567cd35af +
            Ia9f80db3bd889aa11f43f6aa371715d6aadc7d3aeac0e9519f79b787da6e545c +
            I0543957798ccd8923b2a5b736175c6888eb71c1466a1e9cc7d7635701e103823 +
            Id8a5ef9ce42d57c3feb442ca091604f1fc51e648a89794ea3fbe4b30537fd286 +
            I67874ca15a0723ab01392f527151dd5a60a71a0dd16cbbd572fc50a343c684de +
            I2a9f642cd74521fb661e381a3f57eaf539ca18ff62ee2130aa94da51cd13d4c0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 <=
            I96248ed668211f13555b4a086e7534b958b901242794b9978d673726d56286e0 +
            Ied8c84dd66ab8e8fdeb83c6156b8a6f8cbcbee27c41ccdd8c4d199f70ea67e8a +
            I592170f431e8a8e15769fe2e5f3bc43a7c514290149bf9b93a8f3d3a748094a3 +
            Id8cd2e026867692af509cd433fda0fe6a8b5ccb8ed91bad6530d14172dbf7375 +
            I95b908a4845eb4b14e8f933057bab27e44c6a867e4bb02d87417740e3150e018 +
            Idcc1ce57eae666070b5b9984cf69d5d2409ea92b36718906218185325b5611b2 +
            I114dd7172ac111bca494cc4230447a2dc167f12f198288d34cb5311c279a73b8 +
            I30a86fd347fff855a807034e13d6e751b35d4330df8436470af7bb42af947668 +
            Id56cc1c8a7f6213208fea3ab1298a107ea854d908609dbe2358ba954989e1784 +
            Ib1e8234d991235274c74ac026c33d868403b3d03a18a0c674e07dc4f94d614ff +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec <=
            I6d0d8fc19811812bc80267dd50fc4742e9efceded7a9428707fac605fac90368 +
            I9989d555a1c808f108dd152608d93b00d7a396de9492733ffd5165700c869840 +
            Ibf9f290605da4b6295c786c6ebc135cffc80a3352b42e1d841ba5f6fbbf06cc8 +
            I2fef37935343317384b1d29a04765327533fd87d4fe82a74f24b8196b3dffc92 +
            I1a6ae2cf67f356fae1ec533488e09c6696277823378b06751db7ec97115d9c00 +
            I9fc15e538a85dde7207e48d484f796d96ac712463c802b6995b216e71fb74d93 +
            I3c03db46b6474bbd284be2e345d2fae9939f0925a62da2ff9b1e2f3632740b0c +
            I7ba56fb0b187c50e86b74d8dfa7d7b3a1e2bc341cfb56a6343de1e7bb60742ac +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b <=
            I78023336da442165a8be56b4ebf7b41f4bb48bbc2b05c308dcd344c8f36c476a +
            I3464299c3a5abaf050c7176e4c0e17ade3cd5d6d86e82addf3e12d662def2b86 +
            I1ae7d02f524c03ca060c3dbc879653486c099ecee485690ce40a355fc1ed843a +
            I3efcac0fab0af81582237cdcd612c8d22eef1a6534816484190db28f3e7f3a96 +
            I877734e2edefa267510037759c9490dae213d2e046beccfe87e16c1aeb5583c4 +
            Ie6ccfd08b7627ae7cdfd608c7054781099d7df5a0f133672db189134161f76bb +
            Ia261f7672256403997417633102f8c1332ae17195bc38faf0fb85c4e4dd14da7 +
            I7f31f363b408908ca5cc070f150594db404279b7c5326f5da9abe8f60138bd51 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e <=
            I03527e99f5c488d7864664f339e2094fced797e4b46101f3c2bbe0b892c2d299 +
            I7def9ddb7ba2e414a44523f17bbff45806f0100ef624a52e91b03022877a7771 +
            I453d1e19585e0fb4fa66d684f0e6b37f56990cf101cc3942d5d4fc7e2313710a +
            I9c3d0fe7d767050217425eadb8e780e5eeeb31239f2f517ae5d122bee4157180 +
            I87c64e9e81da569414617b07e39a7f67b0b76c71643cf7257b7374feb6fc9750 +
            I90a0e50a5730714abafa98a7ad70e64903062bfe6f8deeb528bdd7008958bd11 +
            I2edaebf9e3781f53167708c4854b01219957ff020915c8d2fa7b68e50ede1d66 +
            If0d87a6c6a4dd34bcb5411a845e6e7bc7fbeb0e6a34933f64283c880ca5d3d8e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 <=
            I950415762b14dbc0817ccfb0d09d95d700be57ecc9f8011c6163f84336da6e43 +
            I7b25bf7d9020a7dacab3d15cd039a86780e41ed33520f5272ee788252efd1b9c +
            I465489f86885351586de73a0aed556821e0ce34d1c2cebb67227004b4503eb3b +
            I6f7a9d597443df1a96370dbd5e1c1f9cb563fdc4db1d00fa66e8a287fca9bea1 +
            Ie72b5524b212840dd1e69f4fa41b4955ca028c1ea7fd2f3440843cc2ef6d4be2 +
            Iea55b5544c098ecff239cee665c2642cce17d3b546df6ea3d0c832a118c535bd +
            I730afd6404f505477b32f86185baccd692e9e64865f66f048a93e33d1cac8df6 +
            I567366a85ce4a20ac4125a297426463bc2f2c71511a97bfe2f4a01f6e8da6403 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f <=
            I305dec30cf8323b9af4b0a6d285a31b3f5afb2e79c1a2ea77ce70a4409a7c765 +
            I81c612bc8b32254693a4a0c89fb21865b161dd1673f5610732b31dd5663f160a +
            Ia7d01a6ab6c0646f75030a0bd04a711a9c50dc4674c921680034012e67a0c3ea +
            I2ad4afbffd2865f5c89feff965381fdaf73ac9ba4bc6e802a39014fe554b09ea +
            I600d6bfc6bdecb80f4f9d6020bdba9b4c04bcb359e66e793a3bd6732173d0b17 +
            Ic4c53101c741f07c928018af5696d83f45a29d0e5a9f766bd2f1f1404f3eb59e +
            I481cb000cdc7a32db6aa5a6b0da57b76f53f5bec6ef93d4ee25557e1b12064f8 +
            I9ccd1f3aa9f849bfe7dd9ff5f9de6fff64a444bc5286321a1f0e73e990d6a996 +
            I8029c5b828acc50a3a785cab42ada7d51c82647934a9dac7f4a738920f1a332c +
            I95d408de4742f651f694ccc8f61d215af1e9b9be2b3860dca46c143e03b3ffec +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 <=
            Idde70a085816497aa92518899b882b67eb7989897509c445847e24204f5e978d +
            Id3bae057e39f6549ce13910da61dbb41693ff87efebfd241bd1410d3da7195ef +
            I6ffb18ff0417e140b26d84cece8d23ea507516ebb60dbee4438e9433713c9f81 +
            If6592aef798f1b26c5c6593d99137d00bab8e8631070e89dbc6a3e11c89b3e92 +
            Ia0090ea9b75c69dfca34ac43abee88b20734f7afb9c1d88f95eda3df6aab27db +
            I54feba5563ca84d4a04e3ff7ff5ecf689d26961daf0ce27f0be8988087296fc6 +
            I8b151ef6b3125cf983140726d775d948a253c13f020d3d1e75b585afb979bc8a +
            I8bddc257a28da31b71dac60701bade264fbf14f8377b1f504ef874c72e0d45a1 +
            I96ba46d5aa5ea6b2cc6a43df70554584d43f49a6bb171722373d28a2b0f1caa8 +
            Iff8bdf9ea44924628e777925357dcbe728f0ef4be0a3574965c811485fb57689 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 <=
            Ibc813c005ecf7c077ea48779116cce31bffebb300fab262a78d166c4e270e3b0 +
            Ib33ee0ec338d1389ec9010793383d24de32231284e86a9b03fd2902743dc8a00 +
            Ie57f94a45eba4db3826b22e3eb6acfcfa04b6d0669e22e5b78dfae4e7659b205 +
            I123d4c26243478ad4cff3406be39503c6b378cdefa50bf60249ec03d3a44270f +
            I8954b3335e6848eaec70a960b632233aff75de56bd0bb895e2b4ae49095fe19b +
            I0011eafd50b7df59be2a4f143443c0ca8ea87f9a93586d07292ba02fdc2b9b4e +
            I931537d878467c473ac81aec8f9a7d79f286024e62ada1e5f363b93d6887070a +
            I6ec3df474c20bfab5d99aca971523dec8454a5ad4536765f4f9bcb0c31978cd4 +
            Iff82ae02f527d0eff3c9f8bb9d8fc818cf9bb7e3fac1a127849eea6ba27a62d6 +
            If8c51307ae2c537425caa18b7c3dbbf0530e94ada2a2a600262f57f93bf60d24 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 <=
            Iefd5db28023cae3483fe3f0f1dcd5e302d642a0b5750cfa9940a9a8d6326cdb8 +
            Ie11729721562e4a52a189a242aba934be636847d35de867cf00d26690c69abd0 +
            I3f5dc950ac82420b73e1bc98c8c412f7e91958fbf455413c6a0ea5b2569e078f +
            I8cf1c2115398eb404050fcfc654b198694d3c54eaa592d0d725b15e7937d8cd5 +
            Ia9160306dcccf07d591c6c85cf86175408905d5e1bdfb36206d9c4bb5b917dc4 +
            I390750ab5fb20d9be34ce0e294c95ca61ab6e511578b636301037a34f9bd9c07 +
            I8b5d8146640c84b84d0d6bcb2362fd5bc7e7462e1905b32b998b1f00f2da3645 +
            Ic3d44900d87d02e6912d962514abecacc6e1f20fb71c052d58a896c5524e1703 +
            Ide09a550a1cc61dd543f2dd7a6e38af908474f7c815ab70318871dece429d0bd +
            Ia71d81a2779b6eb5f39fad80ee4e7bbcf394b97657cb094aec163180224939e3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d <=
            I9c110ac43d6a359d54082ce347cfc9885dba985b743aeb66bf25962b4539a6e9 +
            I58ea58692cbfa8283ab19d6e609fe472aeb9da51d3f3616a9069eacfb18b0bf7 +
            If7454cbad692d8d1ed806663944dde3d846b241d1f69736da66374c5e54b8de5 +
            I0217d8dc004467c4c431dbe27dc564c042c33d06a5be72a29ceab927708c4de5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf <=
            I9841a5dd86a1b359b25fb293e74cfbd88b34e11f22bb61170ecc921048620dc9 +
            Ic98b2baa4c4b3d4541ae5e7f9ae0b032d4dee98ebd73901690f561438ecfe5ce +
            I6483bb2ee2f7c35aa35adc7fcb6cf8cd426e048f4aff95cb9f4f732f97adaabb +
            I14102f52e9c6fa58677dbf1260a5049a6c2807b245f123cecfc3f1a413badded +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47 <=
            I15e7d6b702e93b31ac4e46f9ba4cf63da33641629eb9cd414d1e2c8cf54b750f +
            I8ae4ec097c879009d8316e76b0a2ff9f4228310728d8b4dc196543a3976d26e3 +
            I1f749b245e6db4722494bb36009a7da73ca94f408d8a0ca7829b6d5258f78e4d +
            Id71b753d1cf473f4f4bb7718f412471692e08afc0ae9d25e617c2360df79ceda +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804 <=
            I05a7291b0f3122dd9941bdd5ce72362b3b0b1803abb126606c82744979184be8 +
            Ied43949ed7bc9c0c92af912b9e283a3e674d42242e0fe8e3d9132738d512fd23 +
            If434186e818b5a899ad4add63d67ba1dbed823165df4559ee78b39d8c758c727 +
            I443558f78c6ebb16bcd49ca586ea62d2ba12ed3bade0e54ae9bb60f83d2598de +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b <=
            I44089ced0a31e79af650baaa02274890b1f60ac7398745a0e4da4b2242f849c7 +
            I18e4b7dc3295cc6f5968878bde7abe5447cebc77dce83fce47db55be2237efc9 +
            I0f75d5771cfa314d28e188de297b4bb53c2cb732724a630e10580ee5fe87cb23 +
            Id60b48bbf346bf95a242f425de7f456aaba5b3ed35cf16a07ac541ca8f480319 +
            I9d23867d2eb5d9dbcc21e9242aa71e141a2ecad61f5ad2bb69d798b2fdd1873c +
            If5c2310896ae5dfd3f83de1affe79fad0f0b6b2b673efbceb7d296b33a6900e7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 <=
            I4c8a0d23fea7158b5e99eea187df1d25395edf7df1db8482b41dab7a8bc25030 +
            Ib2fff9999fc00e81b173cdaa0737f3e4f711ccd0034a6611e0e9111acff3893f +
            I6ec1c8ffb963fef21e978fcfd0268bc24dd283819081437974fa5a06caa64c25 +
            I7f3447e248449854eb030c79bc32b602d376441a193e25bfcf9b8a0eda83b57a +
            If550dcd8751a8725d597ff3b723c6b5cff949b2e3087c71d36782ea291f7bd3e +
            I7d078740e07b48774c64f6dfd7bb0f56821dd685e014f0b9d4e3b7da45383e34 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 <=
            I26e6175466ec922073d5092cb4168f87cd1289008e4b99400c5b6c2fec3eaf5b +
            Ie6d2cd42fa78c1cbf17c7f18dfb4c0cc5f79f1fb0bda02dc92192252f99dd047 +
            I31adf91b5f31b4232ee24f82af27e02a7ed1f8535c552409f353690340b64b2c +
            Ief01c27ce040b3f50c19615a8f5d9bc8b467c0f88a778888fe186887b19fd580 +
            I4dcd8811ecf9d39f66ab4cf1e07e739c7972e9cf2ef9ff6c0a948336e22dcc90 +
            Ib3562b77830a64f31728e11cc54a6d19b55344891eb82355e3fb4491086e8808 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af <=
            Ia2952eb350b07a9cd76752e1a5f76814ed095eb0ee2a284f221b1c74e38d822e +
            I123e1ea1b1588abf2d5d4ede7027783bfb20d60ce3fdf365b86c9f5c84956a72 +
            Ie14918150ed723163714038f6ffd2c64b07d62079dc03ac8fdeacde45633def9 +
            I4b15e4ecd6a6f2139463d94eb4061a410569136410e469abc38dbf8cc03948a2 +
            I843cc48bafe9c4d2e4647f2909064999da8c2f4d8dcfeaf533fcd12c32c37ce0 +
            If7d42431922752de30d5506e1d501f65453a4754d7cab03976695cdee9c0c9a4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c <=
            I1308b215c5082a0407de73f2273fc035460ca21b553479402290c244cdedad76 +
            Ib96bae85b07ff95f5a6716cad97c765010937888a28ad63b16eef3b6ae93b3d2 +
            Icd850fa1e932d19313713c2d376413e7b81faea883442278fbc700a2238f6779 +
            I02ff320cae73fe5cc67804e552bffba75496861f085869eabab140094a18fe90 +
            Ia6ddd4cda9a70e95a6ff1a9369bb2851b90588337f2cdad6ab43fdd6c6e32fdb +
            I269a90aa42086a30a9b03141bf37e3abea46a1f1c06710baf2d052a5bb404248 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a <=
            Ia6f33a5c8baa6ea053642148b8e414d0b9d17a66f4e71f6e44e1f6c6e3e535ba +
            I5a03d267642091bb2d177a6689d91b995983fde126d703c6474d730b455ab56e +
            If377629f88304a78a44bdac612907792b54c49caf9dbaf85b3061be5baa2f5e6 +
            I225da3a8a67ccba14e13c78ca2ffd83b37ac9a961371f1aa617f5752b1bb337e +
            Id4f16cdf2e148fb2732fdbe215ff0edd44d29c41dff8c5b307ffcb8305832972 +
            Id88de8b0cefd527c486f8239ff6f61d6ff86085e420d2be56ce58f4d82d78a7a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 <=
            I97449b979933d41c6555a04ba5ba6cae73e44b040387a504f6f7e2ecb763ad08 +
            Ib6f695414c34a124de17de5cee8798a33f0968f7eca5143f21f88c228ffa6345 +
            I8e89f3937a947ff09fef0df8085edc1dc09a36d7bbb39027d358384d54088060 +
            I862b7b7769e1ce1579c40d6363e23230c9253630d97fe8abe72b80e8a8b5440e +
            Ia810fbec78dcd5215c217347900257a8f892a4805dc2365ea79eaff74af7e64b +
            I107db18dddc718b9fe7354d0f352f72df94ad4653ab0712d5765a495ec29242d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 <=
            I9f0d592f1a57b1d3e2c206ffe5a79185253205dfe7b20be53091145aa16f9719 +
            I781bae0d109036c417f71e00a3df3440df3cecd691fe1f67c147c4d2de217f7e +
            I288ddea916663f74bb339e7a94ac9c86412f39671ca69dc7ec1da05a1800092b +
            Ibdb62dc1ed705231a9d0a9e819d824f81e62746fd6d9877557622a8293c7cc3e +
            I48c76be33e4d7a127ef1f7eb5f4952f81439eced5be914ff90aac6d963267659 +
            I642c0e5f0768f835a6ca3ee6f65875346121b502770acb1ce833e9aed46d4ddc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 <=
            I4a91f2655f96c11b03fce33601bc8f71a0fef4dc1782f7158126cd8cc5a1d690 +
            I10ecf0f58ee2fd15e2b4135dc03cb4053c364660c6d2e2bd03cfc37aa6d6621d +
            If023ae056e9b4b370bc83a2d5604602f45a01a005bc19a769c874536faf4abbb +
            I32a7df875889c28b6d8f86a42071ad142efd5a66d6328669bcdf1901a225079f +
            I446e1574b1d7bd427fed19be1920c5c29a3276d9ec816ebe1e4465cbb762b1fb +
            Ib699efc076bd227e0138482c43c5fc8cf0d0d87078e063262fc4b537f554697f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 <=
            Ia441ac067e28123cc7cd9d005d0f5a1628da5628d4473db60d61b85c61e8d9b1 +
            I91cff501b877ec0153cf2d85abd12870d65d1aa997a6bea7d653bf387813998b +
            I5fa215eca11a15c7ad85760cc87a0f8e883d02472c7af460b13cbe214a596c62 +
            I5e14fc93aa39853d74e7844854278275828d0f5428f2af96c00c8b0ab141c868 +
            I0d58818dc0f3ed67f1e3a10ddc7cd0592bfcb8cb3db1c329edea24dfb0ffde5d +
            I8e0d77d4d38cb3b1e5ece19e010043e9a4f0802819f3e70f0ecc9440f65eff4b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa <=
            Ibbcaf468c4ded9be4d2d82d059bfad5174f330444c98aadb71831769a32f70c2 +
            Ib6dfa3959980c5d348630e2edd81fdee8429a3003b0a21369b99343bda03e2a0 +
            Ibb72bc519d54383d213250311085f6368ead1c943881ccc23f944e652f934063 +
            I1a1149d160ca76d7b9db443f5095737e563a7b75de7375f9c148f4f4dbe7e7f0 +
            Ifdcd4016757d0cef222265289850476e0e2a6547732f999ca0cd8449f7134bbd +
            I3eaa094e28f19bdbec184b0ba0f3792f90e67c77bd8dff9af6042c5002735505 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 <=
            Id9d184571e769ba27b0a5a10807ba8da3e6ba57ed7d66aad1cd984ddf5cbcbd0 +
            Ib43a705a217dd9f2321c3e61ee116d257d8ad59bff5b4f80435f9dd96a8d04fb +
            I800a86b8eeb247f39df85aba37dbaa93060858c235c6ac6b0912fca85af95477 +
            I0cc63aa921326ebb19427e9e06862cc0a42b375a328061bc7f6580bf3f1d3b12 +
            I9beeb3f92470748db1e059cd6c5a929d1eee2a3ecd0ac097032c74f4134a22be +
            I62b9322a1d5ff38480981e00d8469983588d084289f2f927f3339250b5c35985 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5 <=
            I62d2fe36d10e598efb7f38f4f57e4511d08c366d7df7f51bfbc63eaaf216035c +
            I58aad5a5682b85bf58d67b9b00883f015e4093979fae9138f7dcd813618e26dd +
            I2f928325d150ab718f3b764d3fc4e15d88af5567b4554ef8bbd02f4c3984f544 +
            I2af0f38cbf134ae07c76f06d4aafee537bcdfe91b1c4aff1ae27898e18da5113 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3 <=
            Ic0561c97824b9d5b0d84c33cd05cd4f95b9cacab06eeb5e022b0cecd043c6a75 +
            I17e36eac60eec64de05cb738d1e6055086891ee6fd7d8fb300df4f98a3405276 +
            I30b6c3fe760f221d2861a5b6061034f6dee7320a04cbd7de2a3c728427f927fa +
            Iec6be5ba578c849ae0e4fee9c059ff88c36cfa7c14cfe218cad7f7f1d6744024 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf <=
            Id7d51984757deb5794eccbf50647e7535041a18dc506aa16b4ba0ad36bc66b0c +
            I05782c612bec6ce9c2707bd6cb6efd55e1da4d234be502ac88cd02453c61ca60 +
            Ibc35679e4c52c119bb0ab5c5a485b11a4bd43ceba90f9998d9704d08ca3285f9 +
            Id18c335cef6d5d988e55f6fda5a09a24ee80f4d4755f797a11ee94141b69b97d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d <=
            I272bc7cf289752b36b9811d4ec63f5c17cb40399f39607b00ba51817fad59e1b +
            I343c495ca033301298c16cbb81a11a7f9d50dfa8b93ea9226caa182c6fae8737 +
            I4d6d60296569a9b2a811f8064057743f13fdc60379669472d28df97061ccedb0 +
            Ie85ad3f88a177d67b69eb3a03e4a9d92f7431af9de9ccd06f2caa01f9d144f33 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde <=
            Ib8956dcf80473ed75d04e9fcc74400f54ee0b840fce7500bcd68ea6dac6d4473 +
            I57ae0fac4bc1fada55e48ef9952dd7b81a55414196fc22fb27a20b723832aa84 +
            I1a54a485e54cb6d528feed952641c7e5350f3d386ceb62ddd2778ad179aef345 +
            Ideafcce97c26d412480370ab40d8261f37e8bf0ba68bf7d04f4099a517195dfa +
            I53e788aafc97015db67a8363c91d81d369d80c4d24542fa45faf7833fa4189c1 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 <=
            I0549cd0fd3abf1658d503a09b0baa63d09b1411eaa524e56fd30b12f8498e549 +
            I23f5e95dbae4b1223d603061df9b75b9a9ae8409c6bc4ad1fe23d3f5c7a68bb1 +
            I4df045f8dab91c2eee20a03bcbea586a003659b77d8a6e941bd2b2ead3006d04 +
            I8a5d6a4832abe68ab6e9ae33b1b6026805c5db0d186df37fe623a2d9931b2534 +
            I8f74cd611f5df70ef183e9d4a86b5ac23349be8cb99cd470c596fcaa6ec95248 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 <=
            I451de528c384521cbb78ae32b3d4640b0cb8d507c10e11ff59a74a9caadd2117 +
            I72329ad9fd98258074b92a7e88a88c68f8db57e7d6460e9c29ec7f3cc251de29 +
            I1edf83d193e0825c58f470cb0d4ccd85e3df4652ab68fe3a701a6ee0e8a0658a +
            I67e66b155579d855e0c14e91d2ce1fc6fe1d2f869e4f56b37de5f700d84073fe +
            Ief3910aa326e0d9782566c81ab1cbd09faf46d3552f78d7ef5fc9de1d9c245d6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b <=
            I511b38f7ea620301cc3bfa759ab56a2dac9061fc83fb1281673a6cf276abcabf +
            I61e7244c25e176443b24d592ff4299482d572c1705c3e0a6b44698b5366ea3ff +
            I1d5563063ac8386b450a3a36bb3d0a3586cfd6d11471071685e3f7f897d8eff2 +
            I0c92cee9eb9e3c8300210834a106174a25005d9a468a481e0f594a960b5995ab +
            Idddd98e139a087c7aef3922ea2542dd364c9d30f70665754f751ed88dfbd3701 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e <=
            I533b2cd0b272eac7c3f9005cc355cf85ce73803134a0fe0ec194628c3af0ed91 +
            Ieca82bcdc6bd68dc2a28a3b203d8adaa09f89fbf0df6cacd8656b54b141d758a +
            I207af234897ed272d784f4a9f8850eaaa2fbf47f583ed1f0564201e33dccfb66 +
            Ic336cf50b44edc74db080d1127ba09a4313c0972702200ac5207aae8ce6b1062 +
            I474f7c67e6159d041be6d6f4f96fe58f9b7086757936ebbc86340bcd9cd9962c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 <=
            Ib8b4f3fbd26b51974ecee1565c3d0c8fa7abd94e467a7369a62ceafa7ea5ddaf +
            I0b2c4982c217189306b4f5d3bace84daaa25f2bcd089f5de092f9a7900106c6c +
            Icc13ce9fe63ee1c11fd5dddbf0a294cf6ab7ae703f742a92150b7a77868a5a16 +
            I91e90d84eae561663a2e9e59f79782a78095807b98187add5501500b8c1cb126 +
            I2a1c16f7d4c3261619c325f4b5cfe98993d5957a2ff466bae11c9cec6006cac6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 <=
            Iff259e6b8d77d06a8354c4d1662328284ede633f1ca4ec4731dcdae94e869f66 +
            I873ab672a8d92c69b75cd8e627aaec129f1cd371c9f863a6bf88e3965909a6d6 +
            I062483fac022c2d74cc4bb84d57c636a3bbb67d68dacf0da453e3b5f71ff8846 +
            If4b0b6bcc29aecf6816eab93edb0cb358730913253ae72d15db63ae06b19c52a +
            I881a2d7025d422202455bdff165dd982c2f4953b361f29688e75ccdf9e04d476 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 <=
            Iec33764f14e5b0a736fa76a2313325240a520c065b59c6cdd0f2fc5dc36a975b +
            I19123fb30bb6e02a13f39e3e96af227e63abb1351e53cbb91b8d9a79be96053f +
            Icb88d7eda8505d92744b075a1c229e3c0f6a9ff062bf5cd35f6f84467b451e9c +
            I48ffe541268d63545fa48263d8df3c288af7b2646b4dca546a4dc521aa247651 +
            I8245c1ad016aa3d7290e1097eb966b09c8a38fa5bf62bcb7ef179f448104f47d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 <=
            Ie282d05ceadb0d075cca024b7311a5e477e903295d7928735a3c338287734846 +
            Ia81ab6d41925460c11303075dea72c7fb3fe533d88450c32414823fc5b10bfaa +
            I1ca12951f309a25752defa88fa366a90a13ce83b7fb40610c01a8c11a3c2e59d +
            If2f521cf64a5e19b1f744d41d929a37a37689534d0e564224b128866d853b043 +
            I10206e80304f6e623a256b6042ceca13c691a34ef5b6d67667ab4bb11f0b0087 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 <=
            If787a878ae1cab622e44a13190d301d15d0c7ed9271dc50e997c926071f1cd02 +
            I19b5f6ad3c2f2551b49883fbab077c8e3d76392fa42a5030b1f832917bc2641b +
            I1fd78c97c2a03a51b8d2a3dce2a553514aaeffdc051bfd3820d409da4b8189a0 +
            I16863fd89fef9bef09bbfec8d23ba6d42f4de7902a5928e9b43546b4078fbb0c +
            I50f15058dc2e50a994089de4a0487158352c882d4639449d9db322a05ddcba3f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f <=
            If4cdb00eb64cb9e80d78f3dedd797796f44f471b76f5ea3ddbc6f8521257e4c9 +
            I7af411084739689195bff036e9d5e9a950a7691f7d771d4d406aba4c32d95116 +
            I6eba99f7e39a1779ace2db8cd1806d099e7cf0678ec385baba570209f784b5eb +
            I27737e1ab6f67dba3964412127cf6c91c7a58f6ba77e5b6a9808e2775069ad4f +
            I0604d25b233f4206fb580d729452e9694d4b795553a4a788f993c992bc433b0b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 <=
            I9e89eff507c5a2386876f56afb505a22f00d8c0f8a32635a00501ef8d56ecc6d +
            I63132df742cc353a39f27a7a5a00e0990e9e9e023f5c2a8bd571fcd6dd2d760a +
            Ib9855ec95d5c99f93ad4c5565e622dc1c2d1c4a3b5d0937219172d97ac290756 +
            I387ea75c114fd752ced502cc147dc9ad385dbf69607c04edf81ab74b6867f2bb +
            I5b2860f88d7cbdbc92264ca1bd0f97c610e7b1cf340e2b65832553a1762fc865 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd <=
            I206a4b82a444ed76c846a17eccf6c9ad62c42263b472949cc97f838f6a416073 +
            I37646f9ba79338e88c3d793a27911c88d573dc5c1cceaeaf565606c5b61495b6 +
            I3e73f999bb1a0c087c2d4023920d56b1525bcb43f9d1bbc1b49b57d6c9c55127 +
            I62f27f0dc53be101d8fc7f026a673fd33a5397534153859f45c113e6820e9c26 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54 <=
            Ib5d22b614e704f01c688034adcd70603b8e69658cb66c96fe3ea76bdb323c222 +
            I0b2f8e7646b38057090faea20bf55e51f17d23baa4daf0c16d00e75e4c5f0ebb +
            Ie3cada5731ce9e6c51353952cfb87527bca19aa77436766bdcc843dd92f1cc60 +
            I92cfa50424ddf1ada795366ac6c7b31cbb1b1330486911824b881a1fda443c25 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979 <=
            I876c143c75e838720b2a1ee393f5da5ba08822ea13fa1ff459d68d7b0c0e5cd6 +
            I43bd10e4f520ec08b30e8474404cf62a6ad869cdd1d280a2d221e0d76f228091 +
            I00c96393d166280a0d866d1999d4306a650507c7bc407202924f6684f61e219e +
            I1d996fec699e93fc4ce63060990c6347d998a81f0b3aefd88339d5d620fd152d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1 <=
            I3dacdb67f2492ed12375b671dc593349c75562e936401def91b4391c153fa572 +
            Ibdfea3d72843376261dc3e06e3f19be4556508098d1b4d37c1c4cf6928860719 +
            I67a45b7ce414632252362c1556be0e627757c871c136d8570d4300fa316205d3 +
            I33546fedf41dca9168afd7d6916823e8c24aa3c4a855b93820215c68c807a56e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be <=
            Id8832e8e711bb3e7fe9136084b9832a2677803cabec7f2469144eb3b6d4ee3ae +
            Ibba131ee71ced96650ce76aa4695641a089046f8b8345ba312d6868dfbfb2787 +
            I16778a093510ae433495baf9d2b7a74ad4c5315403d0e8aa39eb09cf508dc201 +
            I72e85032ae85773b79f3a3dab895c9667cd32c6aeb44c000096ddcbc0f7be0d5 +
            I8617f958a4de5cf233240840c770360befaafe599fbec1e351b24baf301ecdbb +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac <=
            Ifb337611e63cb9cee9828aa75fcb6d978249e65bcc8770d51fb4dd1644c96a86 +
            I428333658d20f4417e24a58fe364d5a647332ef76ecb7f15d83dcccf1aeb3d11 +
            Icdad18f8878b4e9645b4f2d2434f913a6e0f732a20a6a750e25c2398a086ac2d +
            I8d10cf5dcbbd1a765ece13156db0ad4651b41cc5ee286720226649a707accd16 +
            Id824ed4e68ef3624b9a4d6c5924b08a7b727df62fc9135c973c5f79768c627fb +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 <=
            Iac435cdd22e5425837ad24bd6141cb357c302af7ee7637e1cc2ac25474cf7506 +
            I886fbef883afc3146952de2fc934131aeb38bc2134c096497981d303594f1f37 +
            I3b3f53fca961a376010d1a5b0c49f91d58b351d0306b8433ac22a70f5a1f1673 +
            I58d3b6391c1720bf6ac7458ce499fe3b0573e8f7f324db1a796d1126e42e57a6 +
            I3d71ea5bb4c4be8ea80abe59367519a071132c913eaa5c6538baa8c3faf243d4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d <=
            I0d6546f557347e1d72c176a40dcb077c9c4c78ed89975154f5bbb3875eb1131d +
            I88e5fe043e16a274d915245b02d2094d05fb7710f6078dd6b33c2a21676200c1 +
            Ia2343365eee39c9305def2bd744d3e44bf20b5bab8a48c6a2d95908f74f3cd18 +
            I1d5510ca99815d74f26804206bac7f1e7eec3727fa89d91b014becb49a815abc +
            I6adbf5489cbaa65213fe0804e7494a2b8be9db9132a6ab7058764a1a53480999 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 <=
            Ifc4886636576352e5307fb1fefefded0d693fd059a3fcdd6b4c9dbab1b908114 +
            I2fbaaffcceb2dc6a4f6d9d34140997b18356dc3803bb0a6c6d5f1b3f980e18da +
            Ic56053af1a36bedb5e1670282ac0a93d782faf76d25a25edab3dadb09a302de1 +
            Ia3690db3bb1809f3df1fcc3a2dd5f807a0ef26c4cf61810b0f9bb590951f8e36 +
            Ib4e392b7b8f87358dd5cdefe7c272531bc6bb1f27bf1411c1a2f4331809a83c5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee <=
            Ib897fb3696e7d68b81ff3c1573f5cc234d32e10d066864ec203487a8e56f4ece +
            I15ba9fcccc2e3aaba7bb5967d35eeecfc3bfa7ce27f82435be6dee9d0a4af829 +
            I2cd11587dc2659cd92fb2c4f894bbd9d252affb93f75c3c691dbb02225b4e887 +
            I241e6ca6efe96759bbb20d710c448c9c322aa3345fcdbedf625e297070af52e4 +
            I6b528ad76bac25170636a86ebaf7efd14ee7159ea2c83500021e39e968786428 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 <=
            I101eb18f34badddefbdefe0c2448e2a8a243e4803ef3244b25365881bf227145 +
            I20ac47b3e52f25ce7858fb7952654107faed4cb5cf3abe1ba915710d1af4c933 +
            I51abe903b403df434eba534a1102cabe0a0e976c047fc5cc97a6c8e73263c531 +
            Ic7abe3b0fe121e025ad7f7802b7800f4097111a1108ad088e869e81e5374c42c +
            I294be7c0765f0d4209d4442136d706edb2080883d5c78a3c71d66b5946116bef +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 <=
            I82a2a0149ccdf627e13b7d422945e626fa268c22b3c30bbaadd0a8de14ddcf32 +
            I0738f605ff9ccae9ae63f8e6fe7a9b537d97e13bf3f23c7b0daa4fc414eb7eb4 +
            Ibfb1cfcf89fe21ebca17ed6bd834fb8567cef4ccfb8f03fd5edaf59000ba0cae +
            I55d5daa0c4cb89aac08ecbaaaec1d6afa2379b277051281d3c15abaa6af05edc +
            Id834a34ad825df7c595e3754b5a5638badf560cfb68ec8de2903e73e88b1a113 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347 <=
            Icefdcbf9ca1f8e02b93f295ed8dbc43258b29cbc0cdf9c9ed5fa60117263d502 +
            I3f3cf1014fe01e02bb46b2e8a19716cfaecfec0e44fcc344107589dc409044b1 +
            I0c851ecaa50ea3e1769828a7f51da7a8c3b0c0a11eb9002b108693f09e60667f +
            I09e3897931014e7bd9540023eb8fe1097e36eb5c51db24357b492a132c3a8805 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9 <=
            Ic3ea8409cfacf50e41b97c65b0440348d06b8f196001ba1fda6348071b47dd23 +
            I99c4a78ad7af699907cae52326915f18ac1a2a6f9d99b2aa71c34d10fa78fbce +
            I4878199f761be0332cf7d653cf1e73cd52f938bf9ca0f32724d499765f313d46 +
            I674ac3fcd5872491a3c412a02e367a9c29e4dac14a8ffe8b6382c60a29fde8aa +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf <=
            Ic9e13fe7c29048953ae3698eb5d214d6b71367a78bf1042dd6b58064a6cc596d +
            I072f20811fc3b3515b7794a416e5ba39cca6a9579de36442fb39771729dffa8a +
            If4f8191d57bfd0311981d36c3836f8da526830c6fe2dae5933650b290075ef17 +
            I9ac796f1901c19aeab344ea2c785af3ce41bd23dffe88b1b5216f8f8c0b16e40 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2 <=
            Idc5ae39b0c3c764ed6d9b7859b7627b97e24c2b4df7d97229a88cfc0c22ccd87 +
            I9e8877d4beab63d4bf103c07e1cd9330daccde2cdd266b2942f56b2a8e8a926c +
            I6aaddd1a59b6e96dd8cdd4a57d8fc03132dde1c5b0bd06dd6f0a240c2a04f947 +
            I0d186e0127f200b704a4585b2fc43ff1a9ab19833a90ac881abde94b2da89376 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 <=
            I18886d5e45fe8011ebcf9a20aebf875a01f1b793a54ccefdbe44a896e92cb0db +
            I786cf639910ac9a90b1abf55f9e3b66d87c4bb98a2c8e38142969ee5aefcf6d4 +
            Ibee0b890887202cb33c8fb07639c7bc536951ce8e661d561d7e7a7355db5f9e1 +
            Ibf0c6b2fd7ba6e86f7cea34ea8434ec5353399651fae6f00cae29cfd32174563 +
            Iae8191d31be3785db5d8e5d328fb2d96b0b5d5ecc7f9d14f0bdd3f61a9bb6781 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b <=
            I5bb2c70350634acbcf64debae260225ea2ef5b67ce5d03f38d56d3db9de687f5 +
            Ide94701dd8ad54a630c6eadc44221ee5786180f247fcaec8a7787f25c4070968 +
            I31d4c202b8434aacebdaf5a60c34d7bf3864a5a7c4707efbd1cc3dd82a9ba59e +
            Ia7c03e6396e5145d0027d0963c1f8b7068636ee262fe31aa442a5512e0d4e99d +
            I4694c593512d9d84542af4ca5b0f3022f9b1433d7d6435ffd4b1e53093bf4a58 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 <=
            Ia249a4e7b5c5f1f4458d969c346e560a28969f33c9b0371c6bb21776d319afcf +
            Id4182b8f05992677e12502bcc058d967481d0dc2c9c4731b657f04696a5b5bbb +
            I9dd21c6b63d36e7dde6f3133ab04263a47559b648e8717de7065e7f140911d3d +
            I9244711e562e8ea7e5e0de1921bdbbc5b64363d51d121922f441d8f36e949c69 +
            I78c5059e528b7671e27f847d6042b3fa707258c664749d857004679c6ff96a73 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 <=
            I7efedd1a063df95cac921f7cea9ceea1ddd1afd3a70289c50ea2a4807310518b +
            I598f53ba5c7ffa41f21af94375843b0b7a911670719edc80705508ae32ac0ddc +
            Icc14287e817338eea415b9f8dae2527d6e71853a49869ea829d1b51aa7013dab +
            I81c33c11a5d878aea61749e54e68c024fda21f27f7f4fcf45e5b042e8ca4c3fa +
            Ic83ed3610853814d7c9d6932b644f9c924fec7d67e303160a3c5b99c625634c0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 <=
            Ib91519b86b75cae1ba5b32dc531cae021a01350f4e184d39373bf5553f89a7f8 +
            I42295332275fc6fcb94c042fbe6b48d3d03038fc27c535c7e63674f58da60bf0 +
            I3db60bf522be36d36bdcc35d1d5da9cff2db6e8f89b179726fabca1a7c67b255 +
            Idfb0ecafd00955b66bbc43f1585659b2fd82fa239ab0274450da985354bc4c14 +
            Ie33f8884c8fca47e2055b28f4398f3207f7ea20f8d0858d2a0699ef2da5a8f03 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c <=
            Iecd27d9347b5f52e83b7d0fbf7e51de4a3711cbece5ee265b12663b77b58914b +
            I97f8487b89684c5c6952770b0468738f72682d6230be6a5a31a92fe50bfb239d +
            I42336bb9a452e51859fbc836c4294468aced58a32a221057096f5119d459edc9 +
            Ia50c90193d9c7ee51018451884df0da92f138710bf95fc32e439b39bea3f3b01 +
            Id140833a04f0b4b903ad4e99046b17f76d4c405703fba227d36342b6f1fdbd08 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 <=
            If81604260c143a45d248461563d4d94edd94bb71d791a637dcd30c5c0cbbb965 +
            I3e014fe75658214d8ffa60f966549b131bff6a16020d7858523ac829b0126838 +
            I0a22f1dc32c83db6603459232e78078eac21f865aabe0b9a03923e63cea874ff +
            I157157e9b85b39f2f22c57c4beae22472512ec83319dd9ac30075b4266761031 +
            I90d7a3c4ac0a18444eceec2569cae3d5dcb3d33d2e46c329068b0d35ad063971 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 <=
            Ifd8d2fce7b2a1f0fa487e5be6c007a21b5af1d79da5447d461cd37c189e43561 +
            Ibe646b6da0465c3fb411afc4e03d45f553cf91e67cbcd46674a0051ac1092e30 +
            Ia28734d68fd59a227094e3d5643b87d918753610e867c1d047d8878bd9a46be3 +
            I7fed914efeb5727bba8c1dd0a5cab385a750a2cd9215923b596d1ae914639761 +
            I5c7c7df860c87ada06c17210746ef84d27aabaa26e9cad20397822629716d4a6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847 <=
            Ia49277306313784711d5d8ff63e6a0a77d3fbae050dc1089c734c826be497dcc +
            Ic1034fe189ea09f2aa3b69428828a2b7dbfe9389dcf48dbdbe0f15b9157f7c49 +
            I06414f803df7c8e59f01524020e09627cb11f3809c3456a9a64655062b110885 +
            Ieef9e0d39f2e213f365af4a6a34d0d2c7d50155e8052e9b1944473641922e9eb +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1 <=
            Icf9f5e717c65afd1b3bbc3d6c1bd960155773ec7790543f56c86637a891decd9 +
            I53a66c670d7345059cea712c026fe8c524e74b030af0de054cf6e053bb304248 +
            I0734166e34887037bf713bdf1df0f7219241551cec455ed45881734727f90032 +
            I4771e59053fbd3e261c49e0be7e742e7cf9c5bdad030b67f1b955e13e9bcf083 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333 <=
            Ibf4bbd894f269bd6e6eaf9511141b91ac61b5dd3e77b4ffd07aa88474f251ddc +
            I7c10e2245efc27a4e2a96467eb4e3fd9c28be5f26f65c560653ff4742fa5143a +
            Ia7a158b91a24000cb6211d129d65e781a4e28b8333f897bb401042fbe17c37a1 +
            Ic8c13812ba09457021ec6f39406b1106dc025551c62da4259930c361f19c3a2d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0 <=
            Iba1a21e329197ff5e399aca440cec6d6bd3d9593c332cfcba84d52d541ff1ae0 +
            I3c91639fa462a2a7e65410080b46408b692ca4639ed17637b1d465f38631734d +
            Iee901b35683b34719c33d63d90b8ae11fbc338a170164aac943fb0b495c92b97 +
            Ic7aae8edebf83f3971440fd0e86e7700ac4cc0c087c9996d55cfecea8c489fa5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114 <=
            Ib5a93c88521f26a686316f032821a4e9540fdd8e93570ff35437df7522d34ab7 +
            I0806d1e2ea1771b325ea80b71fe9223f495a3831a560f579401b4e94b6ed172a +
            I7f1329fd762cf679c07aced91992aea071fe128bc24f06ce88bf49e876578a9c +
            I091bf548253a3b22f92aca6479b70ccb74a5f9eda8bd80e6bc1e059021f04b9f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a <=
            I13f5f01dccbdf3df23c5bf603a9657e161c1e2368cb5cb48b212231d2fba7794 +
            I840289556d82218416d7f8652d40586181f7b4ecedd132450594aac1bc47a081 +
            Iaf763109fb82e88c7ec019f7b9b668f88f84a5d4f760592d2dc9172c75be0aab +
            I5c1c30033bd61b271c765ba00b033a58c6389d4bd353ce68d1b193bc7138baf4 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210 <=
            Ife767fdd58724398b336a58803ca328013f3a8228ede0cf108dcae054001de56 +
            I58cee4a472b2fa2f17266cd6ab55d475f304bbee835aac31ac7879d77b8a23eb +
            I3724769b2a595469f910cfcf1f002009d9fc27808df7e59ce728af9a923726d5 +
            Ia4370635785f2b904fb6ab3b8cdb86fba5445230a9d3d02cd908e04d92726f3c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48 <=
            I26ad8ce808bb26201de4f63afd861583af9abc55c7623bf15bd1808c0b0c2be4 +
            I5246ce1dc41e20a5e4e3312a997e8c5be2d733f0cc95f74caa7e668f9ad2f1d6 +
            I1de9fe186e9fdadc6c62a9c6645dccfd3709778f3243d2a4155bdfa20d27a544 +
            Ie73ab4d16ef614a27522cdfd47f670a38ab58f89bc10c74975cf0b30400e198f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab <=
            Ic4e32c1234be0a530c66106794dc1114e4c88611be106ffde42a7ae486560ae5 +
            I42ba6c66d951bbe03a57fa7a4926d6323f30784fe87de73cce065cccaa9814b1 +
            I735ec7a402f471520335d15ee3415e874f56381a2c0cab5c3a5b21f7d6f71474 +
            I76b8cfe5d3985f3c0f249680ed81aa3b21cd7af725925846e8875ef9e98a550e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea <=
            I668775bd016b2384bb3d1cb0a1e89a76d2af15b2307cc6a5d2e0d6c699b02544 +
            Ic8108e830a58b12b8e3ef4897cee70758d1539ae6609d73b5455b94b0eee5510 +
            Ic5921b5017385aa779a2016014d381a982c32c64d1643e79631a8ac842d5b584 +
            I58919d58783467b7ad0108f86d6260f3c551692d00e6639260a68a7a512d8689 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4 <=
            I9075819cc111daeabcc2ddedb4a4297b1a42ceac8b93213f7f76d0fe87c8c275 +
            Ia187792bad45afcf25df25b18a076d255536e94db8d7bac4df79761df5f16050 +
            I424c57a79fc220d56d1e499af6318dd2a2f4a4ebab1c83cc7762658b8c34479e +
            I0d276f9604ec2b8621a86706ad1772058a29e94902e8eece60e3d07948e24cee +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2 <=
            I98ee0d4994c76a87aaef2967ab6cb88af05ab0a7972d2dedbf115ec19c426fa0 +
            Id5eaf1d953b17df3896f9a30f37363d1a69fe3a956b97d307c895065ff32674e +
            Ib5e2defed9b5fe67a6a551e253cf68006aca5e13092f7e9b53f8186c76a156dc +
            I5463c05b1b55c142012470d627accadd8e34924e77ef6d139b3fbe1db1cb91e8 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597 <=
            I7c6ea337917ea8eb0696c514db7ffb66719763162bdd0b7e0ac764c1ae63d24b +
            If2cfdc638b3cfc13d31615533cea59a4bf8123299239956479d3f1d702ef54d7 +
            Iccb7ca5c2ab8a9a4e3776ef42997d1d645c5542c25ed35b161702ce450f90fd7 +
            Ifca2987d8c7f1ca30013ddfcdb82a888ebbd7bc3dc421f7e3d6806f5f3a9aa2d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0 <=
            Ic55bde9a87033c380a5cfe5736d205c15099a2f2cf440f88472d7f6e65d360e1 +
            Iaf14e804e3bb7cda8e67e39af906be2c966fbab4a6e73b8d60ee7ac5733669e4 +
            I5460bdaa1d2a7c1cb2e75baa2c211593afac76ce5160a620b385393217b4185a +
            I5ff269ab544d2b74059a73d0ffe0492473b214d392d8c2ee760847e6c07a361a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7 <=
            Icbbddd7f07e1deff7aacc0e96a33556b62ba127dce877dea351b421ac8d00313 +
            Ica809c2eeaf6926552d9f811bf16c30146853674185c2315876fb5b2ea6d0769 +
            I0583863d43273e6464e5e65a8714be627f867a0320302382d94ef661b21f73d0 +
            I26a6366fb57427f6a0d87d4cff8a293a0752887e71b829e747c27980a1a3dbbf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566 <=
            I91c159ee16a42dcacaebf8cdac4c59d45d2e93735cffd86620ffaf2b859c8795 +
            Iadaa0bd11c77d7ea8c8cfc4b0c805c5afe6b75f597b03729ef2cb704dfe48286 +
            If8ea1abf5aef298950b84058c5e76029f717309fa685556f09c32b72959f648a +
            Ieb5560e3a4f6a9c4543d941ac57bd3805afa7fa17624e5739e8e639e8d0d0c5f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8d320b2d799e480d78887d5a1483ff7fe5f1a986d75e808863a9085bfc3634fd <=
            Id32cba1cfd5a10024378db5089213ad668054033f8614d1ae09b83fd483a25de +
            Iecf240e8fe5f620bf43121455ba23a715b23f53e049d2a36f4bf52e2a061a8dc +
            Id1b9b5118024dfae0e058f5418c9e988e0a5a598ef7553947de6f92cd7399201 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2de3b409715599c65489338e9218150f6c33cd987ece5fdd9c7b2ba5c06d3d60 <=
            Iaad1ab5e7603d5441b228c5e899eea7781b6f486b836a7b662f38ea832c1b8fa +
            Iecf3e0156bbf76dff96948ab7bf67772773b6bd62bd0e0fbc86a6eea8b05d4e1 +
            I50e1a6fdaffcdf8fa99074f4480dcc21971ba8f5747b24a33232f9152b07af1f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I56c293e90676ea7b55934e3064087e3a4ea95a1c6ee3bd4d606afabce05357af <=
            I317bde7e15c3a4d1456e9653a45d4d574509cca539be5c064af2ea89db634f45 +
            I84cdf374f692a63dab22cd91edd4f71e1aff29b51b06f0bca914f92407bea09d +
            Ieb31a59d63544ea160d3934f0e38e6333f8571e77352bdbfd338d68c437f02b5 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If32e43e89968b9f008cb77759dc7047519d200c512cb11c105b74c404603fc79 <=
            I953a4a4cbd4e6c0ccf4880cec5c947f86d6542f9a7f125d7c8cd71f8665b9ddb +
            I5b143cf694d99dabce0cb40d2d689fd7232531ab3a30888f811171b6aa2e024f +
            I81e45b654bee6c74edb5e034c89bed7151c60a69b554a35710d1b173fe45ea22 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0 <=
            If7fb04f8e3e8eaef8fcc0486d12d1e37a887bcdecb366c1e8b53a3e1cce0637f +
            I8e95ffa3fdf70dc76c935f7d4dde6f39dfba8eb795f7ccc55510ab3caf678410 +
            I31734ccacbfeb8a5c0c30cfc84934f8d1636ce4ecae14fe7809d6aa8df35a9e8 +
            I5144a2cef7d82b7a91f9d83ff8fdea356bb01db215bc167f0c498d55d1faa622 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931 <=
            I8fe688adfc161cafc0777f3c3ac9ae27372603ec55cb3865f90f38f9dbb59439 +
            Id2dbd07db2080c14fd0026396339e31183fb5bb6a476999102300cf81f34b93a +
            I8a61ed94b6198131fccf4feb6be7327f59408e9de4def9c4a155167192c5f065 +
            I67484837f2e585fbb85de404cad8f08ba58bd1faa81b9931f88473d7f4a9a06e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164 <=
            I3af3a7e6138910d118e49b29a6de8bb8e6fbd1cfe13549eb0feea6cd07e6865c +
            I7e12dde03af7a5ae0d05cdc9b29f31ef726c7bc51a7f07e374bfbc0846a24f0b +
            I445cf6fbf071cc76e6fc981d7f2f201d0e09d3f47c1227feaac47fb57a14e85d +
            I4404bf7e923ee1bc0230835c00684d298572238aa8b9602dc48e177464224a53 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e <=
            Ib87cc4d1070a195aa8118b92d29d7c836685de2e44ba1b21388677c8e8a5fb25 +
            I39249b7f0d22c6116a7dfd0c0748123ebb6a9b7f931a492a534702157ab28c3c +
            Ibca42a442c971d363e4f848d203d2782af05ddbaad93e8cbf334328d94a8a499 +
            Ied796eff44d61681c5d5de05933e785d387a97b2430fee26d96b0b24a1a54c12 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a <=
            Ib0978aef78ec9b21853831a81aac1d87a2410594c7839432302eb5fa99a4c0ca +
            I7958c747e1ef37e2995c52178d143af6a5f3acdf7c6d1cae518c82653ec18716 +
            If4927b8f31777ef2940c413336113e906e0e3556c31b9b3233107b88b1d71999 +
            Icd8838ebb43dad19fa96e741b32851dbaf5c469e0591a1231898a7aeb6ecc788 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980 <=
            I9d56c14b3465733b5c5fbff528a7a7d85c918a857257ba8e302ae84a0f4734de +
            I80c4eccc6e6be84f8936ed3e9a9457a862eca015298ba2db70745f25a65a6571 +
            I18eefcf5075eee79120ffa0e5875cbe7632d1db84b1c498107413f14b72820f1 +
            Ic6d60bc06b0eb51b5ff4b8cc0d0ccf55fd8e5c53aab23b3994ca8d094920d619 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7 <=
            Ice9dcc5d9ccd6caf90dda22be9ce113c53c7eb492cfd5e0b237da4f92aac2d7f +
            Ia2aece9bdb39e997b99e491171667091adbee475ea9b1c372ebbec109f9f714f +
            Id059fc689baea934a9f278b1066a92d6aff850608c0797dd7257693cbfa40102 +
            Ia0feb2870e46760bd3c58e5af56a40a73fcc6c9611766c77c4784f88c35f440e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6 <=
            I908d977677aa9b15536027b54cf497ddb8741b339748986180944418fd848448 +
            I050437a5474ba60337593b28d17e2bec5c76d26ea8afeac61be93e8ba0ada42a +
            I4c5882b979d1f315e20e4a8fc06c794c0217b97de2613e193cb7a213c2119c97 +
            I60b4f2cd3f513ded6891a6506d0ec74357660440c94e62f4f7e2f886c1233204 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I1ee241dd9ec346bf09b25ccd2f1669be719a1411914d367372a46c8d60cb0f44 <=
            If7c696b260799e0ccd86bb377086dd1be59c9d94754dc52605d659391439d3d5 +
            I96ace764b2f8db5049595445104a408a641999152f2a6c63d22bc6946c27322b +
            I90b9d06240e2a49693ac4ebe37203439a157a38d068e630c45341d7d677b816a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia34cf7cdac966a47b902c17ef799ca34f3c17e4f5a410b97d7f07933b977db3d <=
            I55e293b2d9539b16ee0f135097b8ec02fc9af54fc96ec3a3058af417b0d04e48 +
            I84744085fa951f13f4fef6c44fb0180e543fa6793e89f4dcb14c3da6b27105b0 +
            Icc84144f0fef09379e456de5410487e7882d373874a686f1b61db92511a91e2a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If017b6342521fac4000803837465d5793375e9f4b8c2d9fda18843ec7b9e0752 <=
            I8dc734304648fe3fba1dc7108e8697cb88b61a2ffa704491b2b9df8cc8354825 +
            I701aa61e04d2787a36f529185ddcc94c832834d38ff92b37456b64ce46c69b2e +
            Ib5ba52b9ecafcedb064e66c38273f7833d0b6d0239a7fff9ef3a0e30d0f77dc8 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8bc9b50c83facba8db598d0c5c71cf811e181fd16038a08f5aa04f00ff2bed87 <=
            I6dd215113f113a81bfa59464b587ae7c95f02c1461664fdb818ce751c240b96e +
            Ia57f6e4dd9ce4389f90c78df4fca73a681df346f58a85f61a74e842427848347 +
            I38a6e64d23e0dc1a449445bf10e786777e978aeab68b3a99dc5335b93c67da45 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c <=
            Iabfa5de761b3413904b919f913ed73bf27f5249b7dc6bf8471a23f06a30431e1 +
            I9f08c1a4053ac65909c96d240c83e15017c81fa41f351b0a707fb7882e49f4c7 +
            I6a5f07e66bbd7e05ab9c5adc7bdc99f269386519a6212431d5793e766239e862 +
            Icd7ce463860bc6f62da8d62b71970658ed2c5d5872a56b8429d9223197ef0ad5 +
            I83b2a186b150fb7290623bd1cbab9d044e9b5c760ed36ae218fb775354e46fd2 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 <=
            I0442e99f7519b58fb576a898b41563a174beef69bb6a525712224f5d767a5867 +
            I698aa30e42ad4f250363d29dfc5117677b19f2da0afa75a013718ac5b9731d6e +
            Ie81fcb1c1ed576d911918860ec73a2b7823bb2d435a0477ef407393052729326 +
            Iba39b0599ed448a7fdb07f6042ef972612b54c7251b256373b30788f64f616e6 +
            I507512179a289ecb7d9ddf5e853bb42798df8129655c06e568e0a4a1d880ef71 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 <=
            I697a55c4cb2dd56ce91465bb6750d05200607607d7eaa0b27accbf7f20ba97c4 +
            I4d316d60bd6537dcf09dd9b7eecd93c86af11ddecc1ee65e4b9d65c136527e0d +
            I0162ff342347e70b1361d5f3ea70c6f872d9b95ede7f80a0a18a69c84b5ebc8a +
            I47d2361b09dd6690b6b0a7827348e9e420d8b97c4b620a4e4928c8cbd84c321b +
            I6182a01d42a30ec5e8883e7d4f5d8f1d657f78052fa4c8ca2c160aecffda456c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a <=
            I7355df30b826dd16e0f1fe3be878df80c2ca672dfd1392e2a81ac34fa3df69ab +
            I4eb359966514f007fea3e135207ab27fc596987f985b8a3ec6bf51dde2ff9e38 +
            I0cdb70836bdb3237ff43b23b1676a274cc0dfcffb214799b78ea02c2b59049fd +
            I4eb03f5790e18ea72980b8c37b602469d6dba5f850ca3721f49279b4e14cb7c1 +
            Id645d98c8a2ba63ba9060280b1810d0ab7120f007f3f174e1a501a1f487190a0 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If15a6d2660b407d89dda6c113578519092d37491671c47feae8a7a68565a9184 <=
            I16ef3abe43350c9096f6c7e597c48fc86ed26a073055b7bcd696c34676529372 +
            I034d52d03f918c91bfc6236c72b0d40b688e2bd353f9ca1f03f4c61449bf128d +
            I6822880688515ff8108fe78fadc5d22b953ce5face9928836f824aad9355a713 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ibc0fdfece0d7aab4a85b2874a047e1bd390aa826df0d979166e8721339410c39 <=
            I3088ff7517eebe83fe5804308d22b8c6190077f576f2e680848092e21116b94a +
            I00e08c73bb2036cde2d53598b9977dd2504934b9ba8b58bfccdd21adc2fd223f +
            I694ec7b5bec025b308c4cb56eefedc2be0842202dfb047b5a94dc749c757bdde +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I09301323ed69c3f202b9693f2db743880d6e7618dd91405aaef90c34e61d1caf <=
            I830406b0cd2e64515811ab932e9ce01d413f0a68ab7939a2fa14e4eee7d04a5b +
            I3adad3708bb709ccb06c77ab54c92b6c6629853f740147fd958e6200aeee81bf +
            I99a4bc7f129030d12eeef0507cf52503af3df70717d1ba9c38b5dd3a5ffcb616 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Icb4397b9bafcf2461e592a0050cf42f2832d3497c940f82fbe98e855a1153129 <=
            I08384d6ff32b692ca710ac4170d45cb5d2e2df509bbc473af140dc50f51fe46f +
            I8a3c94278b7c901702cf1b70e89c1832afee395077555d27badd4e2b6fde0b7a +
            I668aff5da6360f719a2467c5189f3e53e8eeb310f4c4e26f55f8c39e9dcc4be7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae <=
            I257c396883faa57c509e7257bed0829f9ca51f30a1004ce730d48e1e5b40c0ff +
            Icf6fe11d7e6948c0bdb9cd50a0135c3b0fac213aef728b8a6555b7601c51cb7e +
            I3d284d86f6c46162d3e0f913a5a6b0e1f2e34fc7ced6a0c226d5e78da81a0633 +
            I4583579034ed3bcee2ef0ea2b32a4adf0467f78a2770a84da9948e8d366c1f4f +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e <=
            I7ac4d72123feb2b9af1a6c3da5adba445042363194ef471c8761e289178d0253 +
            I4bed271962970c26ab72de275bea4b2fb0565d7e44f15b2a1df631bba9e5d4e2 +
            I8741cd8af2f9c3a548c5c39709d7a186f0953de5af6d09d88901e0083a539096 +
            I86729a880fe730068d538da490087a1ab6789327f964722c9c14bd9b1c2af35b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f <=
            I54b0290e037c2111cfef49e6b33d9a3fbe3e85f8fa8a5c707832cb5477f5c0f1 +
            I2785beda1166504e0b7ea979dbf6c2c5574159cfe36c60fced2dc64ebd05a9bb +
            Ibc54f1c4736e5a4608208441ce8d81831a0b6c7448083d6e6976981f8a38d1c9 +
            I0f8046b4f96acee2bfb4719bbff91b4b1b81c78ac36ec6e95008a3d9cb5ea6ff +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce <=
            Ic0fd25473d5639721dddea090dc037e39e4a0c08776c0a343408dfcfc402fa99 +
            I8f671fbd5e9e240cc2f3a9c60c1340fb4bea46c25cda7ea5e42c7ca0c2360bb5 +
            I4b9dd5299690e88d870ceb4939b7f8fdffc8419431458851a3691de4f78f9f15 +
            If08c85e70828c39162bc16d65747d3d3d0a6176e8db106b262bbadd651f745b7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If999edef9d50e83e5c53e4715e8f0ae2699c9ad1960e7e16ec5049a8ce0068e8 <=
            I113d1ff61779dda7e1209787ba652b8b332fc5811cdc0aae65a304aa89d56766 +
            Idcb8d71f1ea9d314ae8f26e9f4b9e25ed245bad319b9af2f71b035aca6d8fa6a +
            Ia0ee127b17b441cc11d664edf15d370368494e31b52c4865c97a065ef8bc43b8 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I17d1cca0614280eb976be22c9779a9238712e3fd3d27b84bc092911227433180 <=
            I6159ddc580c73acd6e2391f4c6cd9989ebaa8947db61972e4fb97f1e12efd17b +
            Iac102173e8323a836c8f86d266f551fc24ccd14aaf39c7d9ef26c465d38706ac +
            I8c494bcba3ff73ff29d9d388708fa34caa73b883730349aef6c2648a2f5a1409 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I20665258f942651538aba58d63ca7f531a375ce0ad65c83a1aad4cda0815b334 <=
            I2f4a0e474435a97fa5d2d056d9de566288c0624cb094d71685934475b58572f1 +
            Ic96ea379edce04b88c524fd17a2b6fb2283e45735640aa3d8ffc7f1bca77c78c +
            I7ea6f607967e7d251d71b4c4b3dd545a4a9ae8298c3ee2356bbc16ebef06cb2e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I5337e70d66d8fb81df05813fd3a172c8337b5d2ca39976efd9dcaeda77844be7 <=
            I8de3f6aec12696eef7d069510ff25e6e620fc4fdde5f92923a707116da636284 +
            I9c0a341c77ecbc1b3c44afee03ccc5a8f34b1275db9c439eedca9ff61a1a1eac +
            I215148c89dc37a59b3eaf2f38679554281379dc6c8e57718e1c22c091f4d76cf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 <=
            I0b60295163435ae3d3b31e9613d753e7e41fd66c11fdf2e7248d7864e11d9d84 +
            I97a73864c1c919943cec586befbb524fa6d6da6a60e1503bcef8116c646b71a0 +
            Ica10d27b8c94c1e740a2287ef28e5d3fedab4221b391b0a3a1da3a472f094039 +
            Ibf57f9e63049a49e05739966f1ec2fe4520b2959db6fee3a18ead9ca03aac230 +
            Ief3b5e8fee2d099a90990de9303f34d600235d989d25a30b5a7e2654c18b5c3c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 <=
            Ie3806d0fc4177d813aade41ad46537a9a335516135161cb2ef18ce822cb301aa +
            I211a150dd66153a3c2c72be4c24145e4c9f0b2f9a3032fee9233985ca9d2c4ae +
            I60f3a2c7d8e3935c04abc8aa09b0a2ef540f13bc98beefc600fd70aa25421191 +
            I7cd31013bf73ff7f7aafbf06eba3fe8110dc5490a280c2d79ce53c77896f564f +
            Ia2233f4704a9724ec75efe5e31af6807f8f1529f641ec05d053d6a12308f485b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 <=
            Idf57b2bf209c68bfc70fe2759595334fabe3d50dcfc4fef8637586c6623c9c29 +
            I81b8212f2e15845be4d129b192895f659d31a061a3a033bc3ac9ebecc75f73fe +
            I3af491b2352720f2bd378052706f4ce571453d59b0fc78b3cb0bce2d51ce5700 +
            Ic6d228f83da7a1c9a71d8fe70d5adbbab8856e5fd3640d805c4076f5f7d53553 +
            I6754b9c9cc470509e67ba88c2669e1f70666489af9ca14de9fd4e4328d18e245 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 <=
            Iaf95e616f53a061a7bf59bf1128d2cf6a5ef64d24b292671a3124a6e010d964c +
            Ib07af5e0c881985b1aa0698382702f78d3ec7ac69cd0deae7496bc63e519a738 +
            I144fae9c9898630fa027b3237ed3434c76965eef2eb015effa7c8677b19c91a3 +
            I5b480e9176a1bb70ebc65f73af78889d266a8efa7414cb97cc5255a5ca5f01ec +
            I133d5432ba2f64f1ad612b2505fb95ce91962b6ac761dcd0e92f75d1b663d7b6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7214b0ea3f1135ee6e703c8e873696254a514ff1e88c32d42757c8ed40a5b907 <=
            Idaa2e762bb01a89e36234967b22cc76cf290937df9295939bb4c4ad08cb8413f +
            If4c7abf17850a5fcd64bb4ebaef1dc806938542a3bb2b9eee643fdfcfeec23b8 +
            Ifb664074b1a8bb954cb940a11ae4e7de1278edf3614b861ccd83dfaef95319c2 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib9f05dc23ded7e25eec5344da5ea617060c2cb525c22aff7dfc41f86026b864c <=
            I7addf7487638274202ddfd183ba052556f89f82da9e873224c5dddf27d2d5a66 +
            I8952c026089661f4ddd0720f6ab16e46334fc934e6775e7163aad8cf5dec6b68 +
            I76ca3c17438c05fc53f6f7075ff7404c0838f62472ffebd41a61afb1f3ea5dbe +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4d36f91f636848b5418807d5da024cbeb73a4b63a9b55c2b9bf48f22f2196857 <=
            I7925970ac367f8374fe02f6e4c8c339c58808928696f0acaf85d96fb3f202f00 +
            I58db55229ca30218227b598184e85d57a0e3a8b61308f8114cd709232573e566 +
            I27ed900fc3d84c4ab4570c3bb88b5e9a7077389e5fa169cc4e1d606f09c9c755 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I55699a1c81182c259ac531c5587702742eb60c998c424e33a62849441a5a94fe <=
            I46777db6f6f68d76ef34c4a9c585ac04e8a978663fecf72d2dbaea3287dfea2d +
            I6f71faa84bc155810576a85be759d7c06d84dd53b5e2dbc74ab0175e5d64d3fa +
            I3ef4c55a4a3281a468daa3233ccdbe660c46a930220b5c9bd3caf6041008bdad +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f <=
            If50a43f14a383995b16d784cc119d01749fd30928019bea1b7aba0039c4c350c +
            I0e4ad715cc833c775ed97e88f28c4196d28bcee4370205307f4266e1fc572cb1 +
            I1f9214a0b2b730fd678664ec457d15dcc243ba1d68ea198ef2792ac2440608ee +
            I9d323aa17bffd7ea7a66ef99d4d004ce664a0e7e5388ed24a4d45c69a4d9b396 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7 <=
            I88f1c4536adedb4ffea1b595f5fa753329c4aa2187a3245269734a18a122e189 +
            Id9a38b1906060dc5739f9446bb2dd1a6b6603924d4b7889c931988fb52cfafff +
            I5502a12455fae3619e0c2297d5e4a8062415aa3ddd8f0bbf67a73233bb6df733 +
            I8e6a3df905c8c5778e1fd6e75b091c545389651762d9cb3e0d21b20d8dcee6ae +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e <=
            I554ab27e696a028f48da8ad39e2db6668b57ff692603a9562cd7e8780bfa491d +
            I1f070cf569961de917cbd287e7b14a2ad6e04a4474edfb92c095f6e9cea1efdc +
            Ib423f5e14b109a601cf9e9d403a7b5c0ca0de8d665d065d8f317760c5705071d +
            Ic935d033e29fa4baba415347d379eeb1645c65388d3c7c9858ae48f5a098e2bd +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b <=
            I6996b52f42eb9075a634fcdb07fafaf45c5aa99193446869751c4859e7c1f963 +
            I332737561309225f302f64e49e8b3e4aa4dc35344858059b21e146e8cb84a466 +
            I2d2817ad47b56d0a7ff72c326eabc6e2ffb1819a2748ffe3a4a42d3794cf2fc2 +
            I1f212ee134daea9d568f52fcdce6452048326c2dc243c60d25ee71b95ffea50d +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb <=
            I8e8e17839b8f0cf30290c33a60662c784f062950716903854e36856a58f909b7 +
            Ic595c984782ebc89b61fa2a64e994aa66eb4979ab1e30e890886355dc247a67f +
            Ibfb48072643b2cdc460b7a667940129aa243be78b6d57abbd483d5551fa36eba +
            I3a25f0d4a6f0fa33f493d9aec6fc7a318a826b3885a3cccf04e9b1a85bec345e +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952 <=
            I31ea69d26acd05d303178076eb123a7b2bbfeca82c2690c54323889753261f1d +
            Iac3e25273f8b972112775f3aa57274eabadbc2da5eea147328f85a941b959bfd +
            I4b18b20124a63f85e812047188401b685693ae009c87ae337b840a7a3e03f140 +
            Ifbee83b3613941d8ba27021c2fd37d0990a8af8fa3e0399f0f1f8a92ae18d273 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677 <=
            I41b85a49eea9c0d773ecce66f0023338d3ee5a94e14a87c867a74960d30211cb +
            I698accb14122caa36f489e7fc522e39188ee03651ef0c6670eecd60162cf2f0d +
            I26c556de81da143a85c36f6ba98648e110114ab97302046b7aec581a62689a3d +
            Ia1c056993094512262fa3f3d38a2a46cd43eb08114e1af8c48ce2f6705d7297b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab <=
            Iccacefad631e33ec8e54f8261759ca110fefaa6fd9fad08940205708a7180eb1 +
            Idb883f1d90a389f89c3e04f54dac20f205951bba3fd0a00e9432498c4def1131 +
            I5059641c5d09a0369f6237643b75899865bff068e9aa8779d0befdbd53a6b754 +
            I61e29bdef580f4f1057d7b4ffb5bbf37c67d3b8107d7979c2fce643282c7d861 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7 <=
            I6f52a21dd933b23b7565abd508c69070b8cf652dc313689f62c7f04d7acb934b +
            I80c7df909269b691013f9d178bc3e8c896d4d06ef4cc4b0ac42858888ae8b92a +
            I403d7b440509677065b38ca8634080a8edc4c8eae54a9923c50885861866a7d8 +
            Ib07a3587e3bfa70ff5dcb296b8595c5d15cb8a94efb13c3e5cc92cd3be3605ac +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5 <=
            I78d7fbedde9ab5751194c52134dec1b83ea8d48c4ad77c0b3eb952143612ab71 +
            I581a3a40f892233a7bd0dda3bb84e2e46095c27e45d53ed32ef5226f9d25ce43 +
            If15171a1904299c55ffc5b4c9059900188c1c87caca3f4807c4498abe038becb +
            I8c443a2690956ee9d0171ca05534d698f75563cd74ec9f4de33c7e8dabe8105a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093 <=
            I3fe543ea18333fd169c6d6e692a5b42232e8abd2b14072a4daba9bacbe921d2f +
            I7a52610226b8a85bdc6a0b49cd74cc644d2fad0e8f98ee24c46ccd3664d0af24 +
            I9efd4f4bd4d8dfa270cb1c5a2e3f5c6cbfc3c5b672540ca268e0765170e6c748 +
            I5dcbde9462714577263040534f0560b0c126ba001e959add92d0529cbc94bd9b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a <=
            I7dd3baf838ce22ecec10d3c1a3d0dd16582497f9e447038aa46bfd49571fcb4b +
            I0dfd7663ac138a56ce3fe38c03c10675da9e417e38f56ea0fa4f9f1902d725b3 +
            I94ba926e07e8b3cbc5429ff6bf73020e95dda7b7c0059dc10ef646b2980bd80a +
            I3872eb448ad521cf99b3a9d07ecde078320dcaaac45bd387137deaf5dec956b3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223 <=
            I4a4338f7d9bbbf60ef4dc6e821d22619911e41300b49e83d57a0a959218a05ae +
            Id1fb56c160d418b26fe2b51dbe78addbbd2743e7a342e0b6bebd2e8d3cb1ce99 +
            I89b44baf278e7cf024304d7bc6cfa759a735e5da0cf25a96a83e29fa83d12bd8 +
            I144443166f296f7fdfd616492bb4b1fe44e0353fa6b0fc822b3aec0c1ea0c894 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911 <=
            I9d7b0f41f5cd73f907351990b23117fcaae4302a36d194e6953b54d40361f8fe +
            I8beede7aeefea570e5c65a76dbc5ce1f4eb114e444ea9b4636258bcefd9d5f34 +
            I102751a9d577151cf6f780ced3299363623ab308737d8483ccbe02118244d2bf +
            I5445f1e35f9039ef623a77ce395c2a888153749fe8226e9b844b271c1c69d760 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8 <=
            Ib0de9295b071389ca7b6bd34f7c9371614337b0be04ccd9ab9819a8e39ade463 +
            Iae16b002804d17ac9e2c9655dda031f3f0ac10d703bc42079ee2a5fd3ede604f +
            Id9db55519cb1208a2555678410c950b6fb31e5fb04a0ae12d6b0a9de4d750b43 +
            I5d9ebd6a6829c49b0e41f700d29bf8acf06a5dd87192846e5ca204ea8bf563eb +
            {MAX_SUM_WDTH_LONG{1'h0}};
          If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd <=
            Ib398240cd12e68fb5b3ad4842123a4a16f27cfcae3db8bf1f38de24b82e272aa +
            I7e3620302652666ddabcd16531a36e7af51722c39bffc4224f256a34ca33109c +
            I29e9674dcb3b06489c5f9017b95878c6a75503e1dc4e2ba4c9c6a7a7cd74d885 +
            I7e26d67803410d5079a43dbf6053aee09ff9b0242133282679c3beffd05aae02 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362 <=
            I9b494d3414d329e4419da30566795e7b36627870c521c463cefbeb7b48196d3c +
            I3390b463514e772ff0afe74698bc4850014fbe363d105ce3d0e8810706977682 +
            I49a96e94f51c41ba36bb7a8d466771682602e2dbd6f65e13d7e858a60b554f3b +
            I685960b47e49f3ff64eca0e1f26387605e48d325d533550beca6bd6d0f3abbd3 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c <=
            I29d04420073229582b38d6b3f7d9d638351e92073269d5528b09b080e5fd5670 +
            If07308cb71758beb15e4a33e3770aba8021bd5572128b9bbc1c8db48e7f807b4 +
            I4e556f27c558f3d1f76d2ed4a3f0b1a68d74e5c0ce6370b9eec599e7f76f8bbf +
            Icf75218ad23cd1505d2d69d09c0305642a8be48b8a3b7aca4aa4d01a564ddebf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7 <=
            Ia55512c30a26e336794d389f3700b9153cea83619467b731571ba72a3a9374bf +
            Ic46278073f42d4eba79499cd6293cfcb33a74310e7b2ed4bff06f5cc63dc9ebd +
            Ife11a6b34a661bffcf9f0147459d2f5a23d6c5460c59142668ee0f0506755225 +
            Ic9adc8e66938cafc1f6974ab9e2fd71a29bcd6520e6fca93ce7bab4815494ed6 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13 <=
            I0421a9a7aa72d6f574071ffb4c65878f997e6dc2b605f0d8b351358b08c47ce3 +
            Ia84ec437292f1ad3e702b4fa896a4f545cab7253574d294243af0c1e7de47155 +
            Ifc38f7d8250994e5e62716048122eabe81722a32478caab729cfb06aacfc09c2 +
            I4f8e5bee14ab1e584593fc15140a36cf071f2949f1bc86fc3fb7dbfdeea7343c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Id6e462224a7c7f18670d48e3a7c6d35465875f9638395e7dd87b3c494985d418 <=
            I6efd033a5e005d772ae427cab43bfeacb72354d6905822aaf8d484125615d0f5 +
            Ia6058d7a3749f21a827ae6a0f4e792d6cd62ab37d668d607861bdf3985489d97 +
            Idbadcb95f603dca2fe62a931973c10429cefef4d6cad0b8e46cf34b2f7c7907b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2c0782e7324e49c90f18114dc327f50948f9bf80b906f202a50b101832a88baf <=
            I73c8c2e52e23d992ea9758a361fb9550f0ac7f08bb93b6b26c6fab3b234720a6 +
            I3a8f6218aa06df768133a9b95140db0cdd600a5d1a04a2004479693cecd87571 +
            I9f94e32610a6e83f5ca5d8eb0ad81277c7226ae8ffa7f1e734959a614bf1edd1 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I3d8ccc88024eed4b5d118a6c3b8c06553fcfc8645a8569278e7e7e8d3b41597a <=
            Iedb10f981e08498950a50589d8c2fd5dbff191f233da39d5819ddf2dc5172651 +
            Icf3a16773d04781aa96eb511825cc59c609fc887b464a86c7839c57ddbba37db +
            Ie023df7145a8643ec413fd62bad9e4dafc719f7c882ae969eaccbce255ca7748 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ice2f6ae40746fa0bd1c5b2db1aa0bac608899f3ec311d6e8459e126e446f7947 <=
            Ic24e91afb654a0ee04d27daccc66b42d5e001a5962acd08aa73c3e962e1f2c88 +
            I4408d142165f7f5bcee86e820e4ce79b4ecfe2134d8e50809080e0c27e4e2df9 +
            I3a210f2cb408bb61efba033b0ea8f1cda9a3341500248e1443840c24dfe04cea +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec <=
            Icf6cba7551eee2b4d2b53263af6fc190558f5b29af52c060adf5bc9116d56341 +
            I5aff0a6c62deaff6e9d15280ae8c3cc326ae7f9ea6959dfa41a92c770b592cce +
            I6853348c8635a69100a45e6b2b255d6111daca84f2eb28629edd64f8c36f014c +
            Ifd9d392bdf654a9146eebb9a670b75f4d74807786708350ceef7c79d54805ccc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8 <=
            I9df56fb9c7b812f3ca5949962100efeb5889d69ff60754cb4eb3e0dd18376d45 +
            I6c8cd97a5a950e00f0b9892a96d99ad1e5bae6c2db215bbb532060b753233aff +
            Idd51d2eb571b7a35413e786a8a9437a5ef34a13b84d269e29c3319a4bb7531de +
            I3cf51d0ae95d4e3f7d0809785f84c5d25153742e5dd0d370235828d4f9c0d1cf +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421 <=
            I5cbb1dce1049c737c8e052dd6b84121d353e3ee02202bcb8e5fa27261029c96d +
            I20a501f960ccd425135a3fcb8e667d68940a5950d939bca37d107d479984c038 +
            I5c29250eb53f0eefc2332419b6c8e82f97741659657c08af97f8443954a5385f +
            I4fc7c4344699ed94536cb79d86f697e9da22498a2938b10360763aa9bad9da33 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e <=
            I8d463b693ea969ef3023c411c0c9a1fbc49f81d348282c031b963bd8ce0527a3 +
            Iabd5561747d288862c0b289a28572fb5b0159a3fff7f79c59bf60f1612ec1e3f +
            I4e6e6be5d9a7a85cc07a42c3a252e38fad4229a40bd68bec6728e7efa85984be +
            If7b4cbde972a67fae839c5bc9ddfd64dc244041f6dd60f95c5329105ae08e460 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf <=
            I60b41ade4579462091cc59f1faf9f78f236a3bef12f893facebdf8e6b00096e7 +
            Id73bbd3c91f1e5fe13f11e8849f77aad2ddaa35d1399140ceb5e133da8e11227 +
            I8a3b07f660ad94b304ffecabf47d3378d3ea73b1deccd771fd1982cec9f23e39 +
            Icf608ba43019dffad0c708d49076088f2a4b5e126e76b3b2fefa5a0f1edeac7b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2 <=
            I8060bc4cf825f705f2218152b6a7a8600692076ba01123cae35feec231f128dc +
            I47b18bf83ed7f7e8a2c69814aafa41a66b6838a5a997d036c634f488f1c584f1 +
            I55d6bfb606269d9d01dc348f732caf9cfdc7042c845744b7a25c0a74d0afefbe +
            I0a5867bf6971ed11db3a6dc9af8cb356352990bbc3032878e82b6cb2ca8c402b +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987 <=
            I8090d844610f0d62cc25a9c72c2d76d9d6783a067de9c9ea9d5a1f5c48744c70 +
            I79d13cc47977ecb1fb0ca304be8c225a427063b4328cea4c4a227521a1f26018 +
            Ic3f066b6b8dc09e89e9796c2b739b37e64af709758029ee21800f9fdf02c533d +
            I56253c88487a75fb5f830a66c0dd3172ff25795a2509eaf5367fe045f9e12b61 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3 <=
            I799968e729d7842ce09a838203458d89b96fe9d2d7a5de0cbac32eefbf834898 +
            I02962ee90b42f9b95262049bd2dcb7da2f43333787a578d5f5721681773db287 +
            Ib36374f40465c181d1b8d65f23001a10ffaa250f0fd89077848e6a49a19c56dd +
            I199abcfe7a0dfbaa58ab1dbbb16223bd434b4ce5ed3a65633d506d668aa76f8c +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96 <=
            Ib1101385e86160606eeb12ff49ee86ca465f227b19c9bcad4811c6a0183c0ddc +
            I44445d003eed631dd6933d4ade176469fe9a4ef0b21b0ee20067b5aae73704d8 +
            I7c843a280d8a673e3c59a22f8bfbd5860c3284b189ffa281759aa44233eee225 +
            I2ff52a8e46c22b626ca488ae87c88360d413ad08dfaa6701fe7b237d42c2cbe7 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d <=
            I52cf6523f0dd5f666334b2646768fe4499c699c8f6b27ec32ae325cc0981a515 +
            I289b4317d3472843dd49dc75a39395f8c39b9fc0c70000205510d08404d824a3 +
            I5eef24c8de2049e0e8bdd49346b6be22708a135d56c096907e50ecfbf3affdea +
            Ide088b881c7dabf6e2fab61eb4e5db3ea3750d7b72eb26cb79877bc23429efbe +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a <=
            I3e5c11a25b8726c787dd0ffc08e93b671baf84832d9413eb7031a6fc17e8ad76 +
            I2e063205340c315025edf32a4ba91e5f7cd39f37fc5800906a3862780cdf7d9a +
            I29141cb56b9f52d74c42d689b180cfcfe7daf23ce573c1f4eaf21525370e5376 +
            I5df56a6a00d4d8ca1c6b1a79e5f0e674482cb9541d86dd49c2ac361d86dcea1a +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df <=
            Ic2bb8293812351030940ea0e0a882994714d60a4963e82e2291f6f2d386fce8e +
            Ide8930fe855e6fb7dd5b689395a121a16f491421d448454c9c021f62753732c0 +
            I405b2f517ad52ec3c94eb9d1d695f6fb9700fbd32fb49fca23588911b5dd0ef5 +
            I16b3b3cdfef91e9cd5ab763bbcbe2188e61f45183118f5c735eff60965fe4138 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481 <=
            Ib4d2bee91a2ab56208d3d1f484e63f085a162ab9d482690dd3c5891a2a34d808 +
            Ia4205a1d01cb014ebf8e1d539dbe1c7270bf9bfa8eb7920b136417bdfb9f498e +
            I0bafe9c7cb10e6696f6b6dafb74a2113145f7ef1cb70496d068a61ba1de1bea1 +
            I78e49a2727c2f25a14e0f8937e6241f54246c8f42a643dc569f0249384909fb1 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0 <=
            I6822ca486e86051ea654b41b63bfefc12a2218ec87a88d8b5acc3e3c8a604c94 +
            If6fe8b42d897a8c92c628edac7869deee179622fa52fa779f2d9a0279791afc0 +
            I5b2b2323ba78f198e4c86b284772fed82ae708af1da14bfdf215a7b34f811204 +
            I6563fc7a6bd595720441778baa975487126f50343c92ccba99218e274cf40336 +
            {MAX_SUM_WDTH_LONG{1'h0}};
          I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219 <=
            I01a734e70411ca4d260541915dfb0aa0eccbb88be6043a4a46e412d3b9f1e778 +
            Ice95c4df972e8e6a31901269a2d291a70fe4e8dd1d86ea5ded5a16cb1c169890 +
            I4a55baee8cbea583890824bd3ab4c4391b9d44203332575c030077c6e0e9f862 +
            Idc94a4d308c2e301c3d3524f1e20817f9b666827f340874b5adc763970f2efdc +
            {MAX_SUM_WDTH_LONG{1'h0}};
          Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884 <=
            I93f4f945a6dfc45c0a002e0bd9251f56c68570c71e862e222a853f8855fb1165 +
            Ie28b77da5cb0eae41811ec7dbc5f86111d64b794121eda9f2f0515324579f844 +
            Iab63efeaac16bfc91c71a1a0819747c4576111221b2e355300a6e02adddb1aad +
            I3167835472a3c4db7f1b7fbc1895c44e547122e9ad273066e6bdd43bccde11cb +
            {MAX_SUM_WDTH_LONG{1'h0}};
       end
   end







always_comb begin

            Iea34a791d9561118f20388c1982e96791b9c45c8d09efe2e56ce981faa134d13 = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~I435bc44b4b8aac5fe9ba3c30a74d51a42250154c16d5750e075057d1743ffd69 + 1;
            Idb963323153058965c1bb1f6793ee1ed532b856329d971179c54c8172ba1b677 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iea34a791d9561118f20388c1982e96791b9c45c8d09efe2e56ce981faa134d13);
            I893355bf7ee2fbac8f9873385982e6b24128db3c9934e37db7bb8b576a4ac41e    = Idb963323153058965c1bb1f6793ee1ed532b856329d971179c54c8172ba1b677;

            I4c8eece46c2e28444c6f5c37e2e5554529d6939601f8ebc810fa90d8649ed6ee = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~Idf3bd173aa5e956e898d5800f3317a1ef71e334901db42b94f9c6aa41c87c2b8 + 1;
            I623f2b3e99120e8f406c94a41831d851401dfcedfea86f4b34e5ee38b1273b14 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4c8eece46c2e28444c6f5c37e2e5554529d6939601f8ebc810fa90d8649ed6ee);
            Ic1d44b04503cdaccd5821f80e822659de6f6e305c3206e603ef6e23dd3dad3ce    = I623f2b3e99120e8f406c94a41831d851401dfcedfea86f4b34e5ee38b1273b14;

            Ifac89ff7eb9686dcc27ac30cf29859815ca420f6432a51b6f402333f0683a4ee = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~I04257aade4809f3b60c5cd618c5a29008d1b3d7041330bd5c8db7df720da3694 + 1;
            I6e72afb03410a9a976620d722e3b11b93681ed53351a88a8fa3590f65bc2843c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifac89ff7eb9686dcc27ac30cf29859815ca420f6432a51b6f402333f0683a4ee);
            Ia02e90fa0c6b93819416a3059cf6adaaee9c396532e724c47648f414a16679b6    = I6e72afb03410a9a976620d722e3b11b93681ed53351a88a8fa3590f65bc2843c;

            Iddab3676c92e4641120c33849987a24c0d6ce40830d17459f0535c40cc1bbce5 = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~I0e7725af7e163a3f4ee8bf63bcb825b6d62f4b9260a7c68d0beeabf35eea9391 + 1;
            I8bade7cf8bdd5128caf2415690cff8ade1815c1a93e3d7519333c170fecd364b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iddab3676c92e4641120c33849987a24c0d6ce40830d17459f0535c40cc1bbce5);
            I43f540ed8151f48307326f27534afca5105989e179c37e992cc8516996b10bd8    = I8bade7cf8bdd5128caf2415690cff8ade1815c1a93e3d7519333c170fecd364b;

            I0136c7d988171747d52abfedc779c36c470e40bd8043ae469b0c1beea8a077ee = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~Ia718f1fe0157bb564650d817f5ea7960bd0698409dd04d9b31d54c95a3f90318 + 1;
            I1649cd92dddb73a78816076a829f1c12fb8877cae9ebd080a61259a1d2709c8a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0136c7d988171747d52abfedc779c36c470e40bd8043ae469b0c1beea8a077ee);
            I3d7d9699881b5d4d42cc19d1489f8116cf6f3eef7781b1fdc8cdedda72233a32    = I1649cd92dddb73a78816076a829f1c12fb8877cae9ebd080a61259a1d2709c8a;

            Id1218ca0034b49373a64117899424a661aa27c96a30d3ade1da1893fc2761be3 = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~If0025a7dfd37802d1a1fb43d82ff871c2867504735093f0ffaa8b0d85fcd4d1e + 1;
            I2fd0a82f26ad0db034e9db0a2904a499de0ae72c5d12f6263aec7a213bf72335 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id1218ca0034b49373a64117899424a661aa27c96a30d3ade1da1893fc2761be3);
            I1b0a3f720c3ed13e66b1c568162495031330a4369a4d0ddf65848c307e1d56e6    = I2fd0a82f26ad0db034e9db0a2904a499de0ae72c5d12f6263aec7a213bf72335;

            I3e76241b601228fc46605a51baba2f1651b23918015bd484399022d97f09bd92 = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~I35ddc6b67ba559d53bf4b297c2cfd82bcc814a88095ccdf7d6f22fb59113ae98 + 1;
            I45c3eb9c92ff10381f7483843440f1f44e1bceac56ddee98e6bd46c1bd77a1e4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3e76241b601228fc46605a51baba2f1651b23918015bd484399022d97f09bd92);
            I1927b4579e43362f62245cc1904e0deea9705e4427e3bbaeece21a3e36820df6    = I45c3eb9c92ff10381f7483843440f1f44e1bceac56ddee98e6bd46c1bd77a1e4;

            Iced807c14e21b11607cb94ee75e9f432fdda810c34b30a39aef1e50f8ab0e30e = I7239bca55f4296e1befdd8cafa455f8cc6b8a101e498f12fa9a2b9027f8f9d94 + ~I8be8cfdcda8c42fc83b767d9cdd6af256d434d307b8e324bd533b5b016383bfc + 1;
            I0a47b8dba409dae870aa2446c4c554596287cb31f07039a3c01ae78038ffcad9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iced807c14e21b11607cb94ee75e9f432fdda810c34b30a39aef1e50f8ab0e30e);
            Ia341cb94dc5268759917bc49586f20130d999dbbdcd5f1b34e576770d6d063bb    = I0a47b8dba409dae870aa2446c4c554596287cb31f07039a3c01ae78038ffcad9;

            I5ec4520bbe75dff595380b5e3dbc662e1e5193efc9e5b282d68a1bf00585f9c1 = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~Id60b432b19836d2e0919dc2e0201d162d7446434080aff7165fb949aba097f7b + 1;
            I24e4f15f94203d5d70544e5f8b146fcdb89e835acfb8937067299f0b440f7a34 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5ec4520bbe75dff595380b5e3dbc662e1e5193efc9e5b282d68a1bf00585f9c1);
            I34d68a357aa2b44cf3a3b08384498af0e4cc195b0c725a67769d62e36877cb7f    = I24e4f15f94203d5d70544e5f8b146fcdb89e835acfb8937067299f0b440f7a34;

            I107c1cc34b3e7fe3f69400b3e6f18745b97d257839df7315d1f12f3cb9256812 = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~Icb9b19c9fb878af708bd3b433b656104d0f1ae64cb5d5a3f8dfbac08da1fdec6 + 1;
            I32519f336568f17bae9f4135fd77eefd67f37ef3c5b6b624521209fc8a69ecdb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I107c1cc34b3e7fe3f69400b3e6f18745b97d257839df7315d1f12f3cb9256812);
            I48a2995df1784de9dc4a3b951d711905f920ed0b9fc0e20ee48f8838a3ba6502    = I32519f336568f17bae9f4135fd77eefd67f37ef3c5b6b624521209fc8a69ecdb;

            If0a186df3c3fa86b38c53f061c5f78277ae3d14992d047cc5594125a73b50dd6 = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~I4bfb42a957ed14280a129921d4d635017b23dab77b121f51abcc5e738114e446 + 1;
            Id6f531c71e2af56ad8f4d452827d89b82d866570bface8425648576edf2dc62f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If0a186df3c3fa86b38c53f061c5f78277ae3d14992d047cc5594125a73b50dd6);
            I45e3ffea730c76c713d1e61276b644a026af54458af4d3894e44c4416f9e4867    = Id6f531c71e2af56ad8f4d452827d89b82d866570bface8425648576edf2dc62f;

            I16f0af67f0951998267a540be535b5431ed5e6ffd14355109089885e42fc7e38 = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~I1ee3ce036ac0c878003d846cdc3fa9f6b5854855789ea575f0005a9c9937c58a + 1;
            I37d72f048ee656b44e4e465e7325741ce519f38a7c033cd596a312d8e12be42b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I16f0af67f0951998267a540be535b5431ed5e6ffd14355109089885e42fc7e38);
            I573b8edf32c67a0863b9e9ecb44ce7154a48ec67472c04821ffcb202bf3b28e4    = I37d72f048ee656b44e4e465e7325741ce519f38a7c033cd596a312d8e12be42b;

            I25c23909ef7300400c6ca2484a36d95fdd5765d0ab9f816f2b7eae40b2896405 = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~I706a44814e015449aad217d9bd9e0056813b075d8e622aaec4dc08a3518cc0e5 + 1;
            Ie51bbbbf8e9ea4467e2c172d3855c3c783c8bc93166f414044020a5f7f45e7c8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I25c23909ef7300400c6ca2484a36d95fdd5765d0ab9f816f2b7eae40b2896405);
            Ic2544a607bb965371402190fd2fe4afbd85977e8360b5f0091a6f11f885909c8    = Ie51bbbbf8e9ea4467e2c172d3855c3c783c8bc93166f414044020a5f7f45e7c8;

            I29c0576bd0d8df0a78aee42f63a6007df95d1b2cabb7424d322627654b6a0bfe = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~I804112f16593c6ce81f6459599203b07642485939c898d78e113353659a62a68 + 1;
            Id851fac0751063b14367885b08e771c57d9000f29e0e529be1106e6accfe4eb1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I29c0576bd0d8df0a78aee42f63a6007df95d1b2cabb7424d322627654b6a0bfe);
            I1a641c18ed7edafaa7d5877ae724860b1d54fa6e6890510d1c7febf66944bc55    = Id851fac0751063b14367885b08e771c57d9000f29e0e529be1106e6accfe4eb1;

            I06f14700638e4bccddacf4896cd90e26b33f1388f0a21678bc35a81fb8973e02 = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~I95b68240d25deb08902e18ba5fc3ed7af68c0a6ae8e629edcf59930ed55c22ce + 1;
            I71ea9226d39bea8f66f1c13855318e475eca4a45fbcdfecb5b5bea94e9895019 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I06f14700638e4bccddacf4896cd90e26b33f1388f0a21678bc35a81fb8973e02);
            I7301f67cfc0739e38aae8830e112df2193600d9581476251265730522284b6b5    = I71ea9226d39bea8f66f1c13855318e475eca4a45fbcdfecb5b5bea94e9895019;

            I07a85d69a58e9ae8356b7758dc0c989aa6bcd71b408c3c7770d0e646bdd5ef2d = Ibfd9f5e041a831de3b7d7a5dcc5b194397e724eb6171e70d4b9dffb5308dc75e + ~Iaae1f131bd6bb3b2fd8e363e97f6f9e680c7ed035a086cdf2bef5cb7e023c6d5 + 1;
            I4211635a82c1f604dfe16daddc0995754675f3d3059ad427ba374cea6f9e36fd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I07a85d69a58e9ae8356b7758dc0c989aa6bcd71b408c3c7770d0e646bdd5ef2d);
            I41ff59a42cce4bf7225d8f9296ec89aab75a0ec2dc10f0c341c696fc2461ce3a    = I4211635a82c1f604dfe16daddc0995754675f3d3059ad427ba374cea6f9e36fd;

            I9dcc9ad0f4591fe0ea9c5196fb457aaab567f5be24fff2b29cf4e61567811938 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~I2e17b8ef0d25ba5beb474e7007ce1fe5f99f6f7cbf24e5241761880a551f3c12 + 1;
            I41e027c49a3c7e7075a937c21a58688cd46356ff9a8ecfd497cc216b1d8df456 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9dcc9ad0f4591fe0ea9c5196fb457aaab567f5be24fff2b29cf4e61567811938);
            I799ec6460c042feab5ece45c8877d0614bfea4ebd97b427e1bd00aaba217c1c9    = I41e027c49a3c7e7075a937c21a58688cd46356ff9a8ecfd497cc216b1d8df456;

            I23c501712a70f0ada92c78d2c0704b55e90588bfea60dd5c3d6dbb0ba70ed009 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~Ie515c89eac4b602d36f70f52a3fd62fee155da2eafac9c1b14bf1917b62bab44 + 1;
            Ic090c90fe7246cfc964e807e465274744fde1c059c1a86c193a553def4295df6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I23c501712a70f0ada92c78d2c0704b55e90588bfea60dd5c3d6dbb0ba70ed009);
            Ibf5e207961c05c6ea8ee1cc657aa7bf8a0fd7827e4e550b65cb9cc20925f7536    = Ic090c90fe7246cfc964e807e465274744fde1c059c1a86c193a553def4295df6;

            I8cc4346951815e7dd3951d1975e1d4529332c497689815c86cff1a2e6bd98872 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~I7da5ecb7bb8a413a5c6c51f0aff1921be97bb5df5d56f6648c27ee4196fa93db + 1;
            I523b27aea266bed319f1eeb7acb39554b6d1129e3c850647d3d0a5f6b4ee87cc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8cc4346951815e7dd3951d1975e1d4529332c497689815c86cff1a2e6bd98872);
            I1ce1761a25063d6ca639d1aa9094a30899744186121a71229f255eaf3542b80a    = I523b27aea266bed319f1eeb7acb39554b6d1129e3c850647d3d0a5f6b4ee87cc;

            Ifb944e4f518bc9bee1423b4c08427b203b24f130be8430fd7afb83bef7ba0d2d = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~I83ded8cd9258de3ae8deb907ae3b813cc228b189df92f42c55a4b0eaf411c106 + 1;
            If3585e76d77927b87fa2b357b5f3755404054e391f29839ba9c3a29c0a1084f4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifb944e4f518bc9bee1423b4c08427b203b24f130be8430fd7afb83bef7ba0d2d);
            Ifa331e88bb390c67efa83efdb978b28023c3f4a74750928415242eff2a75326a    = If3585e76d77927b87fa2b357b5f3755404054e391f29839ba9c3a29c0a1084f4;

            Ifcb9110b05d9709662dcd3a0c985290be9f283f2b76d0a82a60b59fdfae1f116 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~I23d075a3ac353b3deca0a572e9cbec9b1ae24ffc7f134b36c6f938d949bdcb1e + 1;
            Icdb198ad2d4b3ffc14486474c17026ab6c9129e1783a62dfb7046874dc639667 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifcb9110b05d9709662dcd3a0c985290be9f283f2b76d0a82a60b59fdfae1f116);
            I7e5dd2b4a968c805518feeef59ac29c86d9c06c30446f8966bff4b169c65962a    = Icdb198ad2d4b3ffc14486474c17026ab6c9129e1783a62dfb7046874dc639667;

            I4359ce5cccb720df3276f0771c774342c0e7ee09f4e356283023be0a60cd1115 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~Ia61e8ceb90369d4ed8ed86b9cdf7d4e89056cf4fca5c7e223bdd7b2c5656ac9d + 1;
            Ifd4918d774147592104adca1c7b4abe2c20a82553bd5cdbae652d80335fb933a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4359ce5cccb720df3276f0771c774342c0e7ee09f4e356283023be0a60cd1115);
            I9663885f1f636653b6649709c8859bdf9e407c18311f63a0e6677f6671926884    = Ifd4918d774147592104adca1c7b4abe2c20a82553bd5cdbae652d80335fb933a;

            Iac34667e98a93c9bb269f6dbe69d4148df3a55d9ea25098e7630a36b5ab58138 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~I7bbabd42e7ee42c653f61b4bbd72ed2b076dec2c89baaec2b4589bd55b92fa6a + 1;
            Ic935f15a1c1aa2ee20c06cccdc61d9b18929a70e43e44123bbc51e64bf29e1fe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iac34667e98a93c9bb269f6dbe69d4148df3a55d9ea25098e7630a36b5ab58138);
            I9e8163c831756fc1d31bf9bb6e966a5c58738673504240801b73891e606845ac    = Ic935f15a1c1aa2ee20c06cccdc61d9b18929a70e43e44123bbc51e64bf29e1fe;

            I0c29df9d670f78350175d3c013388fbf48c167f3cfc7576f8d56186e227ee2f1 = Icbe34503610ebbe63344491d0ef8f8bc70117e7d4b305f3894920dda30d9b6e1 + ~I0e9e95de14abaad3f4dee2c74242d09121b496fc60f22dd3513b90860e7d03ab + 1;
            Iaaa7217330cfc4c43630903983e580f1ae9eff2fa7200e236b2055614a50531c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0c29df9d670f78350175d3c013388fbf48c167f3cfc7576f8d56186e227ee2f1);
            I211a4aa442cd695ebef8bfdd8734fca64e796eec6eaeae0f7c1c306d89ac50ad    = Iaaa7217330cfc4c43630903983e580f1ae9eff2fa7200e236b2055614a50531c;

            I3b58ebce4a4f16f7271ba1ae7dac9dc9977abd0c90030d9aba39ce0c5d604478 = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~I7bd679f7d7da9dc0742c725247978f1c14611083c7de896c4c2de108c6766fb9 + 1;
            I76857068f374b6f47eda0c4192e95879ea55667a3d96b78003079f89c096843e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3b58ebce4a4f16f7271ba1ae7dac9dc9977abd0c90030d9aba39ce0c5d604478);
            I2e3ac37a60fed64971c398ea5f48490f1a8ba9c0fe63583d4996ef4884aa0eea    = I76857068f374b6f47eda0c4192e95879ea55667a3d96b78003079f89c096843e;

            Ie0a8e687a253c1e072e5d299c180b344586ed28837bbf2b20a2a737dfbb904ce = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~Ib5d526172ae46c2a06c11e15361cb13141d0ba754320f60ce6bcd97a9e495221 + 1;
            Ife34f6a36501f7796b3321efdacf37a75e6cb15cc2276751fd20794654b3c515 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie0a8e687a253c1e072e5d299c180b344586ed28837bbf2b20a2a737dfbb904ce);
            I71f710555439b202404f08c784a66fffed0e12c7dad92ced1b83a6f28245a512    = Ife34f6a36501f7796b3321efdacf37a75e6cb15cc2276751fd20794654b3c515;

            I857c867fb70f76bc0c7d09b8c34d62fe9d558eaf96766b58b776793692b63497 = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~I6b499c648458a2ed0cf0b27d81aeb706a260c5615a8def0ae89a1a44693061c5 + 1;
            Ic269a154a2e6550cdc5270948790b9962936b7fe59e88379d1fb543fd7f9b8f4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I857c867fb70f76bc0c7d09b8c34d62fe9d558eaf96766b58b776793692b63497);
            I458d537d6f291b854051834fc85511253dbd0054f1be7bde7ac2696c4e4424ca    = Ic269a154a2e6550cdc5270948790b9962936b7fe59e88379d1fb543fd7f9b8f4;

            I3c98ae8ef287ba03079f7fd14ee83b588b02cf1b02e362e12737c93f35031230 = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~Iba5fd100311e883873db0c3474169654308059bc4c43d52479a4515fa85e8900 + 1;
            Ieb1ef347bc6ea6aaed4c4763221f318e5b5db3997be4a4d107e338cc37e3a4bb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3c98ae8ef287ba03079f7fd14ee83b588b02cf1b02e362e12737c93f35031230);
            I3e27399b8d9e65418758d9dca1b1cfbcb4d908000611b218f4ad2097da556a51    = Ieb1ef347bc6ea6aaed4c4763221f318e5b5db3997be4a4d107e338cc37e3a4bb;

            Iaea6828ee218d24373cfb8449c584b5806a1a815d7ab34c2a39d76dc3186ca3b = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~Ibdb4937356d2b1cd2091a695635cc7c69b694f775f4c4e8680ea49df1ea6722d + 1;
            I9d8215327a40c9b967e1a5dc8c9e9c390c37bf87f96114a7d81cd08285223c43 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaea6828ee218d24373cfb8449c584b5806a1a815d7ab34c2a39d76dc3186ca3b);
            I38ef2b3fde182cebc6e8265c6e99d08e21e28d55b2eb1b7a161f13e385ac5b72    = I9d8215327a40c9b967e1a5dc8c9e9c390c37bf87f96114a7d81cd08285223c43;

            Ic34d5eef3a8c9a0ff524b6ca5d233209869368afe0266bfa94c6d159c3b4b97d = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~I238b01744b520f8759a7e466290a15b15b96fc95b4b8a14afacbedb1657f7069 + 1;
            Id71a454e9889c6cf7e01d39d50bde9e8bc5850b88ccda4c91eb8266ef7e5a695 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic34d5eef3a8c9a0ff524b6ca5d233209869368afe0266bfa94c6d159c3b4b97d);
            I0f2d9a8f6ab682ae8c5fb31b30d5c11be65370398f373fda27a64bf6d718193c    = Id71a454e9889c6cf7e01d39d50bde9e8bc5850b88ccda4c91eb8266ef7e5a695;

            I92306fea80ed98e3391ee19be59721f0ddf93aff9c5c85a1c03942ab1ddc0b7b = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~I4909110fd7213171cbddcd3545ba2a0d3a135e723189edadc7c64599fd2f1f53 + 1;
            Ib5228b88950d45370aa8a132d3824bd69b574875b1bd9d3783780b87edbc3ced = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I92306fea80ed98e3391ee19be59721f0ddf93aff9c5c85a1c03942ab1ddc0b7b);
            Ie504e487c65a8cf270fcb907ff7a6f204c5afe50af53c0b0279719522b595c19    = Ib5228b88950d45370aa8a132d3824bd69b574875b1bd9d3783780b87edbc3ced;

            If38b0396ad61a4a69acd171a8474d2270c09dc3cd74273589ce39f3cf9c2d9c6 = I0843b40b0650450cc5656d30e0afb90a109189dabf6379f0dabd39016115d0dc + ~I929870fcfce11dff715cf2210ad4a4c30db9af500a8d380153f38f0ea2b7c2b3 + 1;
            I2c860739a98a8e6052efa8701d70df89f34952d6249f7266956ad0a6d6701159 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If38b0396ad61a4a69acd171a8474d2270c09dc3cd74273589ce39f3cf9c2d9c6);
            I7306fa7f8f192749aacf00bcfc3ee6266ad06e373f4075503bf8c7daa963f7b6    = I2c860739a98a8e6052efa8701d70df89f34952d6249f7266956ad0a6d6701159;

            I2aa525f826749dfac72e0a870919582cf43e69ce68dd68555201ca204fad6ee3 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~I7cc2cdc76a638cf4fabcdbd60142d7e4fa11f11486c85b7add7d4f9ba16042c5 + 1;
            I250cee6e4a22b9f9fe50b6acc67a25365520ec326130a11c9c68cce437e6f56f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2aa525f826749dfac72e0a870919582cf43e69ce68dd68555201ca204fad6ee3);
            Ica9704300b0989fb0bb8dd9ddc1807a4906458c6f7f487fb7d7e214e31458eb8    = I250cee6e4a22b9f9fe50b6acc67a25365520ec326130a11c9c68cce437e6f56f;

            I8e300db9fc7aee834809aaf20ac393fc3d046ffe391d61effac8eb11f7daa1c3 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~I9a798d59823ac9a032d0daa203a7bb153e483bbe4fc47083c1d7e4a65e400156 + 1;
            I805133cb6a397bf027d1985ca36380b66ae7d0b33ca30987f825dba8d803488d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8e300db9fc7aee834809aaf20ac393fc3d046ffe391d61effac8eb11f7daa1c3);
            Ic8e52a8db0d0cf4d90f46c2d5b5871d31db974cbd84b5e68f4d872ccb6fb9cf5    = I805133cb6a397bf027d1985ca36380b66ae7d0b33ca30987f825dba8d803488d;

            I7f4e6a672481e296d10f94ea345bbe9babcdadc2e3b447be67ed1cb4c5b5b010 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~If307a1ee8e5164bac03971d07c03c3c0440857c7cc29df11a751b3bef9bb1516 + 1;
            I71c2e463b98044653ab94090116d3d5093fcaaf7ac48bbe2f5b2b26980af991c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7f4e6a672481e296d10f94ea345bbe9babcdadc2e3b447be67ed1cb4c5b5b010);
            I59ef74fe764da43c107f5eb1c48cc198be3cfce3b3c55e0eac3efe7c9af888a0    = I71c2e463b98044653ab94090116d3d5093fcaaf7ac48bbe2f5b2b26980af991c;

            Id1d212084a29e275b0e589f056235a0f87097cb4fe96989ee3e2e8b44b8d14c3 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~Iefca48dd9d0f3c717b0a3b081894e93ac451ed275f3cfa7aed675f58327a2d02 + 1;
            If85b088f394e161ace940e64c404069e394099027a64365e447bebea842a0781 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id1d212084a29e275b0e589f056235a0f87097cb4fe96989ee3e2e8b44b8d14c3);
            Ib33fa9a97b26fc69be1d69ad97dcc345c1701bd9ca2fb0922d724237bd2cf8cd    = If85b088f394e161ace940e64c404069e394099027a64365e447bebea842a0781;

            I0df196e9a75907dc29b66b17b63677adc1d35b6b543dfb5ab01f7beedef65a95 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~I18e5d7f94022748f9a5645c2b0e385407e0f00d6f9ab28a55982fd36330ce524 + 1;
            I92da904919e10cc11e45847a0102a3b8cc6c52cdc4815d7de7a6c949a2024901 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0df196e9a75907dc29b66b17b63677adc1d35b6b543dfb5ab01f7beedef65a95);
            Ibc1655e6f13d450c6beb85bc81ffd4b765ed49cb361ddcae84e6e635e85513da    = I92da904919e10cc11e45847a0102a3b8cc6c52cdc4815d7de7a6c949a2024901;

            I45edda32704ad01d8fa7f3baa6e5836bc669570d223d634ad149ab4580abd625 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~I727007bc323c90e0c264e5b8688898c0df1bb72c976fbc3513439c14f15b5733 + 1;
            Id3bd78d48b87d258733b0c2d0a166e6921566570e0131a68d8dc65eb28ca4a1c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I45edda32704ad01d8fa7f3baa6e5836bc669570d223d634ad149ab4580abd625);
            I170b2f3df88d573e89dcd7abd2e33192d1e08eb33a333dab67be7795d2371e04    = Id3bd78d48b87d258733b0c2d0a166e6921566570e0131a68d8dc65eb28ca4a1c;

            Ia3e1f15e4a1a4c0522470cf8fb86314da400e3e882c97731468b384e9d84e739 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~I739fb2ce1dc1a27f40af1c53d575108539718f9d60f83de60531d7bb201685ff + 1;
            I3833bf9f2a4fc740f72874fec3b21e205b6fbdaaefca4942cee8751f170d55be = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia3e1f15e4a1a4c0522470cf8fb86314da400e3e882c97731468b384e9d84e739);
            Ia554b8c5dc66b7db32a935b99a2e41aa84c6c13fa944f2de90eed8c1d462d023    = I3833bf9f2a4fc740f72874fec3b21e205b6fbdaaefca4942cee8751f170d55be;

            Ib8ae927e56d694255bb5d70c5a6602b13e582f7ec4b06fad5c0f1c623b9bd64f = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~Id29a54af13b6045a8a43f741c229ff88d4aeeffef29065cb29cffbd861479f7d + 1;
            I62f9a8d7e8821466e48058b064f25fe8420acaf3a00a1eafc36103bdeded51c8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib8ae927e56d694255bb5d70c5a6602b13e582f7ec4b06fad5c0f1c623b9bd64f);
            I60e54e7e8d975cee4bf0823ff91ce212f02e407e9e2064ea4ca882ba4961553f    = I62f9a8d7e8821466e48058b064f25fe8420acaf3a00a1eafc36103bdeded51c8;

            I2956ab41e4cda82864182a110ce8b803793f9e0dbcfccfc439f0e473385d9746 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~I31ef992f17daed0e1947c4d26611e7377d8b3049bb8ae2ffb3d56f3db5f85916 + 1;
            Ifb8ea528ec3a42384215586669a0abeab4982d73d76a71c72e4c5c45ddb937c9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2956ab41e4cda82864182a110ce8b803793f9e0dbcfccfc439f0e473385d9746);
            I4470cc46d92649aa472f4dce99afb05681b554782384542942fb243099cfc6de    = Ifb8ea528ec3a42384215586669a0abeab4982d73d76a71c72e4c5c45ddb937c9;

            Id5cf825b09ae8cc8c7c63eec98a9a37fd15767b0f44364dc17e6abde6293a711 = I00ae7a7de011b32cd6fa30759fe7a98468c6e9da295d642d4b364e24a880b769 + ~If51ca9faad7b057d5a086daeaf1118808bbaf90b484e38571530cc3bb497dee9 + 1;
            Ib9a1b462db35f3d9d512995ddb639c3553c22f5020cc3fe7316a605096d8b8a7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id5cf825b09ae8cc8c7c63eec98a9a37fd15767b0f44364dc17e6abde6293a711);
            I9f258a7197af9b66d573a49b5923adec1c8637c53af4c2073805fa31fef73dfe    = Ib9a1b462db35f3d9d512995ddb639c3553c22f5020cc3fe7316a605096d8b8a7;

            I7d405f7f9d952c8a7ca9daf1fdf591b1c0108a683ef3084c8bd0a95d7ce42788 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I11abd59187e2db0058526cb1ea58af9061d439139fa151aaa74184499fcfd24d + 1;
            Ie51c190c3c1827c2c707668d10923b176edee9736a17f532e7ed432af0544083 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7d405f7f9d952c8a7ca9daf1fdf591b1c0108a683ef3084c8bd0a95d7ce42788);
            I52497162427ed0e9f305f509a79ddbdd02f12eebc337f57d63a9e477ce556e44    = Ie51c190c3c1827c2c707668d10923b176edee9736a17f532e7ed432af0544083;

            I88d3389ec9d452ba7af534f1a58d6463b08369c185e66a77bfb6604e6d201916 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I91c40ee5121cd738ba7213df9bda6130b101385a28d8a5fef6544c86f6bd1e3d + 1;
            I46ef2ced2e09d9ef212937cb037346d3309bba86efe06537a39a963d9debb65d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I88d3389ec9d452ba7af534f1a58d6463b08369c185e66a77bfb6604e6d201916);
            I7d53fc143b190930a55ef8fcf893ea0b45d87abc54330c08bf4b4d5c67d4cbda    = I46ef2ced2e09d9ef212937cb037346d3309bba86efe06537a39a963d9debb65d;

            I0d869013e0ccbc57f7bd590ccf22dafd343f209d7a547f1d24b105b31815ba18 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I2976810df2af0dd2879fac8afe975126944b2e40a51dc7dd169051bb5086b3de + 1;
            I37b543101174150d8b288848968eb5974a06d0936975538caab590ec97366a1f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0d869013e0ccbc57f7bd590ccf22dafd343f209d7a547f1d24b105b31815ba18);
            I7f819482e0a2454a58a949963a2600e43477da52fcac968f397cade6b69be570    = I37b543101174150d8b288848968eb5974a06d0936975538caab590ec97366a1f;

            I707948c8eb9a0d646b7d61a3b86b807a4e9962d5f81c582212a6bc7fc58e3c0b = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~Ic45f0213074aad63c68cf3fe879ad5b0e70a5977f282822ab582ab88ae7236bb + 1;
            I36fa36e23de34e375c1e39c129c8aa1f63ed250191e4bcc0cddeb9815fc1c717 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I707948c8eb9a0d646b7d61a3b86b807a4e9962d5f81c582212a6bc7fc58e3c0b);
            I551c9d548f30a033083c22bbd3fb8c0ad11c32fbbf66ccc8d0f6b7a177a49b39    = I36fa36e23de34e375c1e39c129c8aa1f63ed250191e4bcc0cddeb9815fc1c717;

            Ib1b8ba2fabf6c4f6336045bd785ae8b52ff275740fc54346295ee42b9ba530a1 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I3599299f7f89ed3c6b11b31caa26e6b30553b9dcc1d5968283085959f822a4c6 + 1;
            I0cb9d359df8b98e0323b9bb85a1efa6ba10fd2478777accabfa9e658d8e02dbf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib1b8ba2fabf6c4f6336045bd785ae8b52ff275740fc54346295ee42b9ba530a1);
            If00a6af912a327873844b41dfbbcb9b7383e07272e5eb09cdf9b4a4a827b4f1f    = I0cb9d359df8b98e0323b9bb85a1efa6ba10fd2478777accabfa9e658d8e02dbf;

            I8fc3cd3e94bb31bff1119828a5ed77af969c8ae0ad80901b9e6303491db001b1 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I2d89506b7ec0311db709c4aba53b749ec1b531bf4bc7867f3866c39a73aada38 + 1;
            Ie53bff4851def180b28f22f53a301b0e7c0e897bd637a0045221b0e969249ddf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8fc3cd3e94bb31bff1119828a5ed77af969c8ae0ad80901b9e6303491db001b1);
            I770b9333cb3aebf6d60d58661bc3282c1fed64de0824268f9f7aaa2dad91efc7    = Ie53bff4851def180b28f22f53a301b0e7c0e897bd637a0045221b0e969249ddf;

            I70a05485fe3663a0704c166ec4819fdd34b5b705623ae6f1c76a783449f04af6 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~Ie3e85438dc476813cea40910227c7d63eb275948fbd481f56cc51656c1bc8b34 + 1;
            I735d477462d8bc4faf83227feb6433daa37d331e95657535b4e8db091cf9b315 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I70a05485fe3663a0704c166ec4819fdd34b5b705623ae6f1c76a783449f04af6);
            I27a121a528b8c373659d1b04c8b5eaf5856b441ddf1b24331855326f31bfc492    = I735d477462d8bc4faf83227feb6433daa37d331e95657535b4e8db091cf9b315;

            Iab0a5fa6bdfbb14163473868e4651dbf1098141c464648018316844fa71bd877 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I24dbfd322139e6a1964e587f89b06274c35617e961a5f61f90c67ee3b20ff208 + 1;
            I9d907af9ccf3e40047d3c7e02550caa8588212f478714ba92e91482893944968 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iab0a5fa6bdfbb14163473868e4651dbf1098141c464648018316844fa71bd877);
            I044870873609a6dc7acef74d59eaea493c553cbcc3eff5b580dfd6a8f176d987    = I9d907af9ccf3e40047d3c7e02550caa8588212f478714ba92e91482893944968;

            If86295d92e67aea78f792b994694f74fef76cca427defd79e2368750b480156c = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~Ic1711dd767cbb72abed2584c5bc27d5422882cb4299da3914c684696eded290d + 1;
            Ia588f9a4cffca8b6d433336ac4fdf52e81a27bdbeed8cf2a5d733183c7aa86f2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If86295d92e67aea78f792b994694f74fef76cca427defd79e2368750b480156c);
            I1db3917cd01f808a2a2f4c78ef1ed3328ca804093065a1cfb9e15ef210bb8c93    = Ia588f9a4cffca8b6d433336ac4fdf52e81a27bdbeed8cf2a5d733183c7aa86f2;

            I7c78ad362cb79bd72205c943398381fa981d5b2e995582c7b16089de4bba9b27 = I67c636b3ff5f49cf428a737b6c3e7faf66e61d2f08f877cba359e21c465f1722 + ~I8e6aa1d0b76cee0ce4862aa5d01ee91caa123335ab19a2150e8c4315c7d958c6 + 1;
            I06e5c848aec73e10515e09f5e32ac2db3c5a972a8084519617121e18c27f4bbb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7c78ad362cb79bd72205c943398381fa981d5b2e995582c7b16089de4bba9b27);
            Idd38249645258d9f8ef1e5cfbda4f15a700ff3b6d78b9c202bfbeca278528f57    = I06e5c848aec73e10515e09f5e32ac2db3c5a972a8084519617121e18c27f4bbb;

            I5a70e23cd0dff70ed6ed5b227d239f56dcd214cbb2fdb0286c2e154f4e450ba4 = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~Ifc131936849b96a3bcc7bed4c38ebe94d51c56feb4e96d25dfbbcc3670568a16 + 1;
            If809ec52b215e06373de8da5e7b6b16db8490684dab7ae07b39bc7440e19f4bc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5a70e23cd0dff70ed6ed5b227d239f56dcd214cbb2fdb0286c2e154f4e450ba4);
            Ie2757ee84c5d0e87b17c22db78eec37478ff53ed9383587a3afa0e3270afde8f    = If809ec52b215e06373de8da5e7b6b16db8490684dab7ae07b39bc7440e19f4bc;

            Ia7ac2e243e12e18eb1233f947496d37da38950a0a2db140cd51b6e3ea075848a = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I89ca3ef99e4b84441ed3cd9f386109125b6da2d23485fc22513b1d8ded87f894 + 1;
            Ifc9e721cab51c6460c44a26b6803f4cbd505fd11afe41341e3ec656fe2698779 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia7ac2e243e12e18eb1233f947496d37da38950a0a2db140cd51b6e3ea075848a);
            I85ce012ac5bad111ae4ab945035baf1b2820c82822f28a7b7c314515345af8a3    = Ifc9e721cab51c6460c44a26b6803f4cbd505fd11afe41341e3ec656fe2698779;

            I2c9e693d898458dc309fab7b6d2492d5b78b53f9c89ef8e7bf3f8038972b2c24 = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I4c871d8c6a677ef8fa6c955524def78e8df6f9f3fdafb141d43db76d4569104d + 1;
            I0b55c5a4fc86bd53678cc688a8577a636d79a0d9b0f515135007234a4a807541 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2c9e693d898458dc309fab7b6d2492d5b78b53f9c89ef8e7bf3f8038972b2c24);
            I89db4b6e1da27586c9fb92f89e492af68c0497029c97adbcdd5e3facac07c213    = I0b55c5a4fc86bd53678cc688a8577a636d79a0d9b0f515135007234a4a807541;

            Iea4dced4cd8775da052c065ef31c3abf4aab1d0b2654d5f7e904bda36ab05ec0 = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I10a223d797492c10ad8f6aac1cbdae83833e701ae6314ed988ac117debc98c33 + 1;
            Ib378ca85da27dec3042e6f79bfea73ae2f099d548d5ea58fd3bf61c2ff85a4bb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iea4dced4cd8775da052c065ef31c3abf4aab1d0b2654d5f7e904bda36ab05ec0);
            I3bdc9359c749bc85fb3a7fc68446c47edf3565e167d9a28caf4bf5010b95a575    = Ib378ca85da27dec3042e6f79bfea73ae2f099d548d5ea58fd3bf61c2ff85a4bb;

            I5a5083c658290744b00a18aaa5fc88ff90eb17aa0c06746715f76592608ace49 = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I95e467521db517b858e59156f95992ddc522a7d038ac6bbe691a91b567cd35af + 1;
            I1bb76da4e4cc33ffa0f6f61ee985779f4f7a02f8e336f7ee969bf4b4d1599fc7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5a5083c658290744b00a18aaa5fc88ff90eb17aa0c06746715f76592608ace49);
            I09a731c0252003cf8c9e4848c2e8ecb6a86e0bf4d76ed8fe028e3a609d639aaa    = I1bb76da4e4cc33ffa0f6f61ee985779f4f7a02f8e336f7ee969bf4b4d1599fc7;

            I5e65da8fb9465ec0e386cc33ac36903a3dee2c59151adc9c83091591a0bf554a = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~Ia9f80db3bd889aa11f43f6aa371715d6aadc7d3aeac0e9519f79b787da6e545c + 1;
            Id1fb2ff888cbc4ad3ddee50de256240ef2be853fbe54f51092a1bfcf26ed4fcf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5e65da8fb9465ec0e386cc33ac36903a3dee2c59151adc9c83091591a0bf554a);
            Iae3ca8fe4281bb23b5ed7e87317e7aea52a130420731529f44179ea0274a58f5    = Id1fb2ff888cbc4ad3ddee50de256240ef2be853fbe54f51092a1bfcf26ed4fcf;

            I1911ec0cf18a635f5d524a57281219443e1eb9eb4cb4f9b5c5f07dae014ead9f = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I0543957798ccd8923b2a5b736175c6888eb71c1466a1e9cc7d7635701e103823 + 1;
            Ia03c4f3191a16f379150692d47660685ffb0b79d91fa4026b8410e2c02219dbb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1911ec0cf18a635f5d524a57281219443e1eb9eb4cb4f9b5c5f07dae014ead9f);
            I38f8f9e2731f858a15a6f2f3a375d0d29634c0da467767e21318213ae7beee7e    = Ia03c4f3191a16f379150692d47660685ffb0b79d91fa4026b8410e2c02219dbb;

            I09c8e5480f9759a5e59d4ef582789a986f66929ee1e1cc030f6f1a716339d4d1 = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~Id8a5ef9ce42d57c3feb442ca091604f1fc51e648a89794ea3fbe4b30537fd286 + 1;
            I44aef1d958b6a776898fe8f0f0a8ebc867154b9d4605421433b66f6832c2be1b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I09c8e5480f9759a5e59d4ef582789a986f66929ee1e1cc030f6f1a716339d4d1);
            I01eae75c6d18bb06d82fd21bc1aaf1cb883bed514f5497fbc433fdc42d217535    = I44aef1d958b6a776898fe8f0f0a8ebc867154b9d4605421433b66f6832c2be1b;

            I29e4efa13123958a82952155cf24212b7f04fe94bf1aa7579617cabcdfd49d03 = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I67874ca15a0723ab01392f527151dd5a60a71a0dd16cbbd572fc50a343c684de + 1;
            I1659da800cada125cbe3b104cf7d512523aa5616f7c9ce70ac7c72fd92403027 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I29e4efa13123958a82952155cf24212b7f04fe94bf1aa7579617cabcdfd49d03);
            Ie5a56b54b520cb4b1b0e5509ed4b3fa804bfc0be8566ed98b455a29b7148d291    = I1659da800cada125cbe3b104cf7d512523aa5616f7c9ce70ac7c72fd92403027;

            I24cce2dccb4540ed239adc5602a5cfb9a2a480bdfa780124b0d05dba8946730a = I12ffd423da118421e4cc1bb1c4706e7c5a5090acc19d6785552b7bb7fe288e3c + ~I2a9f642cd74521fb661e381a3f57eaf539ca18ff62ee2130aa94da51cd13d4c0 + 1;
            I09149397adf0c3b57e577b66b5b3a58bd1396ade0ab7cb174692b182e52141d5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I24cce2dccb4540ed239adc5602a5cfb9a2a480bdfa780124b0d05dba8946730a);
            I0a4b485210baac225fd3f32b36be68140468a6c307f3f91de4416553421e3db5    = I09149397adf0c3b57e577b66b5b3a58bd1396ade0ab7cb174692b182e52141d5;

            Icb9ad5b9e222f215f848ff5fee922a8dc526f16eba35decb2cc80395c848903c = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~I96248ed668211f13555b4a086e7534b958b901242794b9978d673726d56286e0 + 1;
            I15d75a1d3038a54892de000a31379baa7cb9de5538a2823c1e52f64fb061b914 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icb9ad5b9e222f215f848ff5fee922a8dc526f16eba35decb2cc80395c848903c);
            I172389b084abec531bf617713612fa0d8b27b0967bb62a6514aa873f609bb5b0    = I15d75a1d3038a54892de000a31379baa7cb9de5538a2823c1e52f64fb061b914;

            I181f8d112163d3cd54f1842ed88acdee6575a19ff24c4702f463ec4642361196 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~Ied8c84dd66ab8e8fdeb83c6156b8a6f8cbcbee27c41ccdd8c4d199f70ea67e8a + 1;
            I21909db4fda5a886100a19a744a9b172b3d171ccd1dddcb5c47b0d3488a48f6e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I181f8d112163d3cd54f1842ed88acdee6575a19ff24c4702f463ec4642361196);
            Iff3e149eb4ce60c9f28638248c33ab96208976458886b1735785c2dba298121d    = I21909db4fda5a886100a19a744a9b172b3d171ccd1dddcb5c47b0d3488a48f6e;

            I39c3950d86099683961f34448fe235f94e87f5b7067a39abaa69732a48c0ba79 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~I592170f431e8a8e15769fe2e5f3bc43a7c514290149bf9b93a8f3d3a748094a3 + 1;
            I668cba84a2aaea84945a6ebb1a72e6668cebbcec3d78bf88246f3872d78abb2c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I39c3950d86099683961f34448fe235f94e87f5b7067a39abaa69732a48c0ba79);
            I1bc8f647801308e33369cc5f2652781230a588ae772b1e53992f2124c17ad5d9    = I668cba84a2aaea84945a6ebb1a72e6668cebbcec3d78bf88246f3872d78abb2c;

            I456e1a4a9412cedb175a75a2c7b65837b127c5f2478a8bad034592dc7db84079 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~Id8cd2e026867692af509cd433fda0fe6a8b5ccb8ed91bad6530d14172dbf7375 + 1;
            I2bb5bd1737da6b4feec1bbd2245644956d6e825951368ab22e426f1662650a32 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I456e1a4a9412cedb175a75a2c7b65837b127c5f2478a8bad034592dc7db84079);
            I4e3be7e07012df2e0a3bc90dcb0b4756a778cfcf9192e3722191ba8be32e7e14    = I2bb5bd1737da6b4feec1bbd2245644956d6e825951368ab22e426f1662650a32;

            Id5d890ac1e6399e0071d7e3ae3f3f6038b5dbbd5ac18819fbdb425cd65d23aa6 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~I95b908a4845eb4b14e8f933057bab27e44c6a867e4bb02d87417740e3150e018 + 1;
            I5a26f98f9f83ddae2958fe17b1b3f0d2f7dc64309a438e2fe1f4b8dc87e5d1f4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id5d890ac1e6399e0071d7e3ae3f3f6038b5dbbd5ac18819fbdb425cd65d23aa6);
            I5c01e607e3f3ba8c06fa54e0ea9fdf0dea25c19c9eb317e51a670199ad40ea90    = I5a26f98f9f83ddae2958fe17b1b3f0d2f7dc64309a438e2fe1f4b8dc87e5d1f4;

            Id616fa98bf8bc6050ebcaa718c98c6dcac9ed2895a71b3a0d6fc42fd71205959 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~Idcc1ce57eae666070b5b9984cf69d5d2409ea92b36718906218185325b5611b2 + 1;
            Ifd0ce5d7e19da5ad023cf65265ce2071eacda4cd9553f0823662bc9569ecf872 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id616fa98bf8bc6050ebcaa718c98c6dcac9ed2895a71b3a0d6fc42fd71205959);
            I38fa842b13449763b8db07a9f91ab3479670dbc6043c1b363df6c93f6d7011b5    = Ifd0ce5d7e19da5ad023cf65265ce2071eacda4cd9553f0823662bc9569ecf872;

            I0e86f93ab7eab1ffc76fcb7a83eed533ad27ce0f06a15ccdbaeeb4c0293317f4 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~I114dd7172ac111bca494cc4230447a2dc167f12f198288d34cb5311c279a73b8 + 1;
            I91855e266ca0be3dab2b079bc241abd61a6724c1eae142ccc58d0a4b46fe2709 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0e86f93ab7eab1ffc76fcb7a83eed533ad27ce0f06a15ccdbaeeb4c0293317f4);
            Ie52aeb4c0ba45662d7f71f542630151f22c1801244258b9c8c20dcaed7f1472e    = I91855e266ca0be3dab2b079bc241abd61a6724c1eae142ccc58d0a4b46fe2709;

            Ie517400824ee7e75e8f286ac888007dc57c24fcb6707f0b369532fa6b0a96b4a = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~I30a86fd347fff855a807034e13d6e751b35d4330df8436470af7bb42af947668 + 1;
            I5a38f537a832431af9ac0e9070decc66ae16f850af8ac9349959011fdbf151f0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie517400824ee7e75e8f286ac888007dc57c24fcb6707f0b369532fa6b0a96b4a);
            Ie995e639d0338c10aaafa2dd930d57c74442bbde282aefcedcc9ac3b1eeee565    = I5a38f537a832431af9ac0e9070decc66ae16f850af8ac9349959011fdbf151f0;

            I4d5e1e1c63d137b4924c9e478035c320ae319e1f2a23433b9eaf3a537db29c2a = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~Id56cc1c8a7f6213208fea3ab1298a107ea854d908609dbe2358ba954989e1784 + 1;
            I180662d06f4e8f2216950660d1078c52394ea152dbfff6443f6983f3493caa89 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4d5e1e1c63d137b4924c9e478035c320ae319e1f2a23433b9eaf3a537db29c2a);
            I3b7705f03e900fd64d1b68f0b4036e5ef40c39722a2e6bc8ea6f22f91fb4b044    = I180662d06f4e8f2216950660d1078c52394ea152dbfff6443f6983f3493caa89;

            I93f155f57d9443e4b03255cbc0718355e5bec200a58bd83eea6bc11ed564ced7 = I5aba0b9a861c7337bb29f15b36c22a8292edfa6cf6a6db707d3bee735f8ebae0 + ~Ib1e8234d991235274c74ac026c33d868403b3d03a18a0c674e07dc4f94d614ff + 1;
            I5093a95294be69b95d3d4e3cbcd6a93f482b9a77f5214ff42a003cfdb5bc34e1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I93f155f57d9443e4b03255cbc0718355e5bec200a58bd83eea6bc11ed564ced7);
            I4656f355712fef190fb3697699fda1c25bbe9f7577a4d1a95aab55550fd7bfbf    = I5093a95294be69b95d3d4e3cbcd6a93f482b9a77f5214ff42a003cfdb5bc34e1;

            I7e0a468c76cdf4b3b95812da2dcabdd9992c595254d9c0a02d815dbb310c302d = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I6d0d8fc19811812bc80267dd50fc4742e9efceded7a9428707fac605fac90368 + 1;
            If6d7b3ad99d2259ce46cd080637bcf973f36b74bdf7b265d793f04aa27305ce7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7e0a468c76cdf4b3b95812da2dcabdd9992c595254d9c0a02d815dbb310c302d);
            Ie53b7792c539fa6f2aac95f09dd4a489c9167cf9d6d749f498ab99380c2e694a    = If6d7b3ad99d2259ce46cd080637bcf973f36b74bdf7b265d793f04aa27305ce7;

            I7f6ac9fe8ed957551d29e18ea194077943be18e78174e93c0ff4f9d3dac8f657 = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I9989d555a1c808f108dd152608d93b00d7a396de9492733ffd5165700c869840 + 1;
            I298771c166c7b3809860fdc01e1ee8e865e1c5f2b6a4492af4a9f2dbb6b0e0a7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7f6ac9fe8ed957551d29e18ea194077943be18e78174e93c0ff4f9d3dac8f657);
            Ie8270cd60cde73d16c5b65134dd393e02f413312f997a0344223cfe05d27985b    = I298771c166c7b3809860fdc01e1ee8e865e1c5f2b6a4492af4a9f2dbb6b0e0a7;

            I46d9e33c21650fad18bb70da588abee2fe9735680d0c187331e081c111bdc4af = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~Ibf9f290605da4b6295c786c6ebc135cffc80a3352b42e1d841ba5f6fbbf06cc8 + 1;
            Id2c03e9e66b771798f4ccfe5a9bebd633ac87eb38c9f211f1ce4d10950e5ef91 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I46d9e33c21650fad18bb70da588abee2fe9735680d0c187331e081c111bdc4af);
            I53d82131f37765f57bd586de5a55e92a697f63f20f366913802549f9ce658e68    = Id2c03e9e66b771798f4ccfe5a9bebd633ac87eb38c9f211f1ce4d10950e5ef91;

            I15d1b221d76c92d20200cadb2f0bb529c3b89164d7f67774ae33b2a01ea39fb4 = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I2fef37935343317384b1d29a04765327533fd87d4fe82a74f24b8196b3dffc92 + 1;
            Ie15e789de7ea93b8fae0ec21d465a7c42518fee4af3e1f9584e08b3563488c1e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I15d1b221d76c92d20200cadb2f0bb529c3b89164d7f67774ae33b2a01ea39fb4);
            I289dc39cab39ac30635179b9cd90bd31489a146c8c026138e1a1f9ef7a0ba30c    = Ie15e789de7ea93b8fae0ec21d465a7c42518fee4af3e1f9584e08b3563488c1e;

            I1f76b9ab604bd37a481f9327251fbb99d28272bea9f03133a4d1f97499a2b4db = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I1a6ae2cf67f356fae1ec533488e09c6696277823378b06751db7ec97115d9c00 + 1;
            Ie6b05d841cdf5f0f96018c49f9a88d21f39875c8f8af17d0dfb16b0d12a670da = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1f76b9ab604bd37a481f9327251fbb99d28272bea9f03133a4d1f97499a2b4db);
            I23d6a001aa9c80161e8b305bf34ef8d675247595457a8326a13fd348a02a1539    = Ie6b05d841cdf5f0f96018c49f9a88d21f39875c8f8af17d0dfb16b0d12a670da;

            If9a6c15537c6ae15c785c8729b2c059a320f316c98f777dcee42050c46990ce5 = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I9fc15e538a85dde7207e48d484f796d96ac712463c802b6995b216e71fb74d93 + 1;
            If3c580027dfedf572f89eb6a3ad9f82877baf03f3d6ddba81a8d868dbab61d83 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If9a6c15537c6ae15c785c8729b2c059a320f316c98f777dcee42050c46990ce5);
            I15c69e4ab6a25a44e8cb3ae11dfdf0e1dcf71c2cd63add1ab315e1d8a2d2043f    = If3c580027dfedf572f89eb6a3ad9f82877baf03f3d6ddba81a8d868dbab61d83;

            I10f9d40381df04200ca994a74c8a8d70730997334d739548351b8bb93dc29a53 = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I3c03db46b6474bbd284be2e345d2fae9939f0925a62da2ff9b1e2f3632740b0c + 1;
            I9edea5dd63fc137c4ea1044296f48581e5d5fc613cab5f0494a13a6241fa4b38 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I10f9d40381df04200ca994a74c8a8d70730997334d739548351b8bb93dc29a53);
            I36dcdce4926fb26d7d1b098549754fdfbc3b61a8947394227deedcb51ef1c374    = I9edea5dd63fc137c4ea1044296f48581e5d5fc613cab5f0494a13a6241fa4b38;

            I11b57b318e1a6ffe46a449f5031d9517c7b51452160307f7c0c414cbce227277 = Ia0863884d470eb62561ef6f23fd30359d70dccc4141e58bd04062afcbb8576ec + ~I7ba56fb0b187c50e86b74d8dfa7d7b3a1e2bc341cfb56a6343de1e7bb60742ac + 1;
            I468b553f5f3c22cfd36667c1c4f5743c10bc1632ebb3581b3f5151e5f79c6a51 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I11b57b318e1a6ffe46a449f5031d9517c7b51452160307f7c0c414cbce227277);
            Ic97aaa16a00e936ef8bd742c1c1c14696a72063ec283fcfd02962ffddc327cb5    = I468b553f5f3c22cfd36667c1c4f5743c10bc1632ebb3581b3f5151e5f79c6a51;

            I7b41563150c1630c478200a5a0a08a7809a1ae2d161450e63f10f4629308ba45 = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~I78023336da442165a8be56b4ebf7b41f4bb48bbc2b05c308dcd344c8f36c476a + 1;
            If5169c101f3b104ad3312dfa6e081e948c3354bc8a884861269c89dd7f8fe5e7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7b41563150c1630c478200a5a0a08a7809a1ae2d161450e63f10f4629308ba45);
            Ia28ac0bd59dbf550e8f75ac42fa8618aef3a8323a0e0cd6bc6dccd79c71fe396    = If5169c101f3b104ad3312dfa6e081e948c3354bc8a884861269c89dd7f8fe5e7;

            I9e477ebbbe435cede26f2d18e939f81f8da88b0089026282010e0f60e8d3e89a = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~I3464299c3a5abaf050c7176e4c0e17ade3cd5d6d86e82addf3e12d662def2b86 + 1;
            Ie88edc9e0f743d11046dfe95865fce6327d2f63bba8fc4911fd93ceba76cb03b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9e477ebbbe435cede26f2d18e939f81f8da88b0089026282010e0f60e8d3e89a);
            I70f499bcd8ce706da16f5d06d481e5197fda5d63b024d9850a34bdaf8f41c2cd    = Ie88edc9e0f743d11046dfe95865fce6327d2f63bba8fc4911fd93ceba76cb03b;

            Ib2254e933b3358a2febe2ee78bfa00d03502945608b8eb00f8b921077315df0e = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~I1ae7d02f524c03ca060c3dbc879653486c099ecee485690ce40a355fc1ed843a + 1;
            Iae0f73413a2fc8784aa61b30e9699da78e56fd7ba2fd8293e32cbc9dfe6bc114 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib2254e933b3358a2febe2ee78bfa00d03502945608b8eb00f8b921077315df0e);
            Ie7a936ed864922de2eca56a7a648d209cef422443181f89ebbbd6724f5bd0ee4    = Iae0f73413a2fc8784aa61b30e9699da78e56fd7ba2fd8293e32cbc9dfe6bc114;

            I92aa5d178a20d871c5226ec40b3c94942f20c06ab5351b9f0bd08586022f76b8 = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~I3efcac0fab0af81582237cdcd612c8d22eef1a6534816484190db28f3e7f3a96 + 1;
            I68165edd77863351062c8e0a09c1efdd3d244841d10f66ed22b25236c10b84ce = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I92aa5d178a20d871c5226ec40b3c94942f20c06ab5351b9f0bd08586022f76b8);
            Ifa54fad7897ca3a5db0d7fdf35cba73823e245f86c54af8a772f1d30f540247c    = I68165edd77863351062c8e0a09c1efdd3d244841d10f66ed22b25236c10b84ce;

            I9261ce4479f81cbaad6fbb8ee9c872d9dfdab45875f0af6c01c479990686fffd = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~I877734e2edefa267510037759c9490dae213d2e046beccfe87e16c1aeb5583c4 + 1;
            I6f3393df8a2c258b1c44d7ae93b7b9ebe39c27cecee6bc2acd3f5c191278d2ea = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9261ce4479f81cbaad6fbb8ee9c872d9dfdab45875f0af6c01c479990686fffd);
            I8c7c890f6f561a9a81130bf7ef4100851c3d86620903cb6b6d648746c0463b46    = I6f3393df8a2c258b1c44d7ae93b7b9ebe39c27cecee6bc2acd3f5c191278d2ea;

            I7def5551ef03ec4cae6129877ec5f900d6d7edbc6fc66f3f80de9a23b31adadf = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~Ie6ccfd08b7627ae7cdfd608c7054781099d7df5a0f133672db189134161f76bb + 1;
            I6189724f652320ab2c3d18de4f35ada1ebff4b32b2d3e86c66a3f2c74941172e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7def5551ef03ec4cae6129877ec5f900d6d7edbc6fc66f3f80de9a23b31adadf);
            I53795a7f407f9dd9d22f6483bbf9efb36313825abbc84c49e1885b01cb2724ed    = I6189724f652320ab2c3d18de4f35ada1ebff4b32b2d3e86c66a3f2c74941172e;

            I9e2c2192b5d360a53c35daad843eb9d5e18e850305732dac35c9213a45ca5d05 = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~Ia261f7672256403997417633102f8c1332ae17195bc38faf0fb85c4e4dd14da7 + 1;
            Ib32260d6129253637588b8358e00892c493347f945a010d24fe897e6a9f2eae3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9e2c2192b5d360a53c35daad843eb9d5e18e850305732dac35c9213a45ca5d05);
            I9d28182f6270a0cad620a562c047b449c03bc2036e855d1842707337fbf007eb    = Ib32260d6129253637588b8358e00892c493347f945a010d24fe897e6a9f2eae3;

            Iecda880e0e0336e9564a1eefd20e2d22e0ee56f103a90a56427a0af52069511f = I8b2a530749074d0c5d99ca93b607e52cf2afea530a2ba1548d5e06198ae9858b + ~I7f31f363b408908ca5cc070f150594db404279b7c5326f5da9abe8f60138bd51 + 1;
            Idce2a9ec74e8909d7514e546c058c4adcd18ae2607f3490cc9918249ce38ceb4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iecda880e0e0336e9564a1eefd20e2d22e0ee56f103a90a56427a0af52069511f);
            I2837d4f41e5abdb0abe8c9282938afdd85015263ad60e9a187ee91944f18bd1a    = Idce2a9ec74e8909d7514e546c058c4adcd18ae2607f3490cc9918249ce38ceb4;

            Ica0e4cafeb0b7c9e6caff0f66b45625890be48216b4a25b0fd582a72e2def407 = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I03527e99f5c488d7864664f339e2094fced797e4b46101f3c2bbe0b892c2d299 + 1;
            Ib8a985708ccedac94fd8d239571a6d5a2fe336ece2d15ee7d0abe9a79dc1e48c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ica0e4cafeb0b7c9e6caff0f66b45625890be48216b4a25b0fd582a72e2def407);
            I832e0057c56a4b0624a8ba7fc95565ff1322ef3b377d21b243c1fa69a9b83982    = Ib8a985708ccedac94fd8d239571a6d5a2fe336ece2d15ee7d0abe9a79dc1e48c;

            Ibdbea6826ae5ea65408f48eac06e1542cd2b3b0e1a4bbeba724c85ee552f1d6b = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I7def9ddb7ba2e414a44523f17bbff45806f0100ef624a52e91b03022877a7771 + 1;
            Ic0ccbd30732da760b3a4fcf87c08c87c22cbf26d0cd50785f80ddd7682b1fdce = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibdbea6826ae5ea65408f48eac06e1542cd2b3b0e1a4bbeba724c85ee552f1d6b);
            I81243c0fe8b8a3ab03ea4a07b48ae230b9783bc2b49006705893387b2eb0353b    = Ic0ccbd30732da760b3a4fcf87c08c87c22cbf26d0cd50785f80ddd7682b1fdce;

            I67619c07a6d53459465f2d77929930804aae53cbb52a97de1d849e532d9ce5cb = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I453d1e19585e0fb4fa66d684f0e6b37f56990cf101cc3942d5d4fc7e2313710a + 1;
            I6d7c4898670ee6aa4eb6fd97e1abacb7e4152c19d5e286e110420d2083a5412a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I67619c07a6d53459465f2d77929930804aae53cbb52a97de1d849e532d9ce5cb);
            I53e079434705c9ad3bf3e5cdf3f1d09bd1b0f7742fab2145a089e823e5c28f30    = I6d7c4898670ee6aa4eb6fd97e1abacb7e4152c19d5e286e110420d2083a5412a;

            I555422dd30763e140e02b9b6385eec9ea18ed35842a4eb56f68f861556d50adb = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I9c3d0fe7d767050217425eadb8e780e5eeeb31239f2f517ae5d122bee4157180 + 1;
            I48ec069746bb9dc6300ac6cacbcc382506e2c77773451d32f4d9fe4cdb43ba8b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I555422dd30763e140e02b9b6385eec9ea18ed35842a4eb56f68f861556d50adb);
            I77f3f1abf296aafc631f7b3d8bec79228071d4097f2083f70dfee8fa6ca52ba9    = I48ec069746bb9dc6300ac6cacbcc382506e2c77773451d32f4d9fe4cdb43ba8b;

            Ib6b064fc5e6213c920e8d2207427c6c27622bfccce85f662b0bb2e677990272e = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I87c64e9e81da569414617b07e39a7f67b0b76c71643cf7257b7374feb6fc9750 + 1;
            I94f08b3dab411dca5351bddf1de6f5e659685e48a5ef632fd7d4e52dc69d3dda = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib6b064fc5e6213c920e8d2207427c6c27622bfccce85f662b0bb2e677990272e);
            I1704967bdd23aca028c7fd652f9a0efcc55a31662c9f9b65911b7c1241205d9c    = I94f08b3dab411dca5351bddf1de6f5e659685e48a5ef632fd7d4e52dc69d3dda;

            I7e5e6e223f3acc5d6f776796e0be8f4806d5355cbe795331b0ef20ad3e12abe9 = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I90a0e50a5730714abafa98a7ad70e64903062bfe6f8deeb528bdd7008958bd11 + 1;
            I80e179604c153f8ad75c1e75837fbd86beec291776ff5363e2302f962998776e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7e5e6e223f3acc5d6f776796e0be8f4806d5355cbe795331b0ef20ad3e12abe9);
            Ia2313572dea3f44e7ec31d1474ed481064164548d3de394b69a6e99f60561388    = I80e179604c153f8ad75c1e75837fbd86beec291776ff5363e2302f962998776e;

            I1a7d235bf70814393dfca5c8eaa078813b915fa814648adc0a6b2d72e24d1d52 = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~I2edaebf9e3781f53167708c4854b01219957ff020915c8d2fa7b68e50ede1d66 + 1;
            I8608849b8538dae3f311153c3c70f026f5bce23c17237d20d192c838f0d890cc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1a7d235bf70814393dfca5c8eaa078813b915fa814648adc0a6b2d72e24d1d52);
            Icb8aee17be074ffae08bde14b025127c77773cdf482aa5fade629781c3488e18    = I8608849b8538dae3f311153c3c70f026f5bce23c17237d20d192c838f0d890cc;

            I4536ef4b6318344733197809b7d7c05af0bdcfb40818c16bbd525cfe55e1eb81 = I7c03e8d475eca2d3c8f4e595632ff2447d75342db24ca83978db801cf973249e + ~If0d87a6c6a4dd34bcb5411a845e6e7bc7fbeb0e6a34933f64283c880ca5d3d8e + 1;
            I530532adc42fb00f7f781e6b1d108a4d2444cddb08da7c6d088ae9f3d6b7f265 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4536ef4b6318344733197809b7d7c05af0bdcfb40818c16bbd525cfe55e1eb81);
            I4b2da3ec326ef0ce2bd1ef54c04f06bb0c9c7fe6f0736613537206d5f5568ff9    = I530532adc42fb00f7f781e6b1d108a4d2444cddb08da7c6d088ae9f3d6b7f265;

            Ic4910d74bc015f92940dfd059f327ed96a95ab01a170d3d00bb266061a7a157d = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~I950415762b14dbc0817ccfb0d09d95d700be57ecc9f8011c6163f84336da6e43 + 1;
            Ia75f7e68c65cb713bde41f32c61fd9b320c8f4474fa8ce88598372c0fe14c930 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic4910d74bc015f92940dfd059f327ed96a95ab01a170d3d00bb266061a7a157d);
            I475e873205aaae01975a2852b3d3d99aeb7ec9aa17759595012bf55fea91ff81    = Ia75f7e68c65cb713bde41f32c61fd9b320c8f4474fa8ce88598372c0fe14c930;

            I9022439743896e55957c8ec574d3e2e14f88e6baf4b65c4126cb39e589a92da3 = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~I7b25bf7d9020a7dacab3d15cd039a86780e41ed33520f5272ee788252efd1b9c + 1;
            Icca7f4c8f454e356434907ebb02b97ee9f5bc1e7cf4860adb16a1dd6a6b709bc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9022439743896e55957c8ec574d3e2e14f88e6baf4b65c4126cb39e589a92da3);
            I9d7892388f5775db1b77de0b60b10ed4f40c44774e1ca7ffc723e5fad503c487    = Icca7f4c8f454e356434907ebb02b97ee9f5bc1e7cf4860adb16a1dd6a6b709bc;

            I52412770a9e85565ac24e94df63da66b761a5e54ec1bc8c5c8b07b621a33a164 = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~I465489f86885351586de73a0aed556821e0ce34d1c2cebb67227004b4503eb3b + 1;
            I4214214ad8fd0512cbc2cdfcd1f1d11139d4a44c71628c5d2c1f00193b2dc777 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I52412770a9e85565ac24e94df63da66b761a5e54ec1bc8c5c8b07b621a33a164);
            Ib459acc97fee8ddd325d7d8b18d5c339a3c1e03c919c750f88070ec8a4f8a0ad    = I4214214ad8fd0512cbc2cdfcd1f1d11139d4a44c71628c5d2c1f00193b2dc777;

            I43c4705413499cb45c94379264ecec3fbf0bcf83aaaaf0110c9f13309682d21a = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~I6f7a9d597443df1a96370dbd5e1c1f9cb563fdc4db1d00fa66e8a287fca9bea1 + 1;
            I3151a9171bac0e6e2edf837e6bca27cffc3df8c9971c3b3a6873cd8169f34fda = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I43c4705413499cb45c94379264ecec3fbf0bcf83aaaaf0110c9f13309682d21a);
            I25711c9c95cd06f19d25d01854fdb8290f4759c9133d1a0c9e88548b886050a1    = I3151a9171bac0e6e2edf837e6bca27cffc3df8c9971c3b3a6873cd8169f34fda;

            I815e9a6b98dc1542b276704eb99ea559b4b34a16131b14fe631575d5fdf64e66 = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~Ie72b5524b212840dd1e69f4fa41b4955ca028c1ea7fd2f3440843cc2ef6d4be2 + 1;
            If8249d9d116a929e5f3c900c84a36d456b162f7fcd71949c88fce1e080cdb72b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I815e9a6b98dc1542b276704eb99ea559b4b34a16131b14fe631575d5fdf64e66);
            If9e2ce38db8f4cb30a3748fc7ee1244c98a4ef3c6dc840123405c585f6a867b7    = If8249d9d116a929e5f3c900c84a36d456b162f7fcd71949c88fce1e080cdb72b;

            I462a0b49cb7c2a4940d2befa6f37a5c2aaed3a81d20ff47d528b821f8f9dd245 = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~Iea55b5544c098ecff239cee665c2642cce17d3b546df6ea3d0c832a118c535bd + 1;
            Ibce79851c8253df32d60965921c117f70bdd9b486aa72bb17bc3ad578bdee995 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I462a0b49cb7c2a4940d2befa6f37a5c2aaed3a81d20ff47d528b821f8f9dd245);
            I6b1a6a399505ffa0312c9c79ecca8d63de6c5a1c9f6c0590296cb316c22d114f    = Ibce79851c8253df32d60965921c117f70bdd9b486aa72bb17bc3ad578bdee995;

            I5f1a06fb6eaeb2fa30f132d4fbbf98080868dbcc827b35e3a3a75945cfa97ebc = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~I730afd6404f505477b32f86185baccd692e9e64865f66f048a93e33d1cac8df6 + 1;
            I6a9121933f24798dc7d6c4671e05f959e4514a894f78f0e6ca37a9cfc0f7a53e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5f1a06fb6eaeb2fa30f132d4fbbf98080868dbcc827b35e3a3a75945cfa97ebc);
            I5454f64581fced198aa8ed832feea4c5a3de221d45b8eb42ae5820d82e540931    = I6a9121933f24798dc7d6c4671e05f959e4514a894f78f0e6ca37a9cfc0f7a53e;

            Ie6a253c0afa00e08e20896c2d4c77582cd8c24ba00c3363830f057a7f321eb05 = Ifbb7947946d760523a399321ff45290bc8416bc5cbfbd3b45bb0ec1a2ea7a1f9 + ~I567366a85ce4a20ac4125a297426463bc2f2c71511a97bfe2f4a01f6e8da6403 + 1;
            Iab3c6e4766bca2055b7c11e462f459c0c69c45c76b11fd6aefe62006c7a1316d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie6a253c0afa00e08e20896c2d4c77582cd8c24ba00c3363830f057a7f321eb05);
            Ie2235e43965f0eebff14c5c279ef56fc3e4055cc263c20f8d993756e7a5d9b2d    = Iab3c6e4766bca2055b7c11e462f459c0c69c45c76b11fd6aefe62006c7a1316d;

            I1aa2c1de85f2c5fc04250c2fc277af4c7fa7072d9c7946dc8f6f240dcfa87c2e = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I305dec30cf8323b9af4b0a6d285a31b3f5afb2e79c1a2ea77ce70a4409a7c765 + 1;
            Ib645fc54982c8fb5921b1dcc8ec4737c61a564e50d7195d4d9214b231fa4496e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1aa2c1de85f2c5fc04250c2fc277af4c7fa7072d9c7946dc8f6f240dcfa87c2e);
            I72979b4880af333f9e67500779c23973ada097a3cd1e2d4dff0eed1c570f299f    = Ib645fc54982c8fb5921b1dcc8ec4737c61a564e50d7195d4d9214b231fa4496e;

            I61539a1a79c4785262e8d239fd7e9f5d8e7f8fee2526fe7b4057795b6e5a657b = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I81c612bc8b32254693a4a0c89fb21865b161dd1673f5610732b31dd5663f160a + 1;
            Ic7e0e378e8448fc365285c0651e01f06536e3adae7e9c95f309e7d9980d5035d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I61539a1a79c4785262e8d239fd7e9f5d8e7f8fee2526fe7b4057795b6e5a657b);
            I4d0c6d6a69f818fe0856050283b987099cd8c7f3c8c22fdc825a01734c4642bc    = Ic7e0e378e8448fc365285c0651e01f06536e3adae7e9c95f309e7d9980d5035d;

            Iacd51e59a644b3ee8d3b73b5c6e6b6b89586e869487aed8e8c3c6b86c5e82135 = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~Ia7d01a6ab6c0646f75030a0bd04a711a9c50dc4674c921680034012e67a0c3ea + 1;
            Ia325319a3b0f63d7d994b0e5ac83b8cab618c9f79ba7f60dfc0c32bb80c5c72c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iacd51e59a644b3ee8d3b73b5c6e6b6b89586e869487aed8e8c3c6b86c5e82135);
            I811e21f3227b2bc3bd72e9b312edf9bf8e88261543c6bdb1bb09607f49b8206d    = Ia325319a3b0f63d7d994b0e5ac83b8cab618c9f79ba7f60dfc0c32bb80c5c72c;

            Ia3ad491fb952d351e2ca1c3b3994976b3dd273509d86e95b341f2b609175cba9 = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I2ad4afbffd2865f5c89feff965381fdaf73ac9ba4bc6e802a39014fe554b09ea + 1;
            I2da0a6fb45c46249fce53133b82906b2668976ad484cce849bf7530b5c0420ee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia3ad491fb952d351e2ca1c3b3994976b3dd273509d86e95b341f2b609175cba9);
            I4e06a2f339c14dfd77c1d58f78598240d08a7fc156a785a8a3fcae2d2d6d0549    = I2da0a6fb45c46249fce53133b82906b2668976ad484cce849bf7530b5c0420ee;

            Ibf8e7c032bde3ca68321b7cbc2e86bfb0352bd5c21d5da458b3f98d751b3f504 = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I600d6bfc6bdecb80f4f9d6020bdba9b4c04bcb359e66e793a3bd6732173d0b17 + 1;
            I1e4f3c6c98d527ad3075a00ecc95decfa07785b7b0c5ff523ae53741ffe019b8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibf8e7c032bde3ca68321b7cbc2e86bfb0352bd5c21d5da458b3f98d751b3f504);
            I167bb55e57f960522bce657a28f3a58bb6d82aec339cd46a3e8c4136ee023474    = I1e4f3c6c98d527ad3075a00ecc95decfa07785b7b0c5ff523ae53741ffe019b8;

            I4d9675ed29efda87fa20ed542d67c88fb1782698b8879fc28e908d27377c939e = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~Ic4c53101c741f07c928018af5696d83f45a29d0e5a9f766bd2f1f1404f3eb59e + 1;
            I4fb260b26ed5bd044dca51e17dc1b4a7902157d61ba92c823b47e375f9944bc0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4d9675ed29efda87fa20ed542d67c88fb1782698b8879fc28e908d27377c939e);
            Ifde56fe010824d9eea62caa160db5bde8de47e31630cd6a8c5e0572df0fa0709    = I4fb260b26ed5bd044dca51e17dc1b4a7902157d61ba92c823b47e375f9944bc0;

            I6292a3c00e5ada17538f4bf8df9a28541f5d080a806e8104c49a89d94abe9ffc = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I481cb000cdc7a32db6aa5a6b0da57b76f53f5bec6ef93d4ee25557e1b12064f8 + 1;
            I2e94b3f49feae361294ef10579f5ddf4cd4e7656029492a1598cd5cb01a85887 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6292a3c00e5ada17538f4bf8df9a28541f5d080a806e8104c49a89d94abe9ffc);
            I1b81ea9b142b222ca4b90724e3c4facaba82a4dea5c9b05c66032b06a459706e    = I2e94b3f49feae361294ef10579f5ddf4cd4e7656029492a1598cd5cb01a85887;

            I96289ce0db8e685e23fe7fc2b1a700a4cc2d1938225bf444c320d7194f1ae820 = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I9ccd1f3aa9f849bfe7dd9ff5f9de6fff64a444bc5286321a1f0e73e990d6a996 + 1;
            I54c78cf957f6d08b1ef46a35ec24b04b3400321d670b4137d64e89399cd3c370 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I96289ce0db8e685e23fe7fc2b1a700a4cc2d1938225bf444c320d7194f1ae820);
            I3e9361e7d30732f3e689391f56f9007c32c2368c9eb9d85b933f798babb0da68    = I54c78cf957f6d08b1ef46a35ec24b04b3400321d670b4137d64e89399cd3c370;

            Ib1e20a0a29f77c9e1e9f5d4b6938ea3dbc0fd30eff663b54ca2a3e255b3075c9 = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I8029c5b828acc50a3a785cab42ada7d51c82647934a9dac7f4a738920f1a332c + 1;
            Ifcc80d9233cbe913ec2813cdf22e5da4f6a463f224ce7db93884c3b49e6a7a97 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib1e20a0a29f77c9e1e9f5d4b6938ea3dbc0fd30eff663b54ca2a3e255b3075c9);
            I1774935be7ae799801f3b949e3a99707c4b32e7b1538e9f63cd8b940295ea6b1    = Ifcc80d9233cbe913ec2813cdf22e5da4f6a463f224ce7db93884c3b49e6a7a97;

            Id5110d84643f22616230397f50ceaf2f51e6c46fb596eea856ad3f29c4385149 = I9feb397e4c5499c193137fd34621721d862974fda4ed9be5b1d102a2f0fc226f + ~I95d408de4742f651f694ccc8f61d215af1e9b9be2b3860dca46c143e03b3ffec + 1;
            I30472f7544755b800fab38e17aa914eca481774221aa925e5fc526aa7431c05b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id5110d84643f22616230397f50ceaf2f51e6c46fb596eea856ad3f29c4385149);
            Ia4f0bde88d8ea45e325a92c25209a97269d31e2e3999ffe83696236b611de74d    = I30472f7544755b800fab38e17aa914eca481774221aa925e5fc526aa7431c05b;

            I10b08e5e9575d53b3c52e32527e38bca0fad4f0ed25bddf20bfd1d454ef836e5 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~Idde70a085816497aa92518899b882b67eb7989897509c445847e24204f5e978d + 1;
            I2968bd466e64c0ebce5448acf7247671f5f669f88bff8cf1ed20b47e29a9f1f4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I10b08e5e9575d53b3c52e32527e38bca0fad4f0ed25bddf20bfd1d454ef836e5);
            I30378eb921b9521d10fa2953f99f0f362b986bac12404a78a5f50619fe3b55fd    = I2968bd466e64c0ebce5448acf7247671f5f669f88bff8cf1ed20b47e29a9f1f4;

            I9473ca20629c79a46dd6db402744d58ce1ad19d823d0f3f9ff6988c22f02dc8c = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~Id3bae057e39f6549ce13910da61dbb41693ff87efebfd241bd1410d3da7195ef + 1;
            I23dc7c83c84d15f94edcdac20ae49442bfe44709dffec43950a95b107b0521a5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9473ca20629c79a46dd6db402744d58ce1ad19d823d0f3f9ff6988c22f02dc8c);
            I972ff0b38d85487454c289292e792035f568f072c33914f87e1f9c981da34370    = I23dc7c83c84d15f94edcdac20ae49442bfe44709dffec43950a95b107b0521a5;

            I26657dbc109dc227769ffb9fe0418b97e1407634c4cb9d19d48337861333cf76 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~I6ffb18ff0417e140b26d84cece8d23ea507516ebb60dbee4438e9433713c9f81 + 1;
            I40480c0b76e0574c82a8375bf6c3c255f6cd5e8d9f3c09c5ddcdae498d43e294 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I26657dbc109dc227769ffb9fe0418b97e1407634c4cb9d19d48337861333cf76);
            I22ad40f4d98f11e2fc7b9a8d56e44092f6e319c4edb2a67c5d9dcacb6a038846    = I40480c0b76e0574c82a8375bf6c3c255f6cd5e8d9f3c09c5ddcdae498d43e294;

            I0867129ec512051e4846e12f23bb824b363561c6e2511511bddad44a934a9299 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~If6592aef798f1b26c5c6593d99137d00bab8e8631070e89dbc6a3e11c89b3e92 + 1;
            Idaf0d98b59e58bf2225f5790830f4162cfa3dc258f0bb9f84e81d33e2e2b097e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0867129ec512051e4846e12f23bb824b363561c6e2511511bddad44a934a9299);
            If52bfa5da5e6508360b34b20a9607809dc732ad7d40860c8677bb6983d8c30a2    = Idaf0d98b59e58bf2225f5790830f4162cfa3dc258f0bb9f84e81d33e2e2b097e;

            Iaa9d2267657be14e58cfc2369f00ccccf2d09b8711e2325c11eb099296260046 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~Ia0090ea9b75c69dfca34ac43abee88b20734f7afb9c1d88f95eda3df6aab27db + 1;
            Ia9202e23aadf215e5e8887fbe86fd5af4410c49d5dcd48ad38664a63e4a52a77 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaa9d2267657be14e58cfc2369f00ccccf2d09b8711e2325c11eb099296260046);
            I2e9200c7443fa92d38415a8988c0a7ae2366612db06cfc84d9de4faf53d7d1c4    = Ia9202e23aadf215e5e8887fbe86fd5af4410c49d5dcd48ad38664a63e4a52a77;

            I08db08fceae6dac922ddb30dc8c5d2ad75fbd5b6aa2f24fb0b42216c988e8881 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~I54feba5563ca84d4a04e3ff7ff5ecf689d26961daf0ce27f0be8988087296fc6 + 1;
            I911a22b33617a35907440f195ef34301e1abaef90df3cf6b455b7aab22aa7637 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I08db08fceae6dac922ddb30dc8c5d2ad75fbd5b6aa2f24fb0b42216c988e8881);
            If23a3c0642ef8cb4b2d375a21de5253ad97342b92d29b8b7417bbd9ad0fb2fd5    = I911a22b33617a35907440f195ef34301e1abaef90df3cf6b455b7aab22aa7637;

            I835263edaf6c3692cc0dbdcd536e403006ebb5becaf77abeac432c98f2a2e261 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~I8b151ef6b3125cf983140726d775d948a253c13f020d3d1e75b585afb979bc8a + 1;
            I8aceeead21c39681b7587f543140d493989947711214df2082211fddbe4467b1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I835263edaf6c3692cc0dbdcd536e403006ebb5becaf77abeac432c98f2a2e261);
            I8b801d7872264ef55cc09008ded93c39bcf86fcd83e472ebc91d27c953520017    = I8aceeead21c39681b7587f543140d493989947711214df2082211fddbe4467b1;

            Ic6522502026653a983fabdc7a97f3a61c6478884ceb2dbe7a61669f09dec40ad = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~I8bddc257a28da31b71dac60701bade264fbf14f8377b1f504ef874c72e0d45a1 + 1;
            I4a9ca51fe9e7ed20f97438fa441c48b74f2520d29c3c6f530f1317d014a4a09c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic6522502026653a983fabdc7a97f3a61c6478884ceb2dbe7a61669f09dec40ad);
            I727fdffb518b29e800d3761e94d33c96bf32b4006f248d8eeeb18a035a7c8abe    = I4a9ca51fe9e7ed20f97438fa441c48b74f2520d29c3c6f530f1317d014a4a09c;

            Ia9b3853d7376f2b3ff71063cab059c2e5b2b888b4bdd3ddf38c5b207fe5978cf = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~I96ba46d5aa5ea6b2cc6a43df70554584d43f49a6bb171722373d28a2b0f1caa8 + 1;
            I84b6567e6638ffe91637cb5c900fb87d964738c80c7a2bc3c02839e44c665bf8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia9b3853d7376f2b3ff71063cab059c2e5b2b888b4bdd3ddf38c5b207fe5978cf);
            I4b5a25e13e61b54b754dbb201add03176d432d0c31f3ee1a4086797eec57cbd4    = I84b6567e6638ffe91637cb5c900fb87d964738c80c7a2bc3c02839e44c665bf8;

            If869318b9b2eea76cb0f28203ca8bca23b5493b21f9dbf176915a73fa7383cc8 = I2c559f7b2937586c6d2d807306df830beca70d92f6fd4d303f17e2c56faeb6e6 + ~Iff8bdf9ea44924628e777925357dcbe728f0ef4be0a3574965c811485fb57689 + 1;
            I8507dfdc1822c3c555877de0a703babb888342a1cd4a5345593c0eb99d72f5c0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If869318b9b2eea76cb0f28203ca8bca23b5493b21f9dbf176915a73fa7383cc8);
            If4413af8c4f8f3dd1f90f00fb5067c95a240f9e3ba7271b134cfda0a1fad603b    = I8507dfdc1822c3c555877de0a703babb888342a1cd4a5345593c0eb99d72f5c0;

            I1f1a7cbe72daa5437fa96abc25ece5bb43cf13aa018be3537e107fad506f28fb = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~Ibc813c005ecf7c077ea48779116cce31bffebb300fab262a78d166c4e270e3b0 + 1;
            Id8bb5f8d242836821aa26e984a13318a5e507c6bca8479e9c2e3ef96bf24350b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1f1a7cbe72daa5437fa96abc25ece5bb43cf13aa018be3537e107fad506f28fb);
            I0640e35183fc639f884fbb98626d0d54556ba20b2a709c1b4eedad0d3e27ad12    = Id8bb5f8d242836821aa26e984a13318a5e507c6bca8479e9c2e3ef96bf24350b;

            Iffca3b5121937820dcc59668b1027b5276cc746cc65b3c8cee5adf9be0e4f33d = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~Ib33ee0ec338d1389ec9010793383d24de32231284e86a9b03fd2902743dc8a00 + 1;
            Ic21b3ee91f7fd6945933b2d6aa6a8136c92b40340e6ce286cc5f592b6d585a1d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iffca3b5121937820dcc59668b1027b5276cc746cc65b3c8cee5adf9be0e4f33d);
            I79f29e0d9e4930c0e8eab1a5fa373778c2663402943ae843e94dc1d3ac60192a    = Ic21b3ee91f7fd6945933b2d6aa6a8136c92b40340e6ce286cc5f592b6d585a1d;

            I0ca8ee6c12c754f4b5fbbbc35b5edf976cd2f3a819a967d4f7808544e759058b = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~Ie57f94a45eba4db3826b22e3eb6acfcfa04b6d0669e22e5b78dfae4e7659b205 + 1;
            I41e581525a6f6f7decc5d6b1fb34553b16517fa79fe019d523dc0de19975dab0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0ca8ee6c12c754f4b5fbbbc35b5edf976cd2f3a819a967d4f7808544e759058b);
            If41e7a25c141c9a83ddd7dbf5bcbb72f579ba7d25231b25ab91ecdd1b8c50af0    = I41e581525a6f6f7decc5d6b1fb34553b16517fa79fe019d523dc0de19975dab0;

            I09701bbd76150af027015cfe8cc976f8bea0834c8b3cb443f11baef2e0799636 = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~I123d4c26243478ad4cff3406be39503c6b378cdefa50bf60249ec03d3a44270f + 1;
            I154a0c43cc16258a8b281935bb29839d099e65ee46bc98787be8aecdef9922e0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I09701bbd76150af027015cfe8cc976f8bea0834c8b3cb443f11baef2e0799636);
            Iabb9a156ffea98c56dcbde6d29fd606deeb21debc4aa2629e41c035547d5a589    = I154a0c43cc16258a8b281935bb29839d099e65ee46bc98787be8aecdef9922e0;

            Ib7225c329ff4c63f38d638c6647b92bb12ee5063dfd2f1bfcabf0272878cff77 = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~I8954b3335e6848eaec70a960b632233aff75de56bd0bb895e2b4ae49095fe19b + 1;
            Ifbd920d2032ef4cd599ba64059574352b60ae0734a6cbed208f65e8c04ab2efc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib7225c329ff4c63f38d638c6647b92bb12ee5063dfd2f1bfcabf0272878cff77);
            I496dabb1a4608940824606478478a3050517d422cfb20c53c37523f34aa08a45    = Ifbd920d2032ef4cd599ba64059574352b60ae0734a6cbed208f65e8c04ab2efc;

            I78da05b970dd2ce30b2503f93922c4281e5daa812cb0aa255120e75ad946cb4d = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~I0011eafd50b7df59be2a4f143443c0ca8ea87f9a93586d07292ba02fdc2b9b4e + 1;
            I7b8c17efb60e592f131daf550ffa3dc4a692cc5892ce1bc726f9024a5a714bb8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I78da05b970dd2ce30b2503f93922c4281e5daa812cb0aa255120e75ad946cb4d);
            I8bf71b880aa8654933f2008a17308e8366b6f6f22f52091e06364bd10004b891    = I7b8c17efb60e592f131daf550ffa3dc4a692cc5892ce1bc726f9024a5a714bb8;

            I0a363fd35ab7009f60fb2c4f96f61326c370defc1103deedea40bf0d0159256f = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~I931537d878467c473ac81aec8f9a7d79f286024e62ada1e5f363b93d6887070a + 1;
            I12b9fcdf2336d8a724bb7131ee096233b51a61fb5150f5a622509303bf56d9ff = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0a363fd35ab7009f60fb2c4f96f61326c370defc1103deedea40bf0d0159256f);
            I1748e381924bfb743c1257d7830da580af261ef967ffdc1adfafee17c67693aa    = I12b9fcdf2336d8a724bb7131ee096233b51a61fb5150f5a622509303bf56d9ff;

            I806f8a32e68e72b07ae9fdb26d41ac1a42bdb0fd4ffcdee68fffd430b0b007a0 = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~I6ec3df474c20bfab5d99aca971523dec8454a5ad4536765f4f9bcb0c31978cd4 + 1;
            If3f507c6e543114ff388cd6b8eaa2ae808c46166e2b8badbadb1eaa37f0c04d0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I806f8a32e68e72b07ae9fdb26d41ac1a42bdb0fd4ffcdee68fffd430b0b007a0);
            I7412e7d6cab6a1cdead2bfb425b79f89328cf155ce5e3b7e8593a4abc457d4aa    = If3f507c6e543114ff388cd6b8eaa2ae808c46166e2b8badbadb1eaa37f0c04d0;

            I70c5e2d6271591901678b8f0e488d737b3cb603b8b8e448024cc9d7e0deba259 = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~Iff82ae02f527d0eff3c9f8bb9d8fc818cf9bb7e3fac1a127849eea6ba27a62d6 + 1;
            I7f46d67075a762da1edcdfcd9fecf3975109a4cc488f66687f81441a821bbabc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I70c5e2d6271591901678b8f0e488d737b3cb603b8b8e448024cc9d7e0deba259);
            I39fc2e50c10ec72f5df6ea43b36d62fae7c1c3cbf6f54e921133adc9d8ca884f    = I7f46d67075a762da1edcdfcd9fecf3975109a4cc488f66687f81441a821bbabc;

            I3546a9ead1e1b810503b6521bb2c34151dcce36548225099755e87bd323b21df = I1be6c47b8009ecf488578c28a9dc65952942baf50e542df3d4048a9ad63b7367 + ~If8c51307ae2c537425caa18b7c3dbbf0530e94ada2a2a600262f57f93bf60d24 + 1;
            I02c96d25df89a3bbd36a7aec220bc13566ead49f7fa02b64b96d46bb7cf8541a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3546a9ead1e1b810503b6521bb2c34151dcce36548225099755e87bd323b21df);
            Ic3be1c01d32bc2fd127d4c4b371fc566b3977bf6f5ecaf4fb7f662f7bdcb36ae    = I02c96d25df89a3bbd36a7aec220bc13566ead49f7fa02b64b96d46bb7cf8541a;

            I5466c771c60a3618aa4866c2b07d5b586e7d7c70934a747a04273c3367ae8abe = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~Iefd5db28023cae3483fe3f0f1dcd5e302d642a0b5750cfa9940a9a8d6326cdb8 + 1;
            I615191537e8873d55c3af429ce9e1019bda129cab124ff2dd1ca60465f185faa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5466c771c60a3618aa4866c2b07d5b586e7d7c70934a747a04273c3367ae8abe);
            Ic9bd71f61271b1ff2f37d36580487d70287b498a51770475819cbfe50d3e48e6    = I615191537e8873d55c3af429ce9e1019bda129cab124ff2dd1ca60465f185faa;

            I83d8a4e44b0c8c27a4ff0338985fea545759f3660b941608878feff2c4208c82 = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~Ie11729721562e4a52a189a242aba934be636847d35de867cf00d26690c69abd0 + 1;
            I33a3c95ff1b26a9158939189358494e93f924d9b8bc3a4032bbc53d5b7b241d6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I83d8a4e44b0c8c27a4ff0338985fea545759f3660b941608878feff2c4208c82);
            I5217a6046ea279ff9f6f40af49af30f0cdeb374e8c2543da9bb27ce89b08044a    = I33a3c95ff1b26a9158939189358494e93f924d9b8bc3a4032bbc53d5b7b241d6;

            Id4e193d0a39e2ff4ab10d577523c3d264b54fa0a698b4ed0aecb5ddf075a4acc = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~I3f5dc950ac82420b73e1bc98c8c412f7e91958fbf455413c6a0ea5b2569e078f + 1;
            I9d8024a69b10baaf37cb9911eb275f1a827b75cc590c9830cfa90f1892ab1a87 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id4e193d0a39e2ff4ab10d577523c3d264b54fa0a698b4ed0aecb5ddf075a4acc);
            Id8c201e2467b255d627059eb66fab4ef48d0c235488dc0f7eb7c350a1d39467e    = I9d8024a69b10baaf37cb9911eb275f1a827b75cc590c9830cfa90f1892ab1a87;

            I779445414027b5e440b1075ad92e9c743a919e539757a4305d3985b57cf1ea50 = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~I8cf1c2115398eb404050fcfc654b198694d3c54eaa592d0d725b15e7937d8cd5 + 1;
            If683ab5a719cfcc8aea312c7be75e5fd3e2dae0d517ee14a136b1181209760cd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I779445414027b5e440b1075ad92e9c743a919e539757a4305d3985b57cf1ea50);
            I89de4a293c5da110f92bc9aa9b6ecc790b2fb3e1d282a6373d5ddaff63ef6518    = If683ab5a719cfcc8aea312c7be75e5fd3e2dae0d517ee14a136b1181209760cd;

            I9cf43907a8c090249537efb3105ef878ec38cf189b1848dda10fa0934cf6f0c7 = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~Ia9160306dcccf07d591c6c85cf86175408905d5e1bdfb36206d9c4bb5b917dc4 + 1;
            Ie3f9871ea280c6b53533e62c3927542a4c4dd28ff2c551ecd1166b9775315390 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9cf43907a8c090249537efb3105ef878ec38cf189b1848dda10fa0934cf6f0c7);
            I66a3806824b2190f9af7e907d1b4e068fa12560233a9a67bcfc8835373d6d78e    = Ie3f9871ea280c6b53533e62c3927542a4c4dd28ff2c551ecd1166b9775315390;

            I946b706dbb3722bc8069bc60a27d6525a81955d0b22d8c06d5730b117bd8050c = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~I390750ab5fb20d9be34ce0e294c95ca61ab6e511578b636301037a34f9bd9c07 + 1;
            Ie07ac76b3131e7a779a284315a5adf27af7b970781350c076b5f5b6d74e7a45a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I946b706dbb3722bc8069bc60a27d6525a81955d0b22d8c06d5730b117bd8050c);
            Ia7af92f6f7d9e7629ea5a0dc73f90acb4cb2dd8694485491a528df10a2b00aea    = Ie07ac76b3131e7a779a284315a5adf27af7b970781350c076b5f5b6d74e7a45a;

            Ifd3de8ffeb5f4768dce5d08e6e10e4afda032d8e4ad7e88f63c50adfbe81afbe = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~I8b5d8146640c84b84d0d6bcb2362fd5bc7e7462e1905b32b998b1f00f2da3645 + 1;
            Ia9746cf96c8460169eb7c522565deb2322a9984aecdc1473193f1cf0ed5542b7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifd3de8ffeb5f4768dce5d08e6e10e4afda032d8e4ad7e88f63c50adfbe81afbe);
            Ia0e8b0cadc0431f58baf6bd1e0fc4ea9babaadf97f47eea75ce07e41cd0e8822    = Ia9746cf96c8460169eb7c522565deb2322a9984aecdc1473193f1cf0ed5542b7;

            I2325959aa541dcc2298076e643b12a8a9656b31c28607ec3204bcb786729b88b = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~Ic3d44900d87d02e6912d962514abecacc6e1f20fb71c052d58a896c5524e1703 + 1;
            I4fb36b8d1dfb44eaa85b9445f8966900fcbe3e895daeb0451d5e23b9df6676de = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2325959aa541dcc2298076e643b12a8a9656b31c28607ec3204bcb786729b88b);
            I5c3df19631206eafab24135f4eff9ad9449c874e02c4fa9770d4fc4ede66b3f4    = I4fb36b8d1dfb44eaa85b9445f8966900fcbe3e895daeb0451d5e23b9df6676de;

            Ib8801db7c3d797fee2cf63037daafac592616e4a958094ac2d7a85bad398c437 = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~Ide09a550a1cc61dd543f2dd7a6e38af908474f7c815ab70318871dece429d0bd + 1;
            If922d63aac5ca5dafe88f6470303e1e0ba23c90de33d4bdc8432a3c81dae9fb9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib8801db7c3d797fee2cf63037daafac592616e4a958094ac2d7a85bad398c437);
            I74ae8440b495f97712924217bb791b022bbfc59b228632b7f96649f2a2fa053e    = If922d63aac5ca5dafe88f6470303e1e0ba23c90de33d4bdc8432a3c81dae9fb9;

            I64e64024cc00dbd7a3a826c0f9d82dacd15415b344d86bda10ed4d0142fd592d = Ie18a8b814a56ece19f87095efe1088cb5a1b4df110b9baab563c6a7fbff5b9f5 + ~Ia71d81a2779b6eb5f39fad80ee4e7bbcf394b97657cb094aec163180224939e3 + 1;
            I759f10838f0b7e3f75c8762cedfbc1cadbd61af8f7ab3a9e7d88bacde6dc9c40 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I64e64024cc00dbd7a3a826c0f9d82dacd15415b344d86bda10ed4d0142fd592d);
            Ia9c79734a6daa19386ecd68dad6da50274ac40a694cfd496dc40736cb4b33da7    = I759f10838f0b7e3f75c8762cedfbc1cadbd61af8f7ab3a9e7d88bacde6dc9c40;

            I658d4c16a7bd3c6d82219fa10195aa78c15698af2fa5f3bbde967e29fb4fa8db = Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d + ~I9c110ac43d6a359d54082ce347cfc9885dba985b743aeb66bf25962b4539a6e9 + 1;
            I7541dae782ef8b038f2768096ba4fff06fa9fcc6bcb72ccd9b8fe5768ea28941 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I658d4c16a7bd3c6d82219fa10195aa78c15698af2fa5f3bbde967e29fb4fa8db);
            I8d71dedf25220f16c883b67bc750a6e3c8886a6238f13693a22b41345296b0b5    = I7541dae782ef8b038f2768096ba4fff06fa9fcc6bcb72ccd9b8fe5768ea28941;

            I2e7b8e10124f284adebc18b9edb14644f54d024c862e86b76f5d4b04aa2bbc7f = Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d + ~I58ea58692cbfa8283ab19d6e609fe472aeb9da51d3f3616a9069eacfb18b0bf7 + 1;
            Ia13360e2c05d42edd07ecca114d163efa53ef77481588add80343fce0a426d24 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2e7b8e10124f284adebc18b9edb14644f54d024c862e86b76f5d4b04aa2bbc7f);
            Ieaea96e9413e940b5858f87f12dd18ef7c88b6e84caea900505a50fe657e21e4    = Ia13360e2c05d42edd07ecca114d163efa53ef77481588add80343fce0a426d24;

            I1a054e117ce979becaab2b848f8b5874cef5611170ed854e8536c94d310b3ba7 = Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d + ~If7454cbad692d8d1ed806663944dde3d846b241d1f69736da66374c5e54b8de5 + 1;
            I611d21feb8ebaeec639386a89b1cf2bf5144303d16d80b557265f9c66a00c1d6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1a054e117ce979becaab2b848f8b5874cef5611170ed854e8536c94d310b3ba7);
            Ic8d159cee07bee92aa9171ca69177796c91fa7542a63970a29d785b3cac2f30c    = I611d21feb8ebaeec639386a89b1cf2bf5144303d16d80b557265f9c66a00c1d6;

            Ic15c7d8a56833e13814c297cf7982b48a42a0d89cd37c0a67ba3c3528546c240 = Id7c762a3e42270a0bbea98a9f7537c85f51e2e0bcb67499c829f45b47020fe4d + ~I0217d8dc004467c4c431dbe27dc564c042c33d06a5be72a29ceab927708c4de5 + 1;
            I2b59fa34c611ba64fd61ffd1ba77f01508c0122f8e8b2e2aeeee753603349e2b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic15c7d8a56833e13814c297cf7982b48a42a0d89cd37c0a67ba3c3528546c240);
            I4aee30afbdf3dfb74a29ea9bc15aa1b0d200331984b528fade3be76c3249e3f3    = I2b59fa34c611ba64fd61ffd1ba77f01508c0122f8e8b2e2aeeee753603349e2b;

            I79f4cc267149652c039a1084e89dec27f52317ffdd1f4e813053380c7f38982a = I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf + ~I9841a5dd86a1b359b25fb293e74cfbd88b34e11f22bb61170ecc921048620dc9 + 1;
            I4f44a415623a311f037559bed8d19a2cd306a1b12af2f9d015adbe009152908f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I79f4cc267149652c039a1084e89dec27f52317ffdd1f4e813053380c7f38982a);
            Ib48fdf999d6a37fee27e903a4581bf51bd4307f83a7a18c3d7fd5ff5e8490a4f    = I4f44a415623a311f037559bed8d19a2cd306a1b12af2f9d015adbe009152908f;

            I7b69470ac56b2ee8391293d6203e4fb6b7a3a605f38fc684f2eb1ff49faaf1fd = I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf + ~Ic98b2baa4c4b3d4541ae5e7f9ae0b032d4dee98ebd73901690f561438ecfe5ce + 1;
            I65abc9fbfc8e631136259f0a5f47d007c810303995e55de1e7e9f7ccde035fad = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7b69470ac56b2ee8391293d6203e4fb6b7a3a605f38fc684f2eb1ff49faaf1fd);
            Ie581e7d5885d31995c15b699ff1c7f397dd32496d88a5a4c77d1c5bcda532212    = I65abc9fbfc8e631136259f0a5f47d007c810303995e55de1e7e9f7ccde035fad;

            I7a670a21ee5fcfc5f08786bd903f1da0c55661633e25495ee189a3dd55244f0f = I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf + ~I6483bb2ee2f7c35aa35adc7fcb6cf8cd426e048f4aff95cb9f4f732f97adaabb + 1;
            I1f898aceb1ec1cc51f6b9f99e3f9d813eca57d9642b5e41ddf6175c6abe7740d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a670a21ee5fcfc5f08786bd903f1da0c55661633e25495ee189a3dd55244f0f);
            I317cbed94b414a879715617065e78d4ac271816f7f331e5545ba55a46bcd9a5b    = I1f898aceb1ec1cc51f6b9f99e3f9d813eca57d9642b5e41ddf6175c6abe7740d;

            I1cb1d387b00274ba18c42d1329f0bbdd5b95e586049a8230d94772d73597b47e = I2f42623859770f5d633abe24dc20ed735a7760a646a011a6d0c09ad2b70890bf + ~I14102f52e9c6fa58677dbf1260a5049a6c2807b245f123cecfc3f1a413badded + 1;
            I8e2ec7ed430c3dc4cd717cc7a6961e5e7c636d451837ee16a456a1d04d6247cf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1cb1d387b00274ba18c42d1329f0bbdd5b95e586049a8230d94772d73597b47e);
            I76b80ce969069fa14c6d7022d6c072434dfaed48bb2b30aae77035d134019afb    = I8e2ec7ed430c3dc4cd717cc7a6961e5e7c636d451837ee16a456a1d04d6247cf;

            I3f002730cfc58d827800579d570d0433b30d2f387e44b0641fd4004f52c01c27 = Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47 + ~I15e7d6b702e93b31ac4e46f9ba4cf63da33641629eb9cd414d1e2c8cf54b750f + 1;
            Ib9ff76d8c63a43b6873b5f305c93676bcd412530b04ebe4afbbbaa27a6b8f25c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3f002730cfc58d827800579d570d0433b30d2f387e44b0641fd4004f52c01c27);
            I732d56627c4f920af6fac9e623551f6c4c0e5e970b37e4d2f3b0dbc0d2491e29    = Ib9ff76d8c63a43b6873b5f305c93676bcd412530b04ebe4afbbbaa27a6b8f25c;

            Ife74c161a8f2dcf48e3a3b07d65523789eb2aeb2cc2aaaad88cfd91683069b6c = Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47 + ~I8ae4ec097c879009d8316e76b0a2ff9f4228310728d8b4dc196543a3976d26e3 + 1;
            Id3b55be9a317757f5c0144759a5adf67c44a5bb4afe4e60ebeb3be4ec94b1fc0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ife74c161a8f2dcf48e3a3b07d65523789eb2aeb2cc2aaaad88cfd91683069b6c);
            I7c758d1653b4abf515df4c565803d4d5130fad01c8b46a5d447571d0fde55bb8    = Id3b55be9a317757f5c0144759a5adf67c44a5bb4afe4e60ebeb3be4ec94b1fc0;

            I9bb3d89cfaf62aa40cae73b77d1a1ac2999465104de1d7c188918432e1a17c80 = Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47 + ~I1f749b245e6db4722494bb36009a7da73ca94f408d8a0ca7829b6d5258f78e4d + 1;
            Ic3e25c67909179600ab8e63f0335fdb849cf0166472fb983fefe68e9f4f9df7f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9bb3d89cfaf62aa40cae73b77d1a1ac2999465104de1d7c188918432e1a17c80);
            If8ee177b4825244aa2459f76ce3cfe5435b03e72d750c440474a42fee5009643    = Ic3e25c67909179600ab8e63f0335fdb849cf0166472fb983fefe68e9f4f9df7f;

            I82aaadd76fa8b5e7bd489cced1bc3b825f8e281accbc496474db7c4ea4d1e1e2 = Ibf3b12352dee4ae53d1113f86a1cf7a593c01bb07575ff33f1a4beb166c56e47 + ~Id71b753d1cf473f4f4bb7718f412471692e08afc0ae9d25e617c2360df79ceda + 1;
            Iabafc2aaab132f1976385bb8e128f51ff86417dd26b96e57df8e56a2b7044d33 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I82aaadd76fa8b5e7bd489cced1bc3b825f8e281accbc496474db7c4ea4d1e1e2);
            Ibbffe343259cc28309085b16cf40fb046a0a7c9d5dcef49182ab8ba0a9acbb2a    = Iabafc2aaab132f1976385bb8e128f51ff86417dd26b96e57df8e56a2b7044d33;

            I790d57f4f5730ea4166cba282bf1350f040ad2bbdb8863311b0f753991858960 = Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804 + ~I05a7291b0f3122dd9941bdd5ce72362b3b0b1803abb126606c82744979184be8 + 1;
            Ic6492e40db63085730ca2ab4612ce1d9b385e004b467ac433bd9dee4b81990bd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I790d57f4f5730ea4166cba282bf1350f040ad2bbdb8863311b0f753991858960);
            I6ab2cbc5eeb87f6f79360ad8b27bcdf5daad4c85f829eaa00ed855099653be55    = Ic6492e40db63085730ca2ab4612ce1d9b385e004b467ac433bd9dee4b81990bd;

            I7f9bc5d4b3aedfd4e192fdf7774ca874dd2973d41203f33deb2dfee1f3d5eb90 = Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804 + ~Ied43949ed7bc9c0c92af912b9e283a3e674d42242e0fe8e3d9132738d512fd23 + 1;
            I697243100d9508441bb98b0849280bf0d47509aa42f7f334968a19113ea5091b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7f9bc5d4b3aedfd4e192fdf7774ca874dd2973d41203f33deb2dfee1f3d5eb90);
            Ib928fe4e8b8da0fa26516833082019238c839091b1fb32c244e57a2aac417273    = I697243100d9508441bb98b0849280bf0d47509aa42f7f334968a19113ea5091b;

            I219aa384cadf0adcf51cc6828ca3dd9781775e7e7986955e6dd5074ae6bf0887 = Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804 + ~If434186e818b5a899ad4add63d67ba1dbed823165df4559ee78b39d8c758c727 + 1;
            I8b4daf5f5619a17e4bb744ddd92d5bb1a30a01e2928a200d796dfdb9f7594c1e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I219aa384cadf0adcf51cc6828ca3dd9781775e7e7986955e6dd5074ae6bf0887);
            Ib59d2666a9c62eea256e01a7e240af2a1c11a86a51058e6ed4034007a881acf1    = I8b4daf5f5619a17e4bb744ddd92d5bb1a30a01e2928a200d796dfdb9f7594c1e;

            Ia682b7cd027239465bf24461fc4d88457ca84c607032663699d76d58992265e7 = Ia3666acc01fa45f4659cfda4a0710e05580bd50a9e632336f82fb21e3c415804 + ~I443558f78c6ebb16bcd49ca586ea62d2ba12ed3bade0e54ae9bb60f83d2598de + 1;
            Ib2534e75a32847d1999b520266575471effb319ae660aef5e38d0aaac66f83a8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia682b7cd027239465bf24461fc4d88457ca84c607032663699d76d58992265e7);
            I0eccf85cb5b32056038d4f13293549f535d994925067f49a8f1abb6253ed45be    = Ib2534e75a32847d1999b520266575471effb319ae660aef5e38d0aaac66f83a8;

            Ie226e795a9a67a0d9984f30a164ecd2aa0692100a18a77337c2efae4395ff952 = I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b + ~I44089ced0a31e79af650baaa02274890b1f60ac7398745a0e4da4b2242f849c7 + 1;
            Ibc4f182435db6e718a7fde25165e26678a904f8d7372ecfcdacfff50c99c0f79 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie226e795a9a67a0d9984f30a164ecd2aa0692100a18a77337c2efae4395ff952);
            I5c11c8d23929c41fd11d326b4535976b5e6ad33e2969128e4ec4ccfb0897a22c    = Ibc4f182435db6e718a7fde25165e26678a904f8d7372ecfcdacfff50c99c0f79;

            I393c6e437a6f283fdacba0192edc09f7a8882ce8c6516d0284b10a6ed2a43a27 = I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b + ~I18e4b7dc3295cc6f5968878bde7abe5447cebc77dce83fce47db55be2237efc9 + 1;
            I4927222cb1738667a383028851b08d20223cac5a89a663b6b443bb2ee77263a6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I393c6e437a6f283fdacba0192edc09f7a8882ce8c6516d0284b10a6ed2a43a27);
            I7c9db5ef7c22e9722e1811495675725bc9367c52f47417ac0127b2ece6c2b6d5    = I4927222cb1738667a383028851b08d20223cac5a89a663b6b443bb2ee77263a6;

            I8ed39202419d4320b8d1fd945da1efe6befa43abd55b3ad1c7917b0587cc3950 = I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b + ~I0f75d5771cfa314d28e188de297b4bb53c2cb732724a630e10580ee5fe87cb23 + 1;
            Id1c743f39e92313845da6e20dafefce9dd80e43c11314962f5fba867c037687b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8ed39202419d4320b8d1fd945da1efe6befa43abd55b3ad1c7917b0587cc3950);
            I3d113258d0831ee2590c286fb25bc418e5c1d0033cfa04428717bc3782db11a5    = Id1c743f39e92313845da6e20dafefce9dd80e43c11314962f5fba867c037687b;

            Ia66d77f2baa846741b30c7f9b8d0f770d488b658b6d2ce6c265f8de5dcdc3af9 = I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b + ~Id60b48bbf346bf95a242f425de7f456aaba5b3ed35cf16a07ac541ca8f480319 + 1;
            I580cb70e24ddeade0ded45cff406069ff648af95813a3d1ffe82fe9916894680 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia66d77f2baa846741b30c7f9b8d0f770d488b658b6d2ce6c265f8de5dcdc3af9);
            I37fbc80705b247541af9b0468d3bb960bd4b8c1908084a570dc6435714c0f2eb    = I580cb70e24ddeade0ded45cff406069ff648af95813a3d1ffe82fe9916894680;

            I939a2a515cd6383018b9d98f9c3b748c75abd1beaa52e26c273eaed8978e9372 = I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b + ~I9d23867d2eb5d9dbcc21e9242aa71e141a2ecad61f5ad2bb69d798b2fdd1873c + 1;
            Id402959580cf99cd1d64f703a31be57b6a1b1eb883b8197096068729df11b293 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I939a2a515cd6383018b9d98f9c3b748c75abd1beaa52e26c273eaed8978e9372);
            I04ca88712e988bdef397bb8c4e680b6709f92094d54013e6d786aa459174baf5    = Id402959580cf99cd1d64f703a31be57b6a1b1eb883b8197096068729df11b293;

            I66a18b0e3441516bc7212f5564b7d2e079b7a73bbc481c67c4b357fa3a766f4f = I3d03f9caaf0a58d6df25f99b394467defca88935158a9cf421bfe2190234e89b + ~If5c2310896ae5dfd3f83de1affe79fad0f0b6b2b673efbceb7d296b33a6900e7 + 1;
            I1e19af5e5f4b25b16be3d56eb0b7bd5261c3ca95a38576983db444d6655809a2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I66a18b0e3441516bc7212f5564b7d2e079b7a73bbc481c67c4b357fa3a766f4f);
            Ie8303e1d3cd1305166144c2a9c72da17dc5ff4c6afdb56ea458d2c017a90fcac    = I1e19af5e5f4b25b16be3d56eb0b7bd5261c3ca95a38576983db444d6655809a2;

            I6e91dbdb1c31ffd16d890119d91969004497b13d180320f54a27b001b8814f3f = Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 + ~I4c8a0d23fea7158b5e99eea187df1d25395edf7df1db8482b41dab7a8bc25030 + 1;
            I87b00103000c17b5d537b5f7fb82eee037c57dc6b6a3a4cd43a19a92efd8b213 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6e91dbdb1c31ffd16d890119d91969004497b13d180320f54a27b001b8814f3f);
            I9c8296a684c3ac2e51841b13d88cf64656b4d2f7ac1625a77e0cbed908eb5f8a    = I87b00103000c17b5d537b5f7fb82eee037c57dc6b6a3a4cd43a19a92efd8b213;

            Ie0b0cb7147d168ab10e2a8d7c9c839e509d8e967d163eb11c4afa8738c06a266 = Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 + ~Ib2fff9999fc00e81b173cdaa0737f3e4f711ccd0034a6611e0e9111acff3893f + 1;
            I57ee78ee192d7bc07ed64d3d42bbf209e954cb023f7725e15482335cbcf402a2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie0b0cb7147d168ab10e2a8d7c9c839e509d8e967d163eb11c4afa8738c06a266);
            I70b00c7b7fd70b24b225260cda2515d3d5df30d630e9fab4b9f85d810f441649    = I57ee78ee192d7bc07ed64d3d42bbf209e954cb023f7725e15482335cbcf402a2;

            I54327a37a56f54ad389401b3e67be69eb0a6ace8d0f5ef507f5edfec4cb60f33 = Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 + ~I6ec1c8ffb963fef21e978fcfd0268bc24dd283819081437974fa5a06caa64c25 + 1;
            Ibba300f2463e7761c495190751b83704f8a828f727ae23b274c153bd605c758e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I54327a37a56f54ad389401b3e67be69eb0a6ace8d0f5ef507f5edfec4cb60f33);
            I891eaf9692501bbe1df2bd2f2470be83664f12d9e6211b5523bd7500a1e9fc70    = Ibba300f2463e7761c495190751b83704f8a828f727ae23b274c153bd605c758e;

            Id6ff08336ff69aeb7c86ff3c649c59079585a9117b8366ff1776938c76509345 = Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 + ~I7f3447e248449854eb030c79bc32b602d376441a193e25bfcf9b8a0eda83b57a + 1;
            I302b994f71bced52060f5016280bade3df63be8e6348e8137dbf09ea339b2ce0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id6ff08336ff69aeb7c86ff3c649c59079585a9117b8366ff1776938c76509345);
            I807e8a0a095e42d08f8682b77d262989f5440738b49f26eda30b3e70efc7a8e3    = I302b994f71bced52060f5016280bade3df63be8e6348e8137dbf09ea339b2ce0;

            I74cae7d7ceb41afef5f215f9e99e5ea1ee0d38efaa91800a240a26b49dec44a2 = Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 + ~If550dcd8751a8725d597ff3b723c6b5cff949b2e3087c71d36782ea291f7bd3e + 1;
            Icdf358bc87f821358185d6b64ed28411a009602f1bf397ff98dee49cb851087a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I74cae7d7ceb41afef5f215f9e99e5ea1ee0d38efaa91800a240a26b49dec44a2);
            I24a328d80a0dd14fa15ad6101cafcef8008c5846474fcd62cfde858dd3d75461    = Icdf358bc87f821358185d6b64ed28411a009602f1bf397ff98dee49cb851087a;

            I73d3f78f124fc07e4dec71f536f875a26946b68478ccd830fe94b24d6dc73f0f = Id5d41bee31f19baa9d9b84d916ca50555f797ed877b4b900e903d80aca077600 + ~I7d078740e07b48774c64f6dfd7bb0f56821dd685e014f0b9d4e3b7da45383e34 + 1;
            Ia74859916985880396078b181652782883d5e69db172af2bd6b5abf5ca55da72 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I73d3f78f124fc07e4dec71f536f875a26946b68478ccd830fe94b24d6dc73f0f);
            I8273973db378daf42a5ba6dc50c960e8433a2dcb5d17c30f95be6bf89ec0f0b8    = Ia74859916985880396078b181652782883d5e69db172af2bd6b5abf5ca55da72;

            I0dbbf32467809debc31db520a1d652a39c6f32927d5fe8e7bd87a0ccaf5dcbdc = I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 + ~I26e6175466ec922073d5092cb4168f87cd1289008e4b99400c5b6c2fec3eaf5b + 1;
            I76b090fba89f431fd007a510b3d1be2527c10360521dfe032cb18928fe5e5e2e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0dbbf32467809debc31db520a1d652a39c6f32927d5fe8e7bd87a0ccaf5dcbdc);
            I7ecba0b25a70555c9243a99717462e9f43cacafcbb2ce9b03d34054858620493    = I76b090fba89f431fd007a510b3d1be2527c10360521dfe032cb18928fe5e5e2e;

            I4bd4faaa74b900831991b7a4ce8511a5bb45c1ba413ef0d2516ae105cc00c740 = I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 + ~Ie6d2cd42fa78c1cbf17c7f18dfb4c0cc5f79f1fb0bda02dc92192252f99dd047 + 1;
            Ie19a52435cba71b7b88711d46eb5d530a9f236e6a6a2a19c9213d0b527e90719 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4bd4faaa74b900831991b7a4ce8511a5bb45c1ba413ef0d2516ae105cc00c740);
            Ied4b1e4e915dc6bf15ce0f505d7ac9fa6c5b8cbcc5831cdf270791ea45402c8c    = Ie19a52435cba71b7b88711d46eb5d530a9f236e6a6a2a19c9213d0b527e90719;

            I7252a8cf8ccfbfa3d707c9f2ff6b0edab9675a6e54f6e03a8cd7f06f77d2eef0 = I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 + ~I31adf91b5f31b4232ee24f82af27e02a7ed1f8535c552409f353690340b64b2c + 1;
            I7541dea08da40dee1671fed651faf2225a9205f04627982312ea6d8eb94ae3db = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7252a8cf8ccfbfa3d707c9f2ff6b0edab9675a6e54f6e03a8cd7f06f77d2eef0);
            I2b2b4121708eceb760e2854c76289daff432118cee2479045dcbd8ebe358e3cc    = I7541dea08da40dee1671fed651faf2225a9205f04627982312ea6d8eb94ae3db;

            I8534ec2afd654d78899e86e2eac05d7f62677fc213d962a50b1fb5d853c5b966 = I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 + ~Ief01c27ce040b3f50c19615a8f5d9bc8b467c0f88a778888fe186887b19fd580 + 1;
            I879436c6762d7a1f92f45aa9d70bcc63e0ca0957f69d2bd417c5a4410f4b24c0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8534ec2afd654d78899e86e2eac05d7f62677fc213d962a50b1fb5d853c5b966);
            I8eba7f46df1f21311e46e2657b38d61800060add0c96dccfa9c45fae66711d7d    = I879436c6762d7a1f92f45aa9d70bcc63e0ca0957f69d2bd417c5a4410f4b24c0;

            I07de1ee4eb883d98b9baf6d4b08768203be9277a5780b0b713b054c67b6e9362 = I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 + ~I4dcd8811ecf9d39f66ab4cf1e07e739c7972e9cf2ef9ff6c0a948336e22dcc90 + 1;
            I1c46edefc42352d5d7c429376d363db5a76ce8d5ddcc76e2da909f07c270a48e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I07de1ee4eb883d98b9baf6d4b08768203be9277a5780b0b713b054c67b6e9362);
            I587e2742d73f804efba3b90efacfca020ee8a5e13c2a490ec60ac494be39a275    = I1c46edefc42352d5d7c429376d363db5a76ce8d5ddcc76e2da909f07c270a48e;

            I2dbb829ee8781d23865b9bfc192543f10ab2839afd1a8f8211259f1248d89f28 = I1e49cdd13dfa3980fc7fbc06fc362431d632e180f21a562c007508dbce5fbfa3 + ~Ib3562b77830a64f31728e11cc54a6d19b55344891eb82355e3fb4491086e8808 + 1;
            Icbda121f4b7c783c142a1034a6b893200c3a974ca08b153ee0ecd6baadd03099 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2dbb829ee8781d23865b9bfc192543f10ab2839afd1a8f8211259f1248d89f28);
            Ic4766de4b982a051c7546be035a94bb07bc822061d5bd46d9a4070d026b7a593    = Icbda121f4b7c783c142a1034a6b893200c3a974ca08b153ee0ecd6baadd03099;

            I1c85612795fc824409767448d6770bcca93caf10fc2cd8659a98eb808c878444 = I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af + ~Ia2952eb350b07a9cd76752e1a5f76814ed095eb0ee2a284f221b1c74e38d822e + 1;
            Ib7a3b0d88758dcc368ea5aa65eb4c638502d363b70ebb303394e701e588d2a82 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1c85612795fc824409767448d6770bcca93caf10fc2cd8659a98eb808c878444);
            I5ce28b3e49d61224902a9c1f675a4032351731bd0d14cf3bcab007b30d7e5c22    = Ib7a3b0d88758dcc368ea5aa65eb4c638502d363b70ebb303394e701e588d2a82;

            Ib2c9dc402fbacb1f26f72f8b1f1578f70d7a69d30751d4e4661514a819b1a974 = I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af + ~I123e1ea1b1588abf2d5d4ede7027783bfb20d60ce3fdf365b86c9f5c84956a72 + 1;
            Idd87b9bea69d81d0c6e4a3901c764fbae4fc8b0795bae1176b2f5b75ce571d04 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib2c9dc402fbacb1f26f72f8b1f1578f70d7a69d30751d4e4661514a819b1a974);
            I07afa69acae532add7b503ba1bf357b95ab120399bc63d32e65af6f61a369f15    = Idd87b9bea69d81d0c6e4a3901c764fbae4fc8b0795bae1176b2f5b75ce571d04;

            I9d10906535c09c58cb10aaa6c3ba524ec6f2bf3bbe58da21edf42dc791662b04 = I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af + ~Ie14918150ed723163714038f6ffd2c64b07d62079dc03ac8fdeacde45633def9 + 1;
            Ifda52cd13144d30d66a9a0fb8b6c68ceee044c33751a0f3864b564eff21bf815 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9d10906535c09c58cb10aaa6c3ba524ec6f2bf3bbe58da21edf42dc791662b04);
            I4c0f888abd9ba96ae660c5a3f6e9c627c5775611d7a2956fa3049c5574fde7df    = Ifda52cd13144d30d66a9a0fb8b6c68ceee044c33751a0f3864b564eff21bf815;

            I2cc9acaff65bd5636a9def070cb29149ff8834daa39d18594d09d6156003739b = I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af + ~I4b15e4ecd6a6f2139463d94eb4061a410569136410e469abc38dbf8cc03948a2 + 1;
            Iee4a4722007fd835cf2b8e7b244a8f72fd79b0f418fae3ef31a50b35769a3b0b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2cc9acaff65bd5636a9def070cb29149ff8834daa39d18594d09d6156003739b);
            I4bb74c7a5d5fa7f8a3bcc33e4aac51ace977350ac258b3af687b215c37407b49    = Iee4a4722007fd835cf2b8e7b244a8f72fd79b0f418fae3ef31a50b35769a3b0b;

            I478e7d5b826a54848c89bdf12a8fa4b7ca31e387d033563784c60c493cc633f0 = I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af + ~I843cc48bafe9c4d2e4647f2909064999da8c2f4d8dcfeaf533fcd12c32c37ce0 + 1;
            I97604434d22669367d9ace3fdacecd4f777dc9759b5940d5cff195fcb0881346 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I478e7d5b826a54848c89bdf12a8fa4b7ca31e387d033563784c60c493cc633f0);
            Ia781a129677ad67c301dedf105bd58147a815283dd2c06d65ca7ada0aca7cc7e    = I97604434d22669367d9ace3fdacecd4f777dc9759b5940d5cff195fcb0881346;

            Ied5920560e9017a8c035f2d6b019f9abc3c8ac6dcf213cd3e422f92510ff38fc = I7e676a02869d4953f3b0703597514cb5de8354a59a7ad9800620920aac8169af + ~If7d42431922752de30d5506e1d501f65453a4754d7cab03976695cdee9c0c9a4 + 1;
            Ib0c6a201e2d38ed7791d229f2df4ce0605197b5edb176ffd5369d85764de153a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ied5920560e9017a8c035f2d6b019f9abc3c8ac6dcf213cd3e422f92510ff38fc);
            Ieff7f5ac404485dc7719d026c898a08cddf9eac3289347c09da180a04400da13    = Ib0c6a201e2d38ed7791d229f2df4ce0605197b5edb176ffd5369d85764de153a;

            I50780605e408ffc7501e94d92284899a4878c5721680a9d734ef276a4c9974e2 = I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c + ~I1308b215c5082a0407de73f2273fc035460ca21b553479402290c244cdedad76 + 1;
            I69f0a9020d4480b3ab0eb58ec235ffa667587b7da910b3854f56cb49e9047d47 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I50780605e408ffc7501e94d92284899a4878c5721680a9d734ef276a4c9974e2);
            Idbea312fceb0d3b89f626dc27620dc564adf927f2587857f0c80926c0f323433    = I69f0a9020d4480b3ab0eb58ec235ffa667587b7da910b3854f56cb49e9047d47;

            Ibf3bba34d932e08687d92505ae09625c8c1cfa5c24d3d52273050b8186ecafce = I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c + ~Ib96bae85b07ff95f5a6716cad97c765010937888a28ad63b16eef3b6ae93b3d2 + 1;
            I9c2b1197b3d0c6879b675bf90f26c3a5ebd1cdfbf6f5eafc502ad622535df53e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibf3bba34d932e08687d92505ae09625c8c1cfa5c24d3d52273050b8186ecafce);
            Id1537778668b48b3115e7b1a3cde430a348b515e592a110c520b33226ecf7f47    = I9c2b1197b3d0c6879b675bf90f26c3a5ebd1cdfbf6f5eafc502ad622535df53e;

            I5af920c58542851ac5891f1f1dce969c57e1e7cd12a302a68528c7c02c86a524 = I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c + ~Icd850fa1e932d19313713c2d376413e7b81faea883442278fbc700a2238f6779 + 1;
            I576f9c047b4db49719b8ef7ff32de3de609df2969827ec22e91d8b1c929abd99 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5af920c58542851ac5891f1f1dce969c57e1e7cd12a302a68528c7c02c86a524);
            I4d749601335050fe4f61b7b9280c1f83ae58f99216ee191f039f6b94b185e74c    = I576f9c047b4db49719b8ef7ff32de3de609df2969827ec22e91d8b1c929abd99;

            I8559dbc457ce562bb8447f1227ae0c59f2566cdd93fd9051488863bb3e4aa462 = I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c + ~I02ff320cae73fe5cc67804e552bffba75496861f085869eabab140094a18fe90 + 1;
            I22d7ba6fcb1a3830055bf29a53984fbb01f70b4f9c309f6dbf0a2cb493f39818 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8559dbc457ce562bb8447f1227ae0c59f2566cdd93fd9051488863bb3e4aa462);
            I2a445ed5096a1929dc2ef74b28f3243c9e05c70b4e0aed9baedfe94c28d8e4ad    = I22d7ba6fcb1a3830055bf29a53984fbb01f70b4f9c309f6dbf0a2cb493f39818;

            I3aee441136da868b3fc343e6eb88d4a48a636677bf1188261315fff1c8898690 = I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c + ~Ia6ddd4cda9a70e95a6ff1a9369bb2851b90588337f2cdad6ab43fdd6c6e32fdb + 1;
            I16e5e8ec4564f64f3db568b15f064d343674e523b9f6ac2ffcdc1e64a3dcac44 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3aee441136da868b3fc343e6eb88d4a48a636677bf1188261315fff1c8898690);
            Iae58883a74ef0111e20be8cc9df222d4e0e213d390b08244a5361328ba38895f    = I16e5e8ec4564f64f3db568b15f064d343674e523b9f6ac2ffcdc1e64a3dcac44;

            I1aa8aad0f4f034c292c7799a12e5f7887263752b5f11909fb73b32db7c6d7263 = I78954020b3f152fca43c2c77d6b1545bd19744b90014d87e2469f889cc258d1c + ~I269a90aa42086a30a9b03141bf37e3abea46a1f1c06710baf2d052a5bb404248 + 1;
            I240e73cf6faba62b6fd94d95cc67aa7703cc8e96875b5dab437e79e7a384ccf3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1aa8aad0f4f034c292c7799a12e5f7887263752b5f11909fb73b32db7c6d7263);
            Ibd5a78278d93327ec1527d2329cb8bdc601611fa5ee53fc37e64259d6bc217a2    = I240e73cf6faba62b6fd94d95cc67aa7703cc8e96875b5dab437e79e7a384ccf3;

            I559ba5b3899cbbfda28e2b04083c4958d942ab0a8577e5e7b9dabc58053b7f6c = I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a + ~Ia6f33a5c8baa6ea053642148b8e414d0b9d17a66f4e71f6e44e1f6c6e3e535ba + 1;
            I3c8e8025305283334b1155f2e020f3909d725f3d656a9209f357f396b345bf9a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I559ba5b3899cbbfda28e2b04083c4958d942ab0a8577e5e7b9dabc58053b7f6c);
            Id1f021d678d21318bd8881474b337f0b540c16dc97a33c4fc3abc12bb662f4a5    = I3c8e8025305283334b1155f2e020f3909d725f3d656a9209f357f396b345bf9a;

            Icb53fd5ff0cc1bb11f4efa51be8b18e0455037e4718b955718ffdf5d6bd24dcc = I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a + ~I5a03d267642091bb2d177a6689d91b995983fde126d703c6474d730b455ab56e + 1;
            I236740a734448318d6759a5e14178c1bfe93f1d1f793768577105ac5ee42d6f0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icb53fd5ff0cc1bb11f4efa51be8b18e0455037e4718b955718ffdf5d6bd24dcc);
            Id4d52f3a7303153d65a86d328d1e7e5dcdd602d284aba3e104ee0528d9b1d465    = I236740a734448318d6759a5e14178c1bfe93f1d1f793768577105ac5ee42d6f0;

            Iee6c6b7151a6d52632c5dd250c0fd5c866ed5e07c96d8ba7ed0fbfb13b5cc9ae = I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a + ~If377629f88304a78a44bdac612907792b54c49caf9dbaf85b3061be5baa2f5e6 + 1;
            I4200e2460844e967c243fdd9ea3e3863aca3b8023d85311149c7b30e2d3ccc10 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iee6c6b7151a6d52632c5dd250c0fd5c866ed5e07c96d8ba7ed0fbfb13b5cc9ae);
            I608fc1c1a500a0fd76e9a326afc6c5a26d1cd78f1b150d970f5ca74d1d7a3193    = I4200e2460844e967c243fdd9ea3e3863aca3b8023d85311149c7b30e2d3ccc10;

            I54cea20aecb1a113601e099b4a28a9582e143bf7b257df21a059c2c561056024 = I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a + ~I225da3a8a67ccba14e13c78ca2ffd83b37ac9a961371f1aa617f5752b1bb337e + 1;
            I831a730b580c0d83322ab8cd6cf78e490b8e104fac72df3a67d75d029a18178e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I54cea20aecb1a113601e099b4a28a9582e143bf7b257df21a059c2c561056024);
            I7b2d4fe3f2c703eace8068da2810bc7bc190900ec3959bfc4a396e72ef5a8200    = I831a730b580c0d83322ab8cd6cf78e490b8e104fac72df3a67d75d029a18178e;

            I127ecbb26b8b54be69afacba0c7c900d1eadb8907e3337013e771e8afd15b8ec = I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a + ~Id4f16cdf2e148fb2732fdbe215ff0edd44d29c41dff8c5b307ffcb8305832972 + 1;
            Ib33753185ecae290a3ff7193c21cb9f11014cd9ab59194b625bd9fb1ddf99413 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I127ecbb26b8b54be69afacba0c7c900d1eadb8907e3337013e771e8afd15b8ec);
            I72d8c9fea747adec725ada83bdebc85126870df2cd2cb9f88d2d043635bfdd84    = Ib33753185ecae290a3ff7193c21cb9f11014cd9ab59194b625bd9fb1ddf99413;

            Ib655fac982e2ba3b34f9be933b8da91c7416d2add55a9225d8354e85b51c66d6 = I159a1fec90e3b4434be00ee0fd264b0879b065ef2783f32ec99ead912243822a + ~Id88de8b0cefd527c486f8239ff6f61d6ff86085e420d2be56ce58f4d82d78a7a + 1;
            I780dd1faa05c0ff00db1b222da69e706fa7d30b9522b0ec2b89f6b23c30366da = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib655fac982e2ba3b34f9be933b8da91c7416d2add55a9225d8354e85b51c66d6);
            I4f237165ee7800d1fd20968d90afd5a858b8ae73675c1a03b67be17159247ffa    = I780dd1faa05c0ff00db1b222da69e706fa7d30b9522b0ec2b89f6b23c30366da;

            I066453fa3220e314882976bf9b0e935d3cd7f5233141a89a6fb00390d245ed9c = Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 + ~I97449b979933d41c6555a04ba5ba6cae73e44b040387a504f6f7e2ecb763ad08 + 1;
            I9cdd258f7d667c4be0a7f3eb13f79628e9bc1c12c8cd9febace271ff54191872 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I066453fa3220e314882976bf9b0e935d3cd7f5233141a89a6fb00390d245ed9c);
            I333abb8de54c2cdc50519fe091024d9862592e0191ef4acb0b6e1b7c45701234    = I9cdd258f7d667c4be0a7f3eb13f79628e9bc1c12c8cd9febace271ff54191872;

            Icc27708504fa373a81980a39fe27a732fe8ed4d3e67838b787c8d633cd1134f9 = Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 + ~Ib6f695414c34a124de17de5cee8798a33f0968f7eca5143f21f88c228ffa6345 + 1;
            I5996255101f1029eab99365af8b51d34cd6ab7e8d3bdf19598c43c5fa910d513 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icc27708504fa373a81980a39fe27a732fe8ed4d3e67838b787c8d633cd1134f9);
            I6ef7e70fed5f181598201b2c2c0002f1251010c752be38c1f229c337e4a66428    = I5996255101f1029eab99365af8b51d34cd6ab7e8d3bdf19598c43c5fa910d513;

            I9dbb69baeb72fc989c784ef8b69a50b8acd0c076fbd3aea250967efda14c7ff3 = Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 + ~I8e89f3937a947ff09fef0df8085edc1dc09a36d7bbb39027d358384d54088060 + 1;
            Ibfece5f844143052755772dc83b99eb3b78ef024232c0d1c1ca251da508d3516 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9dbb69baeb72fc989c784ef8b69a50b8acd0c076fbd3aea250967efda14c7ff3);
            I75665f397a59da51376855f9b737164887c48da916cdadc4b4d1605f3d8e4071    = Ibfece5f844143052755772dc83b99eb3b78ef024232c0d1c1ca251da508d3516;

            I3027ef5a77a2956cd097cebac4348dffc636fa06b156a08dd403916fdf42d957 = Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 + ~I862b7b7769e1ce1579c40d6363e23230c9253630d97fe8abe72b80e8a8b5440e + 1;
            Ib3368641096566227d03c6778a2f243fdb3b21b67dc940542c24f4045931684a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3027ef5a77a2956cd097cebac4348dffc636fa06b156a08dd403916fdf42d957);
            Ie81e5c2a20cacfd646fdc8795e265386030f32624e917b5877a38d9790ed93be    = Ib3368641096566227d03c6778a2f243fdb3b21b67dc940542c24f4045931684a;

            Ia0f10f5c6d9dc1cbb77556836ef659a542681ea3f0bd54d0edbb2259e14e6c0a = Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 + ~Ia810fbec78dcd5215c217347900257a8f892a4805dc2365ea79eaff74af7e64b + 1;
            I2ecfa55d807d1228b72f0ad1afd67133387e87cfa537cf8a7619fb887e86aaf4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia0f10f5c6d9dc1cbb77556836ef659a542681ea3f0bd54d0edbb2259e14e6c0a);
            I9760a21471e149d0c56a22ba9a49f377439bba25562cdba484b355531562bd05    = I2ecfa55d807d1228b72f0ad1afd67133387e87cfa537cf8a7619fb887e86aaf4;

            Ic81c2a6ad2dd6d624ab25855269124b464c2d5dfa31e41fac639a888994a2ea6 = Idbee3f9bd5e4063907482d891afe489a3df56fbfddeb997f6fee01ee98d81f26 + ~I107db18dddc718b9fe7354d0f352f72df94ad4653ab0712d5765a495ec29242d + 1;
            Ieab494ba47e97c3d84f264bf6017276cb149db18ad24479caadf0c8d24ec487c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic81c2a6ad2dd6d624ab25855269124b464c2d5dfa31e41fac639a888994a2ea6);
            Ie9ad099032e87edfcc146b2b8fc401eb78cd1c370d99a7d87b96cffcb2bace7f    = Ieab494ba47e97c3d84f264bf6017276cb149db18ad24479caadf0c8d24ec487c;

            Ifd84bbe3c8b82cd5fcde5db6c40190c17411a69c9502007d0392efb1b0507c87 = Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 + ~I9f0d592f1a57b1d3e2c206ffe5a79185253205dfe7b20be53091145aa16f9719 + 1;
            Ief87170e911c48a4f8f1830ae52e6b34421df444bced0e8746e004999ff5f39f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifd84bbe3c8b82cd5fcde5db6c40190c17411a69c9502007d0392efb1b0507c87);
            I42d22931f7defa6032679880bb907c668d62e4c65343d359f7ee0679bb098ef2    = Ief87170e911c48a4f8f1830ae52e6b34421df444bced0e8746e004999ff5f39f;

            I4ae6345c74a23a9713c9efd40683df95cb7d8f18163ecc526a0188b17f0ff54c = Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 + ~I781bae0d109036c417f71e00a3df3440df3cecd691fe1f67c147c4d2de217f7e + 1;
            Ia1e1fad227b8e563997b52484713aec367521484f20e560a7dcb2780bf2e39b0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4ae6345c74a23a9713c9efd40683df95cb7d8f18163ecc526a0188b17f0ff54c);
            I5d35fcce50496260be81878d7799638cbce05d2afe98817fe9c53a675ee5f98d    = Ia1e1fad227b8e563997b52484713aec367521484f20e560a7dcb2780bf2e39b0;

            Iccfe7f8fc79fb4b135af4cf2a698e9ef2614e7d01d137304a0b51502ba34a79e = Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 + ~I288ddea916663f74bb339e7a94ac9c86412f39671ca69dc7ec1da05a1800092b + 1;
            Idb4e9f7ca3ef03a86dc723495293aaa4ef9783f92a3b05b3344ec8468f9675dc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iccfe7f8fc79fb4b135af4cf2a698e9ef2614e7d01d137304a0b51502ba34a79e);
            I0876112eaaac7d4bd5dda75039d334a15e6d500f29e0c471e8d6dd0ba6cf70e9    = Idb4e9f7ca3ef03a86dc723495293aaa4ef9783f92a3b05b3344ec8468f9675dc;

            Id99854c623c0f1fca0e55e9b6125fbad754c4311497cac1ea4af1471342b7f15 = Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 + ~Ibdb62dc1ed705231a9d0a9e819d824f81e62746fd6d9877557622a8293c7cc3e + 1;
            I677395b9f313591599a7200d68572fa3eb1b30aa5a4bc4476ddd9fd840f29edb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id99854c623c0f1fca0e55e9b6125fbad754c4311497cac1ea4af1471342b7f15);
            I612926c7fd5a7811c91d55336a1ea5a427e4c28826227d05d2e08d501bb032d0    = I677395b9f313591599a7200d68572fa3eb1b30aa5a4bc4476ddd9fd840f29edb;

            Iffbb3bf56ca327afb4dd8826363aa655718ef15e14e5a6b9e55664d0cfc76738 = Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 + ~I48c76be33e4d7a127ef1f7eb5f4952f81439eced5be914ff90aac6d963267659 + 1;
            I6001c8b3acc2e47f7beeda5c633fb76e0f191d6dce473637683c7f6efe4d3b7f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iffbb3bf56ca327afb4dd8826363aa655718ef15e14e5a6b9e55664d0cfc76738);
            I4075a88832d68ad5005c73387153538516b97eb30d8d1bfc9f3d205cf338e042    = I6001c8b3acc2e47f7beeda5c633fb76e0f191d6dce473637683c7f6efe4d3b7f;

            I6f62760d6931ff9476617433db3f760557bf58b267224286d0f1f38777f1c19d = Idf99ab13a9e6b4caa69e639a456c37b413a844acaccfd49198a4d8c27677d326 + ~I642c0e5f0768f835a6ca3ee6f65875346121b502770acb1ce833e9aed46d4ddc + 1;
            Ieff52577c0d3fdfd35282159bf2ce744dc12f879d290abdd6f38a0f8b5241dfe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6f62760d6931ff9476617433db3f760557bf58b267224286d0f1f38777f1c19d);
            I4471c46046bb6606ad97bff8b36a4a9c1643c861791e8b3bf97a41e8cb385220    = Ieff52577c0d3fdfd35282159bf2ce744dc12f879d290abdd6f38a0f8b5241dfe;

            Ib5197b3ded0d4c6cfea1aa9572fc7eb7b3e0afc3b5afff40dc48c2fc2d06ee81 = If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 + ~I4a91f2655f96c11b03fce33601bc8f71a0fef4dc1782f7158126cd8cc5a1d690 + 1;
            I9bbf9a8a49255908ad3f62b8c4a149837fde63060eaa2d01bb382fcf59e9edb8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib5197b3ded0d4c6cfea1aa9572fc7eb7b3e0afc3b5afff40dc48c2fc2d06ee81);
            Iee30715a934f261b8e1fb4814e196f3307e095ec0dbfcb10ac1fcaa1d1d16372    = I9bbf9a8a49255908ad3f62b8c4a149837fde63060eaa2d01bb382fcf59e9edb8;

            I421cb52dd669a636801d3709f62f6570b289aecb322b1afd2ffdcbcb5f1377a7 = If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 + ~I10ecf0f58ee2fd15e2b4135dc03cb4053c364660c6d2e2bd03cfc37aa6d6621d + 1;
            I9ae8a856ac9eb44659cef37d3140bcef8b5253afff93a2b3e54eec5c88b6ebd6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I421cb52dd669a636801d3709f62f6570b289aecb322b1afd2ffdcbcb5f1377a7);
            I8b323499e4c61f57b164a287da64b2f1c933376dc7ec202d666ce57ccffc139f    = I9ae8a856ac9eb44659cef37d3140bcef8b5253afff93a2b3e54eec5c88b6ebd6;

            I44643d87119bfc715397cbbd514f7a75934db3d6fb8308d0874dad36e6ff0969 = If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 + ~If023ae056e9b4b370bc83a2d5604602f45a01a005bc19a769c874536faf4abbb + 1;
            Iac850cacadce02a577a7ae8d4d48b52f43aeb883994730d170d89c9f6255c4af = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I44643d87119bfc715397cbbd514f7a75934db3d6fb8308d0874dad36e6ff0969);
            Ic936076da3dcc6a7f335b0d3b428e8b01cfeb9240df6dd50bcfb2188cc37ae8c    = Iac850cacadce02a577a7ae8d4d48b52f43aeb883994730d170d89c9f6255c4af;

            I016081dfe95a2bab40513c2f55287a990f0b79588fe1b8286174ded6b93bc278 = If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 + ~I32a7df875889c28b6d8f86a42071ad142efd5a66d6328669bcdf1901a225079f + 1;
            Ic680429748da0cb695397674fbfe3bbd5f2b5496795b05051d9a62e0c7b38884 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I016081dfe95a2bab40513c2f55287a990f0b79588fe1b8286174ded6b93bc278);
            I1cbbfb485fecaa90d26f81a89b89c0d778558fbc218268369c32c33117c33468    = Ic680429748da0cb695397674fbfe3bbd5f2b5496795b05051d9a62e0c7b38884;

            Ib70f45a310ffb94185cae456609a25620a223187f0c4c3a9f8c5c645054ebb96 = If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 + ~I446e1574b1d7bd427fed19be1920c5c29a3276d9ec816ebe1e4465cbb762b1fb + 1;
            I617715b25070e943cf4b34892f49447ccca1e24e4182820b36e87194ca7edc1c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib70f45a310ffb94185cae456609a25620a223187f0c4c3a9f8c5c645054ebb96);
            I5bd88b9b16b4fbeeecae426d343179b982f46fe09abc37e1db23e03a43157b89    = I617715b25070e943cf4b34892f49447ccca1e24e4182820b36e87194ca7edc1c;

            I4e13170eb723e9bca567d19c25b56d782987da1f75c5a54ab26d0b1538f779e9 = If2ef14928c7840e037723fd9d5ce95d4162e795000290e118aab16ecd31f0088 + ~Ib699efc076bd227e0138482c43c5fc8cf0d0d87078e063262fc4b537f554697f + 1;
            I1eabd1ad44c5bacd15cba04670f5077da1ea3950e797f2ad5bfba62060a161a3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4e13170eb723e9bca567d19c25b56d782987da1f75c5a54ab26d0b1538f779e9);
            Ia5fcf505c93f7902d4ed6f1877bf51599e910bbcc6002e122623c389e72e2600    = I1eabd1ad44c5bacd15cba04670f5077da1ea3950e797f2ad5bfba62060a161a3;

            Iaabe2ac34f3411032dac139922cf9783f86937c5d525c8730c8ccdb257f94f2d = I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 + ~Ia441ac067e28123cc7cd9d005d0f5a1628da5628d4473db60d61b85c61e8d9b1 + 1;
            Ibd5dbd51229b1ffb3fbc33d4567e89a5b5767d759821c0b4761e8b1cba3fd021 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaabe2ac34f3411032dac139922cf9783f86937c5d525c8730c8ccdb257f94f2d);
            Ib2ed8f97504f1f2331d11107b05d538282eba6248d7d8fc3c9ccbb4a0cfd7e70    = Ibd5dbd51229b1ffb3fbc33d4567e89a5b5767d759821c0b4761e8b1cba3fd021;

            Iaa84c2b3b1d95fcb9ff86fcc68a6049f2c0c0c34101bf5bdecbb6d72bee244df = I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 + ~I91cff501b877ec0153cf2d85abd12870d65d1aa997a6bea7d653bf387813998b + 1;
            Ib59b40982a0fa0730bd4bc1b740c68166cd0db83909258e2d0db220140f7ade9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaa84c2b3b1d95fcb9ff86fcc68a6049f2c0c0c34101bf5bdecbb6d72bee244df);
            Ia2d0125fd752a306fa45115b7d888f2eb705d6f14d3e5d4f5191024ed7b1f746    = Ib59b40982a0fa0730bd4bc1b740c68166cd0db83909258e2d0db220140f7ade9;

            I79cc31e6c010fa8eb54cd33d70364720a3290ac19ba06f27ba05b1bdf24d6314 = I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 + ~I5fa215eca11a15c7ad85760cc87a0f8e883d02472c7af460b13cbe214a596c62 + 1;
            If3a3d8a238fcc1d5703240350b6f311213ce4d203c859b54a8ddfbc6af08e9a2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I79cc31e6c010fa8eb54cd33d70364720a3290ac19ba06f27ba05b1bdf24d6314);
            If45da818944a7fc1d4baf55234b4a8299f0513f6db7e1e8cd87e7b57f72eb817    = If3a3d8a238fcc1d5703240350b6f311213ce4d203c859b54a8ddfbc6af08e9a2;

            I045079845680e722358f1a61dfed5b3758b7d491231d08f6f6e674dea560885c = I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 + ~I5e14fc93aa39853d74e7844854278275828d0f5428f2af96c00c8b0ab141c868 + 1;
            Ie1a01aa1296ed81d5b75478aa0ff85cd0866be9418bb8d44d257087fa4f6b345 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I045079845680e722358f1a61dfed5b3758b7d491231d08f6f6e674dea560885c);
            I18d435d55c2e6ef05cdc85c7c5f1fc2e74307ca98333e485f5fcb8eb038dc3f1    = Ie1a01aa1296ed81d5b75478aa0ff85cd0866be9418bb8d44d257087fa4f6b345;

            I43e364076c55650d4376369dd211f84289220dbda754e9f3475b5d1310d66659 = I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 + ~I0d58818dc0f3ed67f1e3a10ddc7cd0592bfcb8cb3db1c329edea24dfb0ffde5d + 1;
            I01eaac160521c659f8be7398b4b66d448fdd6958d181bc148938a1aa3e3fd350 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I43e364076c55650d4376369dd211f84289220dbda754e9f3475b5d1310d66659);
            I6b9155f4e226a633f272039c862d58cbce7e31a597a37e1be49eb81b0b72cf47    = I01eaac160521c659f8be7398b4b66d448fdd6958d181bc148938a1aa3e3fd350;

            I0b9df0d909722adcf9aa8ee430e388b6f201b7f66e12c3cf72b4751fd4249b6a = I7ad4681c2d1a3ad6608bdb638dece92d45578e30fd5d2b056afc9de24d86fd50 + ~I8e0d77d4d38cb3b1e5ece19e010043e9a4f0802819f3e70f0ecc9440f65eff4b + 1;
            I28e7f4c19cd1f47169d939f8c94bceb96e0801b0a66dad9dcb1d2c3a1e656d34 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0b9df0d909722adcf9aa8ee430e388b6f201b7f66e12c3cf72b4751fd4249b6a);
            Ie7dce49639675176aa767ea6d5b2171e0c72deebe4e007b620860a1f8b177060    = I28e7f4c19cd1f47169d939f8c94bceb96e0801b0a66dad9dcb1d2c3a1e656d34;

            Iec9a71f06ec498907631c7b9709bc6461d2b77efe8493e4815501c56083727ec = Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa + ~Ibbcaf468c4ded9be4d2d82d059bfad5174f330444c98aadb71831769a32f70c2 + 1;
            Ic97e339e12a03eae013d5cd740b137561bde6188c1c9b31f5d39199bcf287b23 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iec9a71f06ec498907631c7b9709bc6461d2b77efe8493e4815501c56083727ec);
            I8043c8446ed3aac742a14c3df20420bdd5f0e6561e15c32f4045e2ce8b6f3330    = Ic97e339e12a03eae013d5cd740b137561bde6188c1c9b31f5d39199bcf287b23;

            Ibe52a5b5286c8d781c590bc26cd000c66c7ab759989f65c747574503e47867f2 = Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa + ~Ib6dfa3959980c5d348630e2edd81fdee8429a3003b0a21369b99343bda03e2a0 + 1;
            Ie83bcb1fe72e7583b427cb92e77a596a158312c89c2ddda3ca5ac113f7e8e58b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibe52a5b5286c8d781c590bc26cd000c66c7ab759989f65c747574503e47867f2);
            Ieb807bb8e9746d06de25556b579e51494e760b3a4312caa4862cbf2776acbccb    = Ie83bcb1fe72e7583b427cb92e77a596a158312c89c2ddda3ca5ac113f7e8e58b;

            I55d30fbaca443183b73eb12a611cece679d3b08098711ee7a74767fdc25d8ade = Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa + ~Ibb72bc519d54383d213250311085f6368ead1c943881ccc23f944e652f934063 + 1;
            I8e634f64bc4def7608286b21abd3f531fd18233e92626d134a8b986175008c38 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I55d30fbaca443183b73eb12a611cece679d3b08098711ee7a74767fdc25d8ade);
            Ie1f84176002d4791b93729913c6021f1ffd76c58ad11593dc088cbcf2e4bc4c9    = I8e634f64bc4def7608286b21abd3f531fd18233e92626d134a8b986175008c38;

            If20f8ce49f49f296f4747ef4388ed862862070b059bc482233542b99c18d7373 = Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa + ~I1a1149d160ca76d7b9db443f5095737e563a7b75de7375f9c148f4f4dbe7e7f0 + 1;
            I0a3f32d46730431a4e8b755f34e45c99a2498f70b0a1a72e30247dc78e20e944 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If20f8ce49f49f296f4747ef4388ed862862070b059bc482233542b99c18d7373);
            If56795023544f4a2942b0910b389ee77a220fffaf45786cb20c1806f3d76f76a    = I0a3f32d46730431a4e8b755f34e45c99a2498f70b0a1a72e30247dc78e20e944;

            Iac1ca36a507d9c411a740df9fea1934e7d8d64695834a37eecb2cde9d03a9204 = Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa + ~Ifdcd4016757d0cef222265289850476e0e2a6547732f999ca0cd8449f7134bbd + 1;
            I6ed20cd620c713a5aca6cc3a4b55daed825a10b3f9d779e6e83f4073130a5528 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iac1ca36a507d9c411a740df9fea1934e7d8d64695834a37eecb2cde9d03a9204);
            Ic9d92acd0f4cc0aa5cf4bc5a5f14bb848cb4267dd6aec78011f70039bf4f7c8c    = I6ed20cd620c713a5aca6cc3a4b55daed825a10b3f9d779e6e83f4073130a5528;

            Id62572be7c49640d6256571053ec24877befc584f4518c67f81dddd33afe02ee = Iaf213c4274d8c920cd0ce8713841466e62cd4583e81b3bdb7f45a84b58f425aa + ~I3eaa094e28f19bdbec184b0ba0f3792f90e67c77bd8dff9af6042c5002735505 + 1;
            I815ea11848fc8d4e5819cc19e041d9053b9f67a76ed786264b86c6d92c97464f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id62572be7c49640d6256571053ec24877befc584f4518c67f81dddd33afe02ee);
            I83b87ecce5b21302ac79a58afdd995b617634440666c2a50df5ba1868c7f81c2    = I815ea11848fc8d4e5819cc19e041d9053b9f67a76ed786264b86c6d92c97464f;

            I8c5856de3a047c2d8cd91175dd65f574230329e0a98bb369bc2f1efde176aef5 = I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 + ~Id9d184571e769ba27b0a5a10807ba8da3e6ba57ed7d66aad1cd984ddf5cbcbd0 + 1;
            Id78afeca7f85a7fd2eb3cbc54a726ab58c640d233f3b1f54a728f64ea1038fa2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8c5856de3a047c2d8cd91175dd65f574230329e0a98bb369bc2f1efde176aef5);
            Ida44179080ae7121a94fa6ddc8d15e57d73d73f15c2007f200eb205bd6c0c63f    = Id78afeca7f85a7fd2eb3cbc54a726ab58c640d233f3b1f54a728f64ea1038fa2;

            Ic3358b7d409c989b0359b4768845d172ff09d2c61bf9d17e51d0323a347dbbf5 = I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 + ~Ib43a705a217dd9f2321c3e61ee116d257d8ad59bff5b4f80435f9dd96a8d04fb + 1;
            I366b27c864334c4667735336cb00a70a99147206b5b080a90f7c73d36ff24f79 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic3358b7d409c989b0359b4768845d172ff09d2c61bf9d17e51d0323a347dbbf5);
            I0708b20a51af5c02051540c2de37aeeca5959bd958280e953a9cdf18c324d905    = I366b27c864334c4667735336cb00a70a99147206b5b080a90f7c73d36ff24f79;

            I4bae23c126c76b438684a2e720dd190ada836cd8aff3a9f217f8fc93dcb5941b = I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 + ~I800a86b8eeb247f39df85aba37dbaa93060858c235c6ac6b0912fca85af95477 + 1;
            I36793dfe7c63681d4c68b218eaed75db71f018b3b9a1902c95a586f9a040e60f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4bae23c126c76b438684a2e720dd190ada836cd8aff3a9f217f8fc93dcb5941b);
            I25510ca31a420de3078e0615a3a9f602e7a6f8698e6a79cb0d2688aa63f8e7cd    = I36793dfe7c63681d4c68b218eaed75db71f018b3b9a1902c95a586f9a040e60f;

            I1c6046860b8c1def57621b5c2fbdeb57b6bb9de1195675a875a1a028ea2cf881 = I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 + ~I0cc63aa921326ebb19427e9e06862cc0a42b375a328061bc7f6580bf3f1d3b12 + 1;
            I5f23f925a53b7246e36a09e80472df08b155e259db2d0ced8963692d36f85c84 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1c6046860b8c1def57621b5c2fbdeb57b6bb9de1195675a875a1a028ea2cf881);
            Ief493235efee1fdb4705ae4a1a0244c57346ff2b56b269552c6b5d64595056ca    = I5f23f925a53b7246e36a09e80472df08b155e259db2d0ced8963692d36f85c84;

            I6f58751fe0a0b377048b39ff9ed4d073ab5205a2ec8c36b93cf8adb44ad81d4f = I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 + ~I9beeb3f92470748db1e059cd6c5a929d1eee2a3ecd0ac097032c74f4134a22be + 1;
            I45bd49dc6c406523eda6bab5c72af5615d2a052f7f43502665d95c616383950c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6f58751fe0a0b377048b39ff9ed4d073ab5205a2ec8c36b93cf8adb44ad81d4f);
            I0a5ffd7c103836e4867f6819fab3096c582f2ce1db2c303bfebf50104b7d496b    = I45bd49dc6c406523eda6bab5c72af5615d2a052f7f43502665d95c616383950c;

            Ia43a684b6db0d7a69334ee35b6e06b35546b75cb48143fe9e7b54773b8c0341e = I584ad2d7fc1bd85a5181a996cbd2fdaa0edba05c6bd2b76336bd8b4307389d04 + ~I62b9322a1d5ff38480981e00d8469983588d084289f2f927f3339250b5c35985 + 1;
            I17013aa37e8e70e1e6cee9d90e8a3d4b07b1ff9122b2ad8c3b4c99deab9e6952 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia43a684b6db0d7a69334ee35b6e06b35546b75cb48143fe9e7b54773b8c0341e);
            Ife97a26fdf22e53aaf139436dd732d1fc8cd6cb4957269b6d0666495a0873c4f    = I17013aa37e8e70e1e6cee9d90e8a3d4b07b1ff9122b2ad8c3b4c99deab9e6952;

            I0d2a131e78e3e0c36dcc971e7ff76990cf1d19e2d90d373db2a81750458bfcc0 = I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5 + ~I62d2fe36d10e598efb7f38f4f57e4511d08c366d7df7f51bfbc63eaaf216035c + 1;
            I7506221ee4a6d544aac3f4da89b28ab6fa9d4ea68075210db51d8c6c0d486af0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0d2a131e78e3e0c36dcc971e7ff76990cf1d19e2d90d373db2a81750458bfcc0);
            I2bb55e3fbb0c342fd0434fbb00b85eae3c5f4075979e290f3d22673c392e3a60    = I7506221ee4a6d544aac3f4da89b28ab6fa9d4ea68075210db51d8c6c0d486af0;

            I7a190a23ac0ecbec7ef85c968ae10b90f7f0d9f5400aeb74109b51caf4caa2e0 = I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5 + ~I58aad5a5682b85bf58d67b9b00883f015e4093979fae9138f7dcd813618e26dd + 1;
            Ibc7ef4ff5d5e894f81ff8cd7b641624a6a898281185b77a1e2ecaa556312dba6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a190a23ac0ecbec7ef85c968ae10b90f7f0d9f5400aeb74109b51caf4caa2e0);
            I7dbeb05d89d3fea39368b48237973c682e796d24aba3438109147cc316b96ba2    = Ibc7ef4ff5d5e894f81ff8cd7b641624a6a898281185b77a1e2ecaa556312dba6;

            I97576b987f44843040444751f4b37c3b5974dfe60b4015dbac8adb962635ed1e = I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5 + ~I2f928325d150ab718f3b764d3fc4e15d88af5567b4554ef8bbd02f4c3984f544 + 1;
            I94f547c68a6f0daca7dd1152b5c9440fb76b34a3a133c8947cf8e1ec151cf3cc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I97576b987f44843040444751f4b37c3b5974dfe60b4015dbac8adb962635ed1e);
            I6e863b3eb7ba8e7ad90945ec76c695330de32ae32b69ae2a03091d1ef0142670    = I94f547c68a6f0daca7dd1152b5c9440fb76b34a3a133c8947cf8e1ec151cf3cc;

            Ib6bcf064fff2ac3dac1a636d200459bce8d2240757710aebf6f5ff055ba808b8 = I5ee55e7e31ad2837760ca081f8f37bdc76814d264ef9dfe6a5c2d691d73909e5 + ~I2af0f38cbf134ae07c76f06d4aafee537bcdfe91b1c4aff1ae27898e18da5113 + 1;
            I80b8de6095d16eb257b9da8adcb999d08ca7412d77b70d50bbf75ad9ceb0ee02 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib6bcf064fff2ac3dac1a636d200459bce8d2240757710aebf6f5ff055ba808b8);
            Ib13a4de6ca8fc3856fdeaa543ff8aae727f62ebff652acce5e23c6c121ee740a    = I80b8de6095d16eb257b9da8adcb999d08ca7412d77b70d50bbf75ad9ceb0ee02;

            Iad4f04d003ec15a32b36b0741a3fc3ee341e7d02d9b7d495d63e26d02d5f278c = Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3 + ~Ic0561c97824b9d5b0d84c33cd05cd4f95b9cacab06eeb5e022b0cecd043c6a75 + 1;
            Ife51a94dad3ebb020992018db5c1e1884eef8a8afa5487a3365594fdabcda2e6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iad4f04d003ec15a32b36b0741a3fc3ee341e7d02d9b7d495d63e26d02d5f278c);
            I22692863c63315b86c8a72a902c88573f4af6aa3b1691f68ed588a38ac77f7c2    = Ife51a94dad3ebb020992018db5c1e1884eef8a8afa5487a3365594fdabcda2e6;

            I71245defdd1d5a15a8c64a0c1bc585fb3a5acc2f6427408b4c526faf77e5668d = Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3 + ~I17e36eac60eec64de05cb738d1e6055086891ee6fd7d8fb300df4f98a3405276 + 1;
            I71fe587ddc1cfb6d7ddd3b8471786134d761d3987128e249992f460a0fabf1a3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I71245defdd1d5a15a8c64a0c1bc585fb3a5acc2f6427408b4c526faf77e5668d);
            I2f18a4d6ae6bbfa53e26a0aa169b1cd1c40ff544f7fd42b9ac493729ffa90ce3    = I71fe587ddc1cfb6d7ddd3b8471786134d761d3987128e249992f460a0fabf1a3;

            I9ce7dc815e30f744716169eabc1fd21116601a539776481e8f75ee17262c7fed = Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3 + ~I30b6c3fe760f221d2861a5b6061034f6dee7320a04cbd7de2a3c728427f927fa + 1;
            I693f23e6d443e1a19036a40851f82c92837e7bc1db7efa4913fd4f4354e88471 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9ce7dc815e30f744716169eabc1fd21116601a539776481e8f75ee17262c7fed);
            I5c4daf848487e7de6d8f95704179a300218ae460e56dbe71d33805739ea61144    = I693f23e6d443e1a19036a40851f82c92837e7bc1db7efa4913fd4f4354e88471;

            I19dd506a7468a183410e0bae3025af7af57306a264f0043f2f9a0635a3a5cb5e = Ife10d633dfbd29a354bd4fbea92cff68e41f4ee4df0bec9761e09394b3083ed3 + ~Iec6be5ba578c849ae0e4fee9c059ff88c36cfa7c14cfe218cad7f7f1d6744024 + 1;
            I43594a967fc4ae5970a0ea8821dc6b91e5de451cd6a5bee90fe8be18dd172caf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I19dd506a7468a183410e0bae3025af7af57306a264f0043f2f9a0635a3a5cb5e);
            I94386cfbe9c6f26a678c961cdb0f15d314fc3e6bd04edc61d5596107adc68969    = I43594a967fc4ae5970a0ea8821dc6b91e5de451cd6a5bee90fe8be18dd172caf;

            Idfc570f0db8ee7ca88a35b7c9ffc2306308ecc26877a75c31ccc436f1e9bdcc9 = I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf + ~Id7d51984757deb5794eccbf50647e7535041a18dc506aa16b4ba0ad36bc66b0c + 1;
            I62053bc27431d9b3e1615fbf5ede27d633603a9bbdde1e6df0eb795ad9a00d07 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idfc570f0db8ee7ca88a35b7c9ffc2306308ecc26877a75c31ccc436f1e9bdcc9);
            Icbf8ff1f03b79fbbdd3d73ba2d399ba98a814ca4db6f6541ce67d8e5558d0eb8    = I62053bc27431d9b3e1615fbf5ede27d633603a9bbdde1e6df0eb795ad9a00d07;

            I4e3b7e54b82af833886fdc3ffcb335189bfd516a758fd9fe96a0f4dbb919ed11 = I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf + ~I05782c612bec6ce9c2707bd6cb6efd55e1da4d234be502ac88cd02453c61ca60 + 1;
            I108b6619ec88853b35b010ac5ab6a5c649973073d8523fbe5503a6ce91a78534 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4e3b7e54b82af833886fdc3ffcb335189bfd516a758fd9fe96a0f4dbb919ed11);
            Ia69053f259b67f0fd728ca4fcd2bd39802adb86be01404890b17989eb74240db    = I108b6619ec88853b35b010ac5ab6a5c649973073d8523fbe5503a6ce91a78534;

            I92b84a136bf952296131c7162a68c4215e69d2cabfd345b29ac1c0bf22585921 = I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf + ~Ibc35679e4c52c119bb0ab5c5a485b11a4bd43ceba90f9998d9704d08ca3285f9 + 1;
            I719ca66a3b30047457c24a43119751ee15bd686df9a03f81885e3d8b2cbd07f8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I92b84a136bf952296131c7162a68c4215e69d2cabfd345b29ac1c0bf22585921);
            Id372f6f6b6b8b583699e8af0deba407a85b166caf3110f896594d222f0114cb8    = I719ca66a3b30047457c24a43119751ee15bd686df9a03f81885e3d8b2cbd07f8;

            I7203b0e25219256938283b8d39adec66610804f8024a63dd2bad2ca9e9e01a10 = I4cc7cb7dcabb05337b18279eb8b04e7d9ecbdd2166f70bf0570f1d8a9a281dcf + ~Id18c335cef6d5d988e55f6fda5a09a24ee80f4d4755f797a11ee94141b69b97d + 1;
            I9a9a7a98aafa77a8d0eac55b80e3c9a4dbc6b79d4a714c249193062b14ab5695 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7203b0e25219256938283b8d39adec66610804f8024a63dd2bad2ca9e9e01a10);
            Id9b0a59eec0b8ceb485b7dafbff07051b5bd44c8b9ee4c3fda3773cef4450e78    = I9a9a7a98aafa77a8d0eac55b80e3c9a4dbc6b79d4a714c249193062b14ab5695;

            I8d5085a98240b391006667ecdde09a3735f02bebf47c3ae2e3f4983183111e5e = If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d + ~I272bc7cf289752b36b9811d4ec63f5c17cb40399f39607b00ba51817fad59e1b + 1;
            Ifaa8161798b18d4d55533a337ff4bbfcba6a94e4f92c99d728f1b9e0a9afd72e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8d5085a98240b391006667ecdde09a3735f02bebf47c3ae2e3f4983183111e5e);
            Ic0563f05659ac941778904304c02575d9c9f2125ee05515ffd05749e20880d90    = Ifaa8161798b18d4d55533a337ff4bbfcba6a94e4f92c99d728f1b9e0a9afd72e;

            I793fbfdab6a3b0b8951196e0a8a76d4844094cb64802cd8d50bc2b7ffbb0d937 = If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d + ~I343c495ca033301298c16cbb81a11a7f9d50dfa8b93ea9226caa182c6fae8737 + 1;
            Ic2f50a4dad9dc0ec10f13868d7a117a26e43b501da77693b309eee3c9c713b1f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I793fbfdab6a3b0b8951196e0a8a76d4844094cb64802cd8d50bc2b7ffbb0d937);
            I81590f464fadabf1667af046de2f41172c36389854de1ad410e32cbe3b719ced    = Ic2f50a4dad9dc0ec10f13868d7a117a26e43b501da77693b309eee3c9c713b1f;

            I62a85956a9fd75b6c1d7f93f5472394fc8d0413995f21a8eab042ec0268e63fc = If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d + ~I4d6d60296569a9b2a811f8064057743f13fdc60379669472d28df97061ccedb0 + 1;
            I92edc25de8e424524b27a64e0970c549d2ee4d232fea857eeb0b9a391fd8a03c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I62a85956a9fd75b6c1d7f93f5472394fc8d0413995f21a8eab042ec0268e63fc);
            Ib2f85bbcac9533694e4da81d1e86313ed14510ac8a37929a6158c888ba9cdb0c    = I92edc25de8e424524b27a64e0970c549d2ee4d232fea857eeb0b9a391fd8a03c;

            I64a047649ca6b299cf603e326db494b30d1eb35725319f172957fa38f00150ca = If3aaf64e865cb485a895082261633ea187493e19d6ab0ef8d2aa24bf655dd39d + ~Ie85ad3f88a177d67b69eb3a03e4a9d92f7431af9de9ccd06f2caa01f9d144f33 + 1;
            I09572043800626670079ecc4ff74ee7ff644d70879ed7598d124a0d5e847b288 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I64a047649ca6b299cf603e326db494b30d1eb35725319f172957fa38f00150ca);
            I6128d022628a70641f03bc8d1508dc00be5665cbb426ab6b2befa774ad124efc    = I09572043800626670079ecc4ff74ee7ff644d70879ed7598d124a0d5e847b288;

            I1da8e393ff7564ba162ca784da6731a8632fc4f6b34d907a52185a8b6a59a2d0 = Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde + ~Ib8956dcf80473ed75d04e9fcc74400f54ee0b840fce7500bcd68ea6dac6d4473 + 1;
            I4b3e88dd84be91d43898b83141459d2ecaa7f53424793691b357a4153fbe885c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1da8e393ff7564ba162ca784da6731a8632fc4f6b34d907a52185a8b6a59a2d0);
            I9eb8c67587f031f7dd6668286278ec62c632eebd218d4b5fca188e6447de8cff    = I4b3e88dd84be91d43898b83141459d2ecaa7f53424793691b357a4153fbe885c;

            Ib1c9e95f283090d633d1a8deac1211672e46383b70ec08ba60820f0096fea280 = Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde + ~I57ae0fac4bc1fada55e48ef9952dd7b81a55414196fc22fb27a20b723832aa84 + 1;
            Ia5947b18a468bba37f977f0c09103b82cda7962015feff03f0f7259f29d77d3b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib1c9e95f283090d633d1a8deac1211672e46383b70ec08ba60820f0096fea280);
            I930d8c08531d026f47ecb265d741cbd6a41286e3898d547ec9770fe114da36a2    = Ia5947b18a468bba37f977f0c09103b82cda7962015feff03f0f7259f29d77d3b;

            I066d165e686a647ec05e381773c53d7bd83320b8abd57693dc5dae88a01fd8b6 = Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde + ~I1a54a485e54cb6d528feed952641c7e5350f3d386ceb62ddd2778ad179aef345 + 1;
            I8e2ad7d4039c25bbd7c09ac2d55efdb8a8660f4949c64c3ddc3729f253ffd9f3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I066d165e686a647ec05e381773c53d7bd83320b8abd57693dc5dae88a01fd8b6);
            I7401c9a97f13630805f89ca9767771302df865505689963bf68db913a151a1bd    = I8e2ad7d4039c25bbd7c09ac2d55efdb8a8660f4949c64c3ddc3729f253ffd9f3;

            Iba95ca83f9a8247abda33f9ae9bafedf0b26e6616d5bfbfd78b02637f6120c00 = Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde + ~Ideafcce97c26d412480370ab40d8261f37e8bf0ba68bf7d04f4099a517195dfa + 1;
            Ibf297726d3ad1a4e50327cce6585b2b5449e95ba1c222311ce9d2fa03c74dd88 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iba95ca83f9a8247abda33f9ae9bafedf0b26e6616d5bfbfd78b02637f6120c00);
            I0533ded3a5c68b582fb4785c33ad5742da4947c904b1a52e05c80a3645f3fef1    = Ibf297726d3ad1a4e50327cce6585b2b5449e95ba1c222311ce9d2fa03c74dd88;

            Ie4936469b1efc82d537631d9126581b917e052838c19db1f8fb4512d7352f6d6 = Id896477101c7d097a577e8a8ad1ef2acacf6b3ede1693101688869982e9bdcde + ~I53e788aafc97015db67a8363c91d81d369d80c4d24542fa45faf7833fa4189c1 + 1;
            I2118c0ebdd9baa8fcfd921632fb1fc58d995fc55e506507087ed673f52693ec0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie4936469b1efc82d537631d9126581b917e052838c19db1f8fb4512d7352f6d6);
            I2616f37126555e344d3b2f904a46af3f8a5fcfd59fcbf0677377f16cd59f3be5    = I2118c0ebdd9baa8fcfd921632fb1fc58d995fc55e506507087ed673f52693ec0;

            I7dae66792f1ba5fc8ff7d7541e3c9fdc44b001e3103715d98c57ddbd35686d37 = Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 + ~I0549cd0fd3abf1658d503a09b0baa63d09b1411eaa524e56fd30b12f8498e549 + 1;
            Ica997f542c175790baa0650ff204f09e387d1e1119096ae7f1bf9b6a683c6b80 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7dae66792f1ba5fc8ff7d7541e3c9fdc44b001e3103715d98c57ddbd35686d37);
            Ia049b06c7b1e457c3ee5643e87fc729a409f2fa943275ce5dda083fb1253c2eb    = Ica997f542c175790baa0650ff204f09e387d1e1119096ae7f1bf9b6a683c6b80;

            Idb01042afb3fe35b5df33f4a990e8d512975c238b7dc146f8c60fe42178a232e = Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 + ~I23f5e95dbae4b1223d603061df9b75b9a9ae8409c6bc4ad1fe23d3f5c7a68bb1 + 1;
            I49b78fc64683b38b3318a903923a2523aa1fd7e2f3e13bfb26709a93fd8ed772 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idb01042afb3fe35b5df33f4a990e8d512975c238b7dc146f8c60fe42178a232e);
            I6d785370057273f67048d3cda9ebfb0c8bc43fc5f34af47935e45302ed66e021    = I49b78fc64683b38b3318a903923a2523aa1fd7e2f3e13bfb26709a93fd8ed772;

            I81b03c11c47391653037bfc546e4abce946e244fe10d6d3746006dbecc9e6dc9 = Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 + ~I4df045f8dab91c2eee20a03bcbea586a003659b77d8a6e941bd2b2ead3006d04 + 1;
            I2965e4d3241186a43f93eeb83b4ec8d7e25faf3502c42556448bcca049d1add7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I81b03c11c47391653037bfc546e4abce946e244fe10d6d3746006dbecc9e6dc9);
            If668ac9edc8047d257ed4f162d07f8f326c0c3ffed244595bc249275f04f02b0    = I2965e4d3241186a43f93eeb83b4ec8d7e25faf3502c42556448bcca049d1add7;

            I44dc65b9b972b02070e5bac23ee64e568adb39d61d0f3ddbac27ad0abf453fde = Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 + ~I8a5d6a4832abe68ab6e9ae33b1b6026805c5db0d186df37fe623a2d9931b2534 + 1;
            I883f00e2f9f6d78ae17d150f6305fed3e16ab0da7c8b4ccea0b9aae62672cce8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I44dc65b9b972b02070e5bac23ee64e568adb39d61d0f3ddbac27ad0abf453fde);
            I8ecda1185b64bb196b1281095a7e3bf01377e6fbc7ec9cb20a3700f458944fa9    = I883f00e2f9f6d78ae17d150f6305fed3e16ab0da7c8b4ccea0b9aae62672cce8;

            I53ea37aef026e5dc7e966fab827b86b9a180b1c64d53801e51d7f2c66c729cf1 = Iffe93e6135842606d7819a94e14e0547e0ea97d65ce7caf250097684e7cc9d27 + ~I8f74cd611f5df70ef183e9d4a86b5ac23349be8cb99cd470c596fcaa6ec95248 + 1;
            I4611a21e5c71e60d5cbf9d62950215aee3679907ef0c908ba375182103b06375 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I53ea37aef026e5dc7e966fab827b86b9a180b1c64d53801e51d7f2c66c729cf1);
            I4b6ef863f3c19600f1325225dfeba21b5e9333dff55ddcf9f0cd8e8ec3581a32    = I4611a21e5c71e60d5cbf9d62950215aee3679907ef0c908ba375182103b06375;

            I7147ae9d3a1f4fda281c89a81e01b66d9db82d9e8f609e313a374cd5aaadd687 = I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 + ~I451de528c384521cbb78ae32b3d4640b0cb8d507c10e11ff59a74a9caadd2117 + 1;
            I58f661e6c3018394127a3cf6fb03e6993ca641adb970d8a7c0c2fe2547a36c94 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7147ae9d3a1f4fda281c89a81e01b66d9db82d9e8f609e313a374cd5aaadd687);
            I2cfed4bfd244233c8d85a9ebd9edd2c03f3bbbeddb7c7a32de444794e9c44e17    = I58f661e6c3018394127a3cf6fb03e6993ca641adb970d8a7c0c2fe2547a36c94;

            I550a8278e2a551834175e8275532965c7204bd2f4d021e0c087eedd5a3fbef93 = I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 + ~I72329ad9fd98258074b92a7e88a88c68f8db57e7d6460e9c29ec7f3cc251de29 + 1;
            I0a660d35184450970491123819f2a1ac18ae2eb7132339cd57e564cff1dceac4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I550a8278e2a551834175e8275532965c7204bd2f4d021e0c087eedd5a3fbef93);
            If7e91102c5105c0ecfc871fce4bfb86900fbfc837d6f06f3229d362d20e51ae0    = I0a660d35184450970491123819f2a1ac18ae2eb7132339cd57e564cff1dceac4;

            If5b5d22613b68a9bad72ca89d654b0a7f9d21914b3d596af6ef7de32b98e66e9 = I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 + ~I1edf83d193e0825c58f470cb0d4ccd85e3df4652ab68fe3a701a6ee0e8a0658a + 1;
            I93aaae3307747b620bdc3ad1ef6bd872c1b4fa81e99664494ff00b4357f1675f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If5b5d22613b68a9bad72ca89d654b0a7f9d21914b3d596af6ef7de32b98e66e9);
            I7643b1d4690f708c2c0d93adf0c5ac9ef99fe85eedc024e505edc74208d0f94f    = I93aaae3307747b620bdc3ad1ef6bd872c1b4fa81e99664494ff00b4357f1675f;

            I749908d9a05ab10736825bc8f1db4b879d94c4cdb920daa9aec231b8b2a26dbd = I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 + ~I67e66b155579d855e0c14e91d2ce1fc6fe1d2f869e4f56b37de5f700d84073fe + 1;
            I1efa5f2029f0dba2f9a46aeafb6ad51afc192458717939428f80359d159e00f1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I749908d9a05ab10736825bc8f1db4b879d94c4cdb920daa9aec231b8b2a26dbd);
            I78f713264010c545a0147149b2fa2efaa92985405649e4c4313a0832e8222787    = I1efa5f2029f0dba2f9a46aeafb6ad51afc192458717939428f80359d159e00f1;

            Id85f8d61522c12b51ada0a5c2f8c492d1a72c4d5ef88c99b2b5ca0c8a885aed8 = I9b0c37ae8193193043c4ccebd0e160646dc9623e2f558e8c6d884c6c1cf2cbd1 + ~Ief3910aa326e0d9782566c81ab1cbd09faf46d3552f78d7ef5fc9de1d9c245d6 + 1;
            Ib4e74743b49becf72add5b8e28261cfde3acda86de12ad6d7ee855668c1c79f8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id85f8d61522c12b51ada0a5c2f8c492d1a72c4d5ef88c99b2b5ca0c8a885aed8);
            I6fc297df8d4527160ce05230a017f3710f7c026c6b11d64babe81959156f3462    = Ib4e74743b49becf72add5b8e28261cfde3acda86de12ad6d7ee855668c1c79f8;

            I7a627bb2c8162e911b06414d590ddfb19a4b1b84d0af6c65f451bcb6cb4978e1 = I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b + ~I511b38f7ea620301cc3bfa759ab56a2dac9061fc83fb1281673a6cf276abcabf + 1;
            I8aed9a4d4cda2feddfa8b481712f5723cd792e834384343bede45a150ec1b12e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a627bb2c8162e911b06414d590ddfb19a4b1b84d0af6c65f451bcb6cb4978e1);
            Ie3e13531d22eb604e4a351dce5ee5512894170b3dd6f87962756c534438688ea    = I8aed9a4d4cda2feddfa8b481712f5723cd792e834384343bede45a150ec1b12e;

            Ica888e39630b6f3eb799326d4046056ef55883125634fcbdf6c36133ba571b52 = I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b + ~I61e7244c25e176443b24d592ff4299482d572c1705c3e0a6b44698b5366ea3ff + 1;
            If5f5d06e01de5ae4ba52dc9f61ddb507f1e34bdd36dceca20c19df859460eda6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ica888e39630b6f3eb799326d4046056ef55883125634fcbdf6c36133ba571b52);
            I10312c661b621655f99ef4c729f81bfd1c6aabf28b2f3372264d69d6d177d475    = If5f5d06e01de5ae4ba52dc9f61ddb507f1e34bdd36dceca20c19df859460eda6;

            I7e0846788926a4b2a76f01957b236d542f43fb90aafc16a952cc502d83f31cd9 = I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b + ~I1d5563063ac8386b450a3a36bb3d0a3586cfd6d11471071685e3f7f897d8eff2 + 1;
            Ia1f7010c7618800ab0201f331741ab58055c31cd72fdd0e3db900aa455703ad0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7e0846788926a4b2a76f01957b236d542f43fb90aafc16a952cc502d83f31cd9);
            Ic4b994b93547d46c87ce7cd1fff323144f9de0ff6e79ef0ce9ecc1db89340e6b    = Ia1f7010c7618800ab0201f331741ab58055c31cd72fdd0e3db900aa455703ad0;

            I85ff081ed2d76aa65ad78d86b7804ea0f8822cd35f8b14612104ec232184c5fb = I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b + ~I0c92cee9eb9e3c8300210834a106174a25005d9a468a481e0f594a960b5995ab + 1;
            Idba5ae25e3ea830381b3dadc351ea69d0e7b2bae1370ecc24dec6d408e7f0e3a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I85ff081ed2d76aa65ad78d86b7804ea0f8822cd35f8b14612104ec232184c5fb);
            I38340f75bcbf775a9e070a528d926355b818091cd8e5c1792450d2713ae436bc    = Idba5ae25e3ea830381b3dadc351ea69d0e7b2bae1370ecc24dec6d408e7f0e3a;

            I2f5cf926d3a647e02544e7839c6e999a0798aa5c810a6031433237932e96602e = I7d038b06bf898a198e97664a3c65a8a947c88a97805c330ba7e2c21dc692200b + ~Idddd98e139a087c7aef3922ea2542dd364c9d30f70665754f751ed88dfbd3701 + 1;
            Icc06285b311fcba47b9670c971839fa401cb4c74f3da347961786337621bc629 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2f5cf926d3a647e02544e7839c6e999a0798aa5c810a6031433237932e96602e);
            Iad0e03f141449cf08d3cfdfcd976e4b5a8401179533f5aa4f8216198b749a4e1    = Icc06285b311fcba47b9670c971839fa401cb4c74f3da347961786337621bc629;

            I5f43984a17fec9b995aac537cfed942b8c61fcb134ba29fc82a41db44d46c820 = Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e + ~I533b2cd0b272eac7c3f9005cc355cf85ce73803134a0fe0ec194628c3af0ed91 + 1;
            I4332a72ae402f4043459e290fc47700a896e6eef5e383e720847ff34ef1cb150 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5f43984a17fec9b995aac537cfed942b8c61fcb134ba29fc82a41db44d46c820);
            Ibc82061cbb8fc5b88d39b5b714381ff331de2b2877376cb96a32d6742f3cac6d    = I4332a72ae402f4043459e290fc47700a896e6eef5e383e720847ff34ef1cb150;

            I7a97a4296eda318163fa6fe4417e08ad1963bb488a6bac31f3b3b6af9e7ab213 = Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e + ~Ieca82bcdc6bd68dc2a28a3b203d8adaa09f89fbf0df6cacd8656b54b141d758a + 1;
            I937131c2de1f55c3990b577d63b44282462abde126ef6a5fbe5ea962d48479e8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a97a4296eda318163fa6fe4417e08ad1963bb488a6bac31f3b3b6af9e7ab213);
            I49af7bf73e330c26c437d8f0447a930c63d4677498d07a28ff9b2b25860258d0    = I937131c2de1f55c3990b577d63b44282462abde126ef6a5fbe5ea962d48479e8;

            I439b2964d8e94fafab2d3cd19e72728d4e763624497e8f44e10a8be796d87a31 = Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e + ~I207af234897ed272d784f4a9f8850eaaa2fbf47f583ed1f0564201e33dccfb66 + 1;
            I83e04a31ba3a09afcd0f223722c2852e314c79d93374a673cfd952bbe94fa816 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I439b2964d8e94fafab2d3cd19e72728d4e763624497e8f44e10a8be796d87a31);
            I5e977efb6007fb448a0cd05362289e5bbace24ff868e4fb623ba54135e53fc82    = I83e04a31ba3a09afcd0f223722c2852e314c79d93374a673cfd952bbe94fa816;

            I6476bbdf545c28c272dffa9640a8a640802826f625e7963386bd6b5309fb3588 = Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e + ~Ic336cf50b44edc74db080d1127ba09a4313c0972702200ac5207aae8ce6b1062 + 1;
            I7258f6d3dbef6e7ae01af1761728fc7b034158f1e7f26b13b21b500e1bf3e189 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6476bbdf545c28c272dffa9640a8a640802826f625e7963386bd6b5309fb3588);
            I98233f63b47681b1d8b5e3decd1ab8ad783734a17e2b27c88234f00b23fa30cb    = I7258f6d3dbef6e7ae01af1761728fc7b034158f1e7f26b13b21b500e1bf3e189;

            Ie4122a78fa86e3e8cc54ebd8e3d1433ab29af18f8d6683a4eceefb4108faeb0a = Ia5da5cf90f0aac9fe15ea133d2ddf64297ddc7b8eb6532c6522231e71ada8d7e + ~I474f7c67e6159d041be6d6f4f96fe58f9b7086757936ebbc86340bcd9cd9962c + 1;
            I3d284053eea1d128eb2703e23589b78e03e04e2b5219696ee3b70b3645c0267c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie4122a78fa86e3e8cc54ebd8e3d1433ab29af18f8d6683a4eceefb4108faeb0a);
            I58660674a5ad4c7022a05e5cfcd03fdc7161e65e8050cc59ae6fefc404b6b310    = I3d284053eea1d128eb2703e23589b78e03e04e2b5219696ee3b70b3645c0267c;

            I1de838959290a975e08aae4a25944f707aa1ed044defb47058acac42075cb7ac = Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 + ~Ib8b4f3fbd26b51974ecee1565c3d0c8fa7abd94e467a7369a62ceafa7ea5ddaf + 1;
            Ia14eb5936f779af58b044db01b8d6d6f89557eaa5deb1b16ddc8f7400351b6de = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1de838959290a975e08aae4a25944f707aa1ed044defb47058acac42075cb7ac);
            I9612c348b28222bc7559977c8bd902d73267c977bfbe179506c88be746830331    = Ia14eb5936f779af58b044db01b8d6d6f89557eaa5deb1b16ddc8f7400351b6de;

            I5175fc2784d1f63752e69a808f26af8fddf78fb8ab1a897fbda883f056debdb3 = Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 + ~I0b2c4982c217189306b4f5d3bace84daaa25f2bcd089f5de092f9a7900106c6c + 1;
            I7a3f69cd5191d002a2b8428d09a32b0572981dfa535a5fe1d4406ff3c5193797 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5175fc2784d1f63752e69a808f26af8fddf78fb8ab1a897fbda883f056debdb3);
            Ifea5f415406637bbe581d11e57aaab23cecc2dc1957f45152f03d3006334d24c    = I7a3f69cd5191d002a2b8428d09a32b0572981dfa535a5fe1d4406ff3c5193797;

            I4056a6197e1723e278afa54ba45c2bcaa2766665f2d405d7f11217213f4af9bd = Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 + ~Icc13ce9fe63ee1c11fd5dddbf0a294cf6ab7ae703f742a92150b7a77868a5a16 + 1;
            I1a2e691f96157814ff15983f1dc0c522dfeccac15ebe1fa25bcacaa461170b15 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4056a6197e1723e278afa54ba45c2bcaa2766665f2d405d7f11217213f4af9bd);
            Ie56c2e96de8be01add59d3005f52661524c2193f6bd0fae2a759d4afe9607388    = I1a2e691f96157814ff15983f1dc0c522dfeccac15ebe1fa25bcacaa461170b15;

            I913a4d3bc811c985c378f0c3ceb8cc0d03637df817266b2a5009fe4e96362cc8 = Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 + ~I91e90d84eae561663a2e9e59f79782a78095807b98187add5501500b8c1cb126 + 1;
            Ifef7ad6de75a930ef9a0fd7a22e35afa498ad3ae74dbf41596b9bd952bb82be2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I913a4d3bc811c985c378f0c3ceb8cc0d03637df817266b2a5009fe4e96362cc8);
            I1744ca88c13acb5d2afa42ffe0ee5823eab5e32cbcf3248db4faffd6fe9e2537    = Ifef7ad6de75a930ef9a0fd7a22e35afa498ad3ae74dbf41596b9bd952bb82be2;

            I594b5684b4713ef793ee902ece02cf083e909b95354d67c351748b2b1ee2599d = Ib13c2a56bb6a431fb040a58ae8bcaabb17df8e31d2c45bfff7d9add874119985 + ~I2a1c16f7d4c3261619c325f4b5cfe98993d5957a2ff466bae11c9cec6006cac6 + 1;
            I680a7b47f68662a83f4298c9110d5e5a04eb459ef379b69a53e7f90d371084a9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I594b5684b4713ef793ee902ece02cf083e909b95354d67c351748b2b1ee2599d);
            I2646e32dd3a69da746d970611fa0a89f96286df22ebdcef1ab746d70c4db4331    = I680a7b47f68662a83f4298c9110d5e5a04eb459ef379b69a53e7f90d371084a9;

            I84f3d2170c4ac381738a10ae95bcb1a102d86d6c96bc9c0eef4a682237cc96fa = Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 + ~Iff259e6b8d77d06a8354c4d1662328284ede633f1ca4ec4731dcdae94e869f66 + 1;
            I343f02bd7da57ace84d1a265307da810c9ef6a56ada6ca3f1e102c8e4d53d89f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I84f3d2170c4ac381738a10ae95bcb1a102d86d6c96bc9c0eef4a682237cc96fa);
            I4c7da80c76f8d8ad9ed1199810aaa919460f955b2745ae54cdea9276ad5e2491    = I343f02bd7da57ace84d1a265307da810c9ef6a56ada6ca3f1e102c8e4d53d89f;

            I386f960be90b491237062d67c19264f36bff56381c3264cd7942a395bba04e72 = Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 + ~I873ab672a8d92c69b75cd8e627aaec129f1cd371c9f863a6bf88e3965909a6d6 + 1;
            I83858f36d2e66e2bb6f4357e978909888d598c4ae084d87a74d06f3ab7c334c5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I386f960be90b491237062d67c19264f36bff56381c3264cd7942a395bba04e72);
            I1e411a908fa94c50629647023bf56aaf275299c8c49933fe67ccf00d3ed68d7b    = I83858f36d2e66e2bb6f4357e978909888d598c4ae084d87a74d06f3ab7c334c5;

            Id25989c592a2848f8881f1ea00c42faaaf70c1571f602311ff1bad99c7cd151c = Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 + ~I062483fac022c2d74cc4bb84d57c636a3bbb67d68dacf0da453e3b5f71ff8846 + 1;
            If9bcfc0a82ffb81925d5e0fb3b8bd0ebd910b079c271c352751e38dbe327f634 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id25989c592a2848f8881f1ea00c42faaaf70c1571f602311ff1bad99c7cd151c);
            Ia06978f4049096a298ffcdf526e89060e8f27418076fa351962ec6f407576753    = If9bcfc0a82ffb81925d5e0fb3b8bd0ebd910b079c271c352751e38dbe327f634;

            Ie224e49b46cb25ecb4a8126eaf672bb12181bb28cb1e7cec7eccc94403d72b09 = Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 + ~If4b0b6bcc29aecf6816eab93edb0cb358730913253ae72d15db63ae06b19c52a + 1;
            Ie08a9d45e117e5fad39310981ed379f876f4330ccc7674752b26bfd2547adcac = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie224e49b46cb25ecb4a8126eaf672bb12181bb28cb1e7cec7eccc94403d72b09);
            I93695abbc93c5e195bbc5a1fee05aa7ceb4c58b273ed67ec6f28538aef0843e4    = Ie08a9d45e117e5fad39310981ed379f876f4330ccc7674752b26bfd2547adcac;

            I4e51e76c5c70e114f648c8715d629503228ea3845a66122c7da381e67e805912 = Ia5b00f703869d540a014c7928a5221f0b022584d8ae5c8302f57f654bfc6e936 + ~I881a2d7025d422202455bdff165dd982c2f4953b361f29688e75ccdf9e04d476 + 1;
            Ice7416e3625bcb882a0caa84958b2d20b2a6901ef7a7c748ada330c86ea41763 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4e51e76c5c70e114f648c8715d629503228ea3845a66122c7da381e67e805912);
            I81b17367c5766001911129ae2370c1dc7b3509565fe78fa6e552b7ef936da360    = Ice7416e3625bcb882a0caa84958b2d20b2a6901ef7a7c748ada330c86ea41763;

            I0261480422708e60435782d1ca5012495ec5345a3decbbc9815bbdc2ac374b42 = Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 + ~Iec33764f14e5b0a736fa76a2313325240a520c065b59c6cdd0f2fc5dc36a975b + 1;
            Iba6cd77ac5adf667b7d229aeec4f15eb6112ab90e4b51c09bcd7c64912cbdeb7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0261480422708e60435782d1ca5012495ec5345a3decbbc9815bbdc2ac374b42);
            I189d5a40f26a8b2893b53242a4ec7613797831a4a2192289df09283c7da753d8    = Iba6cd77ac5adf667b7d229aeec4f15eb6112ab90e4b51c09bcd7c64912cbdeb7;

            I4c4a1c399094746d92937b66958c6695428a7963aa82fef3c8cad424289612c5 = Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 + ~I19123fb30bb6e02a13f39e3e96af227e63abb1351e53cbb91b8d9a79be96053f + 1;
            Ib6cd4feec46af9df7727d5febf22dfe6059c43712e65fc7d982d1a6bcfeeba61 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4c4a1c399094746d92937b66958c6695428a7963aa82fef3c8cad424289612c5);
            I15429bf02bcaf6ac17ed02efb1e65c5c37254aedb9ef6181c2731c3f7e2a829d    = Ib6cd4feec46af9df7727d5febf22dfe6059c43712e65fc7d982d1a6bcfeeba61;

            Ic8f4e82cc2d1d643e87ce3d6da690336e97a779fb6fec983608492c39054b09b = Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 + ~Icb88d7eda8505d92744b075a1c229e3c0f6a9ff062bf5cd35f6f84467b451e9c + 1;
            I65b7c3c6e73e0f305942123f4ce97d6765b7bf86e61a3388774c36aabda5a491 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic8f4e82cc2d1d643e87ce3d6da690336e97a779fb6fec983608492c39054b09b);
            I1807ee521c06cb799faa136864a31c00869398289b0e3b185e702f42cb0e7412    = I65b7c3c6e73e0f305942123f4ce97d6765b7bf86e61a3388774c36aabda5a491;

            I3ecbc44de1811b06b96aedafb731823325898269d3f4d57a164b63cede9bee6a = Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 + ~I48ffe541268d63545fa48263d8df3c288af7b2646b4dca546a4dc521aa247651 + 1;
            I3525fe2422d10480b4caa9b5a6fda0228ffa3bcef28a2592f1eda3194cf30bc5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3ecbc44de1811b06b96aedafb731823325898269d3f4d57a164b63cede9bee6a);
            Id4ff3dcea8b6c38c5288cac263296941b841255967f2f58fa97a49fadb2fd2c8    = I3525fe2422d10480b4caa9b5a6fda0228ffa3bcef28a2592f1eda3194cf30bc5;

            Ib23e10fc2319b575483f38a9a75d9a8b55d394fe0d356c89478844a16504cfe5 = Ibeb8a30cdc03c850c2aedb9de445f49a9f429b2babb33e2fd637c9e9d270e634 + ~I8245c1ad016aa3d7290e1097eb966b09c8a38fa5bf62bcb7ef179f448104f47d + 1;
            Id78e42777220c16c860f907907256a6b28e2c5bb9cd011c71943ada87d30a9a2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib23e10fc2319b575483f38a9a75d9a8b55d394fe0d356c89478844a16504cfe5);
            I3856054a7ed02c524f8816bd8ba22a48935b393ced40e98c693416364ff512b3    = Id78e42777220c16c860f907907256a6b28e2c5bb9cd011c71943ada87d30a9a2;

            I5e6f080405681748ecd82a9b555257d553cc1dfcde4ac5f470bf1d282086b3d0 = Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 + ~Ie282d05ceadb0d075cca024b7311a5e477e903295d7928735a3c338287734846 + 1;
            I9c427f570b0c040928fa6aa62250920306e19e3031494e8933e30766f0c782a1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5e6f080405681748ecd82a9b555257d553cc1dfcde4ac5f470bf1d282086b3d0);
            I358ca9d90eebc0e19c434a7d1070a69b3c20b4f8152adcc45c0b73e8cf2c9902    = I9c427f570b0c040928fa6aa62250920306e19e3031494e8933e30766f0c782a1;

            Ia50f5ef4c28fc1650d46ad29de2ca34971e271c9248f06f24953db1d9f767faf = Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 + ~Ia81ab6d41925460c11303075dea72c7fb3fe533d88450c32414823fc5b10bfaa + 1;
            Id55c37de3455c6ed8da5c25f25a98b0ced5787638a4ac262c1bca6fafab7240d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia50f5ef4c28fc1650d46ad29de2ca34971e271c9248f06f24953db1d9f767faf);
            I1e60aaae452f97c016f3f3929c33637509d02988bea72048f7901a440232a85a    = Id55c37de3455c6ed8da5c25f25a98b0ced5787638a4ac262c1bca6fafab7240d;

            I3bd09d09f4fc3bb758f3c1f36925e9f0504fa342b2d80ee031e4c9665fd4ea90 = Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 + ~I1ca12951f309a25752defa88fa366a90a13ce83b7fb40610c01a8c11a3c2e59d + 1;
            If7049605331e013c95aa5eae16577637a3e8c80f5e4c325675654dcbbed1b613 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3bd09d09f4fc3bb758f3c1f36925e9f0504fa342b2d80ee031e4c9665fd4ea90);
            I312753748b2d173f2dde21bfad8dcf880f5fae94cd73fea4dbedb01c43c99b43    = If7049605331e013c95aa5eae16577637a3e8c80f5e4c325675654dcbbed1b613;

            Ie6ffb8ef3481ecbbf20e52ff7d04f51a024049190a3aa838c398f71bf1862115 = Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 + ~If2f521cf64a5e19b1f744d41d929a37a37689534d0e564224b128866d853b043 + 1;
            Idb9c4b9e280f7dd8b4c34242a9e58352a23799e10c7abf9c3448e8a28af55e33 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie6ffb8ef3481ecbbf20e52ff7d04f51a024049190a3aa838c398f71bf1862115);
            I6f210ff43165afc5b4c3a9a22dab74940c409a5fbdf9c47b9eaa68fa08918f23    = Idb9c4b9e280f7dd8b4c34242a9e58352a23799e10c7abf9c3448e8a28af55e33;

            I7a6117b4c4c11077b066e21819d7bc164de5f4060d1c12f57a9751afbc6fa59f = Iae2aefacb9712b5a39ba0e4d88dd2191edfe8af27b1e2048a444572faf4bc873 + ~I10206e80304f6e623a256b6042ceca13c691a34ef5b6d67667ab4bb11f0b0087 + 1;
            If3f33ea5e4ff428c3f59701f77e6f288293231923203fdc140d147d7ec769295 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a6117b4c4c11077b066e21819d7bc164de5f4060d1c12f57a9751afbc6fa59f);
            I3422d7c29697052f1d70152dce7d92858081099a7bd19bcb2a48add3d660ef12    = If3f33ea5e4ff428c3f59701f77e6f288293231923203fdc140d147d7ec769295;

            I96bf467638c2ab6963f57f29caf1efcda6250dad69e87b2833c6d094112a6731 = I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 + ~If787a878ae1cab622e44a13190d301d15d0c7ed9271dc50e997c926071f1cd02 + 1;
            Ieee64ec5ee871ab61afdf8c73149bb2fa68fcdc0050d80179dd9645b4f14a201 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I96bf467638c2ab6963f57f29caf1efcda6250dad69e87b2833c6d094112a6731);
            I90ed9972249e176fb13ac19818b591acc7f7048588409d394fbbb79ac26b3519    = Ieee64ec5ee871ab61afdf8c73149bb2fa68fcdc0050d80179dd9645b4f14a201;

            I6a9adf149ec3e5da62c6f86b4263910048b212f13e52e6b680386feaab5126f1 = I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 + ~I19b5f6ad3c2f2551b49883fbab077c8e3d76392fa42a5030b1f832917bc2641b + 1;
            I8cab52d76008f7803024c4d66307e41aa48256ae1e9d364c354b4b3e405e5c8a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6a9adf149ec3e5da62c6f86b4263910048b212f13e52e6b680386feaab5126f1);
            Iee565a93d37ce096492969d59077dd347ffeabe00c447298bd22adb6f66926dc    = I8cab52d76008f7803024c4d66307e41aa48256ae1e9d364c354b4b3e405e5c8a;

            Ie8947b0e08f05ed4ed4888467fd64bbdacfd30fcadb77185a75e53a60bb78877 = I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 + ~I1fd78c97c2a03a51b8d2a3dce2a553514aaeffdc051bfd3820d409da4b8189a0 + 1;
            I7acd9d954e3db160301869bcb6aedd5652613816ae8340f271aa4f90b9ca4658 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie8947b0e08f05ed4ed4888467fd64bbdacfd30fcadb77185a75e53a60bb78877);
            I8ef1e4ffe1fdc795a0b74f93f87b834e26e14a3a6cf78496df39c9cbdc70a819    = I7acd9d954e3db160301869bcb6aedd5652613816ae8340f271aa4f90b9ca4658;

            I0a66315056f6207395e960b11c230998d50db5a65f8414eda3a59ad04784a571 = I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 + ~I16863fd89fef9bef09bbfec8d23ba6d42f4de7902a5928e9b43546b4078fbb0c + 1;
            I1e3bcd83962abb7b063abe3da76e0bc387b63894a47a4f50f9ae7abce8b944f9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0a66315056f6207395e960b11c230998d50db5a65f8414eda3a59ad04784a571);
            I7bcdd7375cc16a2a91d81c5608f9953d21293d5121600dc475a15b190967b143    = I1e3bcd83962abb7b063abe3da76e0bc387b63894a47a4f50f9ae7abce8b944f9;

            I0f1690027b69262a948ece04cb1de6d4d7a358e60caa676760118364938210c9 = I9874305dca24f545c2727a64d4dececc7262d4ed5f72064a262cfc421cdc7c95 + ~I50f15058dc2e50a994089de4a0487158352c882d4639449d9db322a05ddcba3f + 1;
            I60f85c5d32cf353d7191d12cc29773a42aea456697214a1249353a6c2d7463c9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0f1690027b69262a948ece04cb1de6d4d7a358e60caa676760118364938210c9);
            I75bab5d1e71ba5ad182fb01cfa39d37572ab33f5f848dd0775e3358154e4644f    = I60f85c5d32cf353d7191d12cc29773a42aea456697214a1249353a6c2d7463c9;

            I97771793dd6517655733e9ced45e7daf0a11abb8377c42ad9710c40651558e6c = Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f + ~If4cdb00eb64cb9e80d78f3dedd797796f44f471b76f5ea3ddbc6f8521257e4c9 + 1;
            Ia9665e417120a907ca7c884c26250701f6c61f0e97c21fc62160f80c74ff05db = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I97771793dd6517655733e9ced45e7daf0a11abb8377c42ad9710c40651558e6c);
            I7f17ac4c0a37a850db6a1d3c1a5b2483c0f3afd684853df30d66933c8c593d03    = Ia9665e417120a907ca7c884c26250701f6c61f0e97c21fc62160f80c74ff05db;

            Ieac377a04bf039ea4d773d3e6e336e32f2cf37f375d79bf0867b5e7b7b269254 = Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f + ~I7af411084739689195bff036e9d5e9a950a7691f7d771d4d406aba4c32d95116 + 1;
            I5de5cb17db6bcb69528e636b4248c6995caf3e9f30dd363ac514f8f68d651ebb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ieac377a04bf039ea4d773d3e6e336e32f2cf37f375d79bf0867b5e7b7b269254);
            I6f8e6ce3128ce55b822fddcc664d0340c940bc85adbb5c93acff37548e3018fe    = I5de5cb17db6bcb69528e636b4248c6995caf3e9f30dd363ac514f8f68d651ebb;

            I887deded16218f24dd4ccc29a870e96b43b256ee62e0bfc6ff19c01fbe5b1ddf = Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f + ~I6eba99f7e39a1779ace2db8cd1806d099e7cf0678ec385baba570209f784b5eb + 1;
            I20647c051506a783956d48236b4a5097f9484e404c42e9176d52d59c8efe6c5f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I887deded16218f24dd4ccc29a870e96b43b256ee62e0bfc6ff19c01fbe5b1ddf);
            I3234faedbd9c50f29c09060c3f7ad76e44648841500b09c499875ea77aad9537    = I20647c051506a783956d48236b4a5097f9484e404c42e9176d52d59c8efe6c5f;

            I2b9966a73da68558c67e6cfe373b58865794a87b39dec4065056da2258197341 = Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f + ~I27737e1ab6f67dba3964412127cf6c91c7a58f6ba77e5b6a9808e2775069ad4f + 1;
            I898c9cd15d2ccc181e81531a379b969a0bcc87d38b0f3a9f9c413606bab42b15 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2b9966a73da68558c67e6cfe373b58865794a87b39dec4065056da2258197341);
            I74189716f0b6628c0d75d54cd0815cd8fa65b9047c3f51c5218fa0ba7b7fc47f    = I898c9cd15d2ccc181e81531a379b969a0bcc87d38b0f3a9f9c413606bab42b15;

            I6ac7d8576312302a7dba1bea496c3dd7b20faa3bbc8972a0e231f4e5ae3df8af = Ida5132aa4bd878e233d7875fb796fbcd9d0ddbc8cd652f60df8590d40010a85f + ~I0604d25b233f4206fb580d729452e9694d4b795553a4a788f993c992bc433b0b + 1;
            Ie75a482f66bf63ff96fb92dfaff210e0e43f91de86567ac2bd323fb0017a9f62 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6ac7d8576312302a7dba1bea496c3dd7b20faa3bbc8972a0e231f4e5ae3df8af);
            Icaffca7436caceaf13fa42e9e496c7b149d5931e08057ec92a73fbeb9e610648    = Ie75a482f66bf63ff96fb92dfaff210e0e43f91de86567ac2bd323fb0017a9f62;

            I5290a020c4e8d95084bdead6e37865decf5c9f5410048322c1f73361bbb49ef5 = I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 + ~I9e89eff507c5a2386876f56afb505a22f00d8c0f8a32635a00501ef8d56ecc6d + 1;
            I67d64752ba4f83a2592c0a83a7ff2773e71e84453dc882c23f8aec987abb6731 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5290a020c4e8d95084bdead6e37865decf5c9f5410048322c1f73361bbb49ef5);
            I13009f7de199aa969d82e233d26476e44aa1bfbb7d8a4fbfa0fe4f1f1e7579ff    = I67d64752ba4f83a2592c0a83a7ff2773e71e84453dc882c23f8aec987abb6731;

            Ia2fc1b624f958681d009ec01ed83d41c0e26c3c16ab0fe1e3ec4db7d0988255c = I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 + ~I63132df742cc353a39f27a7a5a00e0990e9e9e023f5c2a8bd571fcd6dd2d760a + 1;
            I37387450a3e4f68a3f1fb2cd428d54ffa4098528dce70e0a1fe3870830602efd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia2fc1b624f958681d009ec01ed83d41c0e26c3c16ab0fe1e3ec4db7d0988255c);
            I8c7ca4914849b513537d3688dc1b76461348ca06e80e489afb60a2a082e905bd    = I37387450a3e4f68a3f1fb2cd428d54ffa4098528dce70e0a1fe3870830602efd;

            I33974096440683b354b7725f26284e9c76a7d5722885b7ad9adf8630ccfacc79 = I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 + ~Ib9855ec95d5c99f93ad4c5565e622dc1c2d1c4a3b5d0937219172d97ac290756 + 1;
            I7db05f66d2fad420c57a7205c5a1b9d9036f088c64b58031e6fa82617923544e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I33974096440683b354b7725f26284e9c76a7d5722885b7ad9adf8630ccfacc79);
            I9117209a7cbd232356943389578d67bb7d6c217e7e40bdbb904fb46fb00e9385    = I7db05f66d2fad420c57a7205c5a1b9d9036f088c64b58031e6fa82617923544e;

            I8de6b3b4abe26905e4adae37762f35b8d1742281e0d0c5ba45a0531020a073f2 = I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 + ~I387ea75c114fd752ced502cc147dc9ad385dbf69607c04edf81ab74b6867f2bb + 1;
            I62c3f28235cae0fcbc04a55e0e578258ec501e25bcdef661063661346cba651b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8de6b3b4abe26905e4adae37762f35b8d1742281e0d0c5ba45a0531020a073f2);
            I0f16d6ab2d87cb715b071b05ad14fc6be271b1d7966b71c80795894643e6fc91    = I62c3f28235cae0fcbc04a55e0e578258ec501e25bcdef661063661346cba651b;

            If5011d2823a3b17fd74435029ee1469e792ab5a74fddd2d617c4d21b401781c0 = I2cddea26f7b1fa36b7e246e83f2dd4ae7cc47ec1a2a6425a8b05a46567587906 + ~I5b2860f88d7cbdbc92264ca1bd0f97c610e7b1cf340e2b65832553a1762fc865 + 1;
            Ib230966e790f9859c0c85bef2949dd2fb9fdaab81865b0b294036d12648fede0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If5011d2823a3b17fd74435029ee1469e792ab5a74fddd2d617c4d21b401781c0);
            I9fe8ab2f590451df0986a4f7a74194c27699bdfae0f182440f4c1875633cfcf3    = Ib230966e790f9859c0c85bef2949dd2fb9fdaab81865b0b294036d12648fede0;

            Ib4de4fcc7d35169a59e36a3af71a7832f967b7ae3c530c07cad1585784f7edcc = I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd + ~I206a4b82a444ed76c846a17eccf6c9ad62c42263b472949cc97f838f6a416073 + 1;
            I94c80b77b7ee413cd168e55905cfc4beb26ae2f6cbbb944ef335f47cf424086a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib4de4fcc7d35169a59e36a3af71a7832f967b7ae3c530c07cad1585784f7edcc);
            I57876d51522e735eff337a69dc597cdcbb100bb3d3e0e541aad4428637f34e26    = I94c80b77b7ee413cd168e55905cfc4beb26ae2f6cbbb944ef335f47cf424086a;

            Ica1376e18c562fa0863404b998af3c4e320f52008e7287b730de37fdb58e2dc0 = I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd + ~I37646f9ba79338e88c3d793a27911c88d573dc5c1cceaeaf565606c5b61495b6 + 1;
            I6ffff1f75581c6409c82505e1ad4216ff385151e7d592f1d59a1d983eedcbf82 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ica1376e18c562fa0863404b998af3c4e320f52008e7287b730de37fdb58e2dc0);
            I9fc6ec0055cf4788a1f382e41d1bd50b2ee07f2cdacf368e2075fdeef55f53b5    = I6ffff1f75581c6409c82505e1ad4216ff385151e7d592f1d59a1d983eedcbf82;

            Ia6251a913ec7fd4390c5330bbc9f4a983a37c274495a16d05dc96501050eac19 = I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd + ~I3e73f999bb1a0c087c2d4023920d56b1525bcb43f9d1bbc1b49b57d6c9c55127 + 1;
            I979f67eb071e28ab1fea67ea8e52910bd67827cf1dd23c07768c0c237703e23d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia6251a913ec7fd4390c5330bbc9f4a983a37c274495a16d05dc96501050eac19);
            Ib2ce92509ff0447a434264639ad96df47b161136cea1535b3e802c0c4ebc32e8    = I979f67eb071e28ab1fea67ea8e52910bd67827cf1dd23c07768c0c237703e23d;

            If46b3417b1f584a8866028e97e62402cf411792fdddb34faad96f0808ceb6d89 = I7d3811e635419361994befde0cc12bc4ba6c1b679f87a20ce15eea1e905e08cd + ~I62f27f0dc53be101d8fc7f026a673fd33a5397534153859f45c113e6820e9c26 + 1;
            I39e3942d2695061c6bffca3b7cbbbcd0c973e8412976c07d2387e9b05d75246e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If46b3417b1f584a8866028e97e62402cf411792fdddb34faad96f0808ceb6d89);
            I20b66d31e195a0db14cc87da1f6d8810b5f1056c2250bd5cfcb02fb4edc9dd0e    = I39e3942d2695061c6bffca3b7cbbbcd0c973e8412976c07d2387e9b05d75246e;

            I68dd3296bad4509893f3569f8b4e0539af4364b95ceefc0f95e3dffa5b90ac1d = I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54 + ~Ib5d22b614e704f01c688034adcd70603b8e69658cb66c96fe3ea76bdb323c222 + 1;
            If17d9a9ece84d9cfc9fcc430d453155458b6c8a7a3ecaad974c8f29d71b7d440 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I68dd3296bad4509893f3569f8b4e0539af4364b95ceefc0f95e3dffa5b90ac1d);
            Ie7595f637907686de85c9038415609949a80fee8bbb0c4e9f3873225ae6c56bc    = If17d9a9ece84d9cfc9fcc430d453155458b6c8a7a3ecaad974c8f29d71b7d440;

            I7e32c30199d506efaf13a091029320249c5a524f32b0e55deacea536599a92e9 = I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54 + ~I0b2f8e7646b38057090faea20bf55e51f17d23baa4daf0c16d00e75e4c5f0ebb + 1;
            Ia3496c8ef63a7e37f4836fd3f0bec02370cc7614a22a1756e61fa1a536f942fc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7e32c30199d506efaf13a091029320249c5a524f32b0e55deacea536599a92e9);
            I6d41031fb10896690dda6067df08ad914896baaa5f83c46b4051cd5a02f3baef    = Ia3496c8ef63a7e37f4836fd3f0bec02370cc7614a22a1756e61fa1a536f942fc;

            I97f44fd7abe7a43044027a60cc8b9e88d1c474e613b30fb092267b7d8e0d0748 = I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54 + ~Ie3cada5731ce9e6c51353952cfb87527bca19aa77436766bdcc843dd92f1cc60 + 1;
            I79473cb7e5feaef4d80685528a576e134e739af85c92bfc85278f949ae938a96 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I97f44fd7abe7a43044027a60cc8b9e88d1c474e613b30fb092267b7d8e0d0748);
            Idc6c8bd2a37e01dec18007c8fa763941f7016bf299e3cebbbbee3066d4bf8c7b    = I79473cb7e5feaef4d80685528a576e134e739af85c92bfc85278f949ae938a96;

            Ic9b7ae6f6993eeda2a7297af8e3a9301da5055c1031f82fd99451e607ef70738 = I8266457bff8d64b26beb6ff4bb81dce20c26e07e8c6b3c27057818116cc53e54 + ~I92cfa50424ddf1ada795366ac6c7b31cbb1b1330486911824b881a1fda443c25 + 1;
            Ib6f1e860bf50cfc54de5c515cb40c392f0fd1f02c325d52c5e28cb5d3a811a48 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic9b7ae6f6993eeda2a7297af8e3a9301da5055c1031f82fd99451e607ef70738);
            Iac1565ee006c23dca041f0aaff4dd7023b8a22cb72c9f206170be661a66d4732    = Ib6f1e860bf50cfc54de5c515cb40c392f0fd1f02c325d52c5e28cb5d3a811a48;

            Idd55fba0f9374647ac6e708497c4118c4493602ebe8f342e6ffa87b496fb92d8 = Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979 + ~I876c143c75e838720b2a1ee393f5da5ba08822ea13fa1ff459d68d7b0c0e5cd6 + 1;
            If9f2c8dcaceff8232ed4bdc9261d1ee5adc0291873452c335748d5bcca9435a5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idd55fba0f9374647ac6e708497c4118c4493602ebe8f342e6ffa87b496fb92d8);
            I7318d295676d4cc0682f246020963a6411be5cfc2fa525dd7af0f2e651b4f9f8    = If9f2c8dcaceff8232ed4bdc9261d1ee5adc0291873452c335748d5bcca9435a5;

            I94a0208aa6cc55e3ff0c47d436cdbcccce15887177af919270ddfe9096a0a7fa = Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979 + ~I43bd10e4f520ec08b30e8474404cf62a6ad869cdd1d280a2d221e0d76f228091 + 1;
            Ic215b986ae9a8ff5c760e17d5e71da08756ba48d0f8874e35766d0f8fc18b061 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I94a0208aa6cc55e3ff0c47d436cdbcccce15887177af919270ddfe9096a0a7fa);
            I596ee6206f54965079551ffb23aa3c1948f6fbcd48659c4e30b205dd06de79f6    = Ic215b986ae9a8ff5c760e17d5e71da08756ba48d0f8874e35766d0f8fc18b061;

            Iff2621e7d8b4bb5de9b649f5424e482b9dd4f01bb7c5609ce8eb76766e301d6f = Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979 + ~I00c96393d166280a0d866d1999d4306a650507c7bc407202924f6684f61e219e + 1;
            Ic945b809e46ac7f930479330040e1b167e8f5b96a0583a39713a34261e764ffe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iff2621e7d8b4bb5de9b649f5424e482b9dd4f01bb7c5609ce8eb76766e301d6f);
            I7c8c24bd3806dbea5552d386a7363828eb5a822bb292fa0c14ba407a1937d11d    = Ic945b809e46ac7f930479330040e1b167e8f5b96a0583a39713a34261e764ffe;

            I8f5b316fa91d4e39b9eb94d7d051c81e4e95dfa2a2761af7970ff04e6ad1056e = Id92108625a8f677dabc536455746caca3a9d0dd548358689d40358b7d3b3b979 + ~I1d996fec699e93fc4ce63060990c6347d998a81f0b3aefd88339d5d620fd152d + 1;
            If6a91bef840a62f8234c19c7783b8ec5d1910ffcc05eae66cf63c1bd541c5caf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8f5b316fa91d4e39b9eb94d7d051c81e4e95dfa2a2761af7970ff04e6ad1056e);
            Ib7690a963a38d899184e89d3e51ac5cd99cc0ea9b2fca1c2e36e51ea65b893ac    = If6a91bef840a62f8234c19c7783b8ec5d1910ffcc05eae66cf63c1bd541c5caf;

            I1cbe0e864523810adb559c85aeda0f79a1dd57f819e9904d4635023fa1a689a6 = I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1 + ~I3dacdb67f2492ed12375b671dc593349c75562e936401def91b4391c153fa572 + 1;
            Ibd9c2cc79d2377baf6c47290fb8b0671bebedb2aa72b90f8d9fe98d0acfad39e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1cbe0e864523810adb559c85aeda0f79a1dd57f819e9904d4635023fa1a689a6);
            Ie55d9e9e5c4a66363393994597d9138fccd6c11a2a6c939768b63d9cf933ae1a    = Ibd9c2cc79d2377baf6c47290fb8b0671bebedb2aa72b90f8d9fe98d0acfad39e;

            I03c8aad8e9fa3cbae4ea5779a2db031113b6bf72ab3df44995217640c7f52cb2 = I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1 + ~Ibdfea3d72843376261dc3e06e3f19be4556508098d1b4d37c1c4cf6928860719 + 1;
            Ic655dcfe5a7d40fcf2eb0e61961010434f0098e4cb08794fa7963797c764bac2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I03c8aad8e9fa3cbae4ea5779a2db031113b6bf72ab3df44995217640c7f52cb2);
            Id2a5a1513f2b8c1f000f58640c3650ae03d4d56205a8cbd04742be5b91c8c594    = Ic655dcfe5a7d40fcf2eb0e61961010434f0098e4cb08794fa7963797c764bac2;

            I9f9f7fe2510dda62df0c857cb4ae9430a8c435a64bf84a6d94848e53bea684f0 = I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1 + ~I67a45b7ce414632252362c1556be0e627757c871c136d8570d4300fa316205d3 + 1;
            I302186a080a24d93f21320fc1165055fc1a2cdfb86171f35cc5fa8ee98f0e1b2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9f9f7fe2510dda62df0c857cb4ae9430a8c435a64bf84a6d94848e53bea684f0);
            I9a2e9ef69e2c24fdb342d3334d2b71a1bebf10ffe1518dc5f3ebd5ff34dc719a    = I302186a080a24d93f21320fc1165055fc1a2cdfb86171f35cc5fa8ee98f0e1b2;

            Ie596b7fb4376d234eeb9946c5e2d5439cb738fe881235324c8d333cf0283adf2 = I7124f9fd7e7adaaceb485ba5327eeaad1973342ab7415ba4e3c0a6dcdd6803a1 + ~I33546fedf41dca9168afd7d6916823e8c24aa3c4a855b93820215c68c807a56e + 1;
            Ia3900ae4b178203e8a6aab20f112207ecbe30e66c7fbdff63d82e1bc1c9ef760 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie596b7fb4376d234eeb9946c5e2d5439cb738fe881235324c8d333cf0283adf2);
            I8052be48c5148738c00fa7e5be66ac6898d51e7fca2e5905ef028d897d47b236    = Ia3900ae4b178203e8a6aab20f112207ecbe30e66c7fbdff63d82e1bc1c9ef760;

            I44d6eda047420415765497d6523a69b8ba7903ba7a76658dbd8f84d079bdc416 = I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be + ~Id8832e8e711bb3e7fe9136084b9832a2677803cabec7f2469144eb3b6d4ee3ae + 1;
            I4734d2e489a9d1d0d797602f00bbd0e63d76f1ab0bbc514401ab815d5ebeabaa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I44d6eda047420415765497d6523a69b8ba7903ba7a76658dbd8f84d079bdc416);
            Ifc4766e0c1913ae910a794a3de1155638a9352251d646b270e3aba4eac09aa31    = I4734d2e489a9d1d0d797602f00bbd0e63d76f1ab0bbc514401ab815d5ebeabaa;

            I8677eb1f6f7ce797b6e713913227fa9a6d2953074c6b4208dcd3a04a1769b3be = I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be + ~Ibba131ee71ced96650ce76aa4695641a089046f8b8345ba312d6868dfbfb2787 + 1;
            I9d325e738820d37fcdc02fddf7899f4e910dc410218c77432a6e47f1f9a956f1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8677eb1f6f7ce797b6e713913227fa9a6d2953074c6b4208dcd3a04a1769b3be);
            I2322db4da4e5112d362e202ee964c08830d852a01c92f802c1c8bc2978ba25e6    = I9d325e738820d37fcdc02fddf7899f4e910dc410218c77432a6e47f1f9a956f1;

            I1df660831634377e177514ff041dca7c173c608c37c0dec5233ed65899fae519 = I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be + ~I16778a093510ae433495baf9d2b7a74ad4c5315403d0e8aa39eb09cf508dc201 + 1;
            I66cfe3b553e345d01602cf9440774c8383b14922fb66580046e0819ce297b0f5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1df660831634377e177514ff041dca7c173c608c37c0dec5233ed65899fae519);
            If29e3e5b3c3425bf0fd40a98d32046f215032a8ae181688dff1c4a253b0460ef    = I66cfe3b553e345d01602cf9440774c8383b14922fb66580046e0819ce297b0f5;

            Ia5900c9e78693f74b25f0c17c8dd79a78f7187cd79892df701f93314cc71963b = I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be + ~I72e85032ae85773b79f3a3dab895c9667cd32c6aeb44c000096ddcbc0f7be0d5 + 1;
            I00c3f248f180ba740d0d97e10760d76e4d9033a2e4125b04ff783a554db09b1e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia5900c9e78693f74b25f0c17c8dd79a78f7187cd79892df701f93314cc71963b);
            I51e9d69995015664cbb95900d25d26d386de1f49fa7b7d612964802060fd7a8b    = I00c3f248f180ba740d0d97e10760d76e4d9033a2e4125b04ff783a554db09b1e;

            Ie8edff06c26702bf20142c7cb6eb605bfd52076483bbd6e941fddcf87518f184 = I0a453b18c9ddf27bb60fa77117c2b44941545a973e2def031a6fab533dc073be + ~I8617f958a4de5cf233240840c770360befaafe599fbec1e351b24baf301ecdbb + 1;
            I9954c6247025cfb8b0264906e6dc6a703b9dc8d3c4f2736930fe68d278dad962 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie8edff06c26702bf20142c7cb6eb605bfd52076483bbd6e941fddcf87518f184);
            I2af69278f44ee2d81c64b9447b85bd09d2ce2a8dc86bacb9a175b33f72d4f851    = I9954c6247025cfb8b0264906e6dc6a703b9dc8d3c4f2736930fe68d278dad962;

            Id858a113ed0d9d3e0b3b3041add0654aa217c3781cdcfc32a081422edf6c94a6 = I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac + ~Ifb337611e63cb9cee9828aa75fcb6d978249e65bcc8770d51fb4dd1644c96a86 + 1;
            Ifc519e00af8bd07f427774d04fc48f95781295dfe970673d84feca42e324b583 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id858a113ed0d9d3e0b3b3041add0654aa217c3781cdcfc32a081422edf6c94a6);
            Ib82fbfc182e6598a7a8dbae45ea083d2922e3f10e781ac40e1c89f79097f1f23    = Ifc519e00af8bd07f427774d04fc48f95781295dfe970673d84feca42e324b583;

            I63688514e288f5d828f22310d609beb495c809315db245d6cb783e02d21aa354 = I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac + ~I428333658d20f4417e24a58fe364d5a647332ef76ecb7f15d83dcccf1aeb3d11 + 1;
            Ida260241e2192ba6e2a1d15acbfabfce6023278ca1f2be17943bf48d0b95d045 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I63688514e288f5d828f22310d609beb495c809315db245d6cb783e02d21aa354);
            Ie3180a2d7f37d66f9895c1de89329e69ef7e88d0808fce147b25636e639efdd5    = Ida260241e2192ba6e2a1d15acbfabfce6023278ca1f2be17943bf48d0b95d045;

            I402c6bd3528da160ede7f8c92d97a0c27835b1fd267e14fb8d92706f13719570 = I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac + ~Icdad18f8878b4e9645b4f2d2434f913a6e0f732a20a6a750e25c2398a086ac2d + 1;
            Ief91e723aebbfa64c457be6ccd3ed8e2faa4703c627ae36bf868d8d970bc315a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I402c6bd3528da160ede7f8c92d97a0c27835b1fd267e14fb8d92706f13719570);
            Ifb545544cfc26097f08bb8236d489536608fd3ef900015de2da0a8a5dfcd44ef    = Ief91e723aebbfa64c457be6ccd3ed8e2faa4703c627ae36bf868d8d970bc315a;

            Icfdc65f513f27d474c48d7fe42ed9134e668a9b706d011dad7025214c61c5c6a = I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac + ~I8d10cf5dcbbd1a765ece13156db0ad4651b41cc5ee286720226649a707accd16 + 1;
            I53a559b412f643abf84ed01e98377ed96246560bb003bd28eedf2164de2c2db4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icfdc65f513f27d474c48d7fe42ed9134e668a9b706d011dad7025214c61c5c6a);
            I90ba4bf676fa4d1eb6132a37c0b4a580ef39ac1cc44d6111b84d6c7b907922b2    = I53a559b412f643abf84ed01e98377ed96246560bb003bd28eedf2164de2c2db4;

            I59cbaf9b106eecde3385e8d646545284791f53e64fef5d89e72699fdf9d66786 = I1f0d6416c6b6a2754159138b42abe65479387083e0c9d319abbd6dd6836466ac + ~Id824ed4e68ef3624b9a4d6c5924b08a7b727df62fc9135c973c5f79768c627fb + 1;
            Ie685d62aec7093c42c2c432f32fb1bca42a9af0ceff50f2ff2ffe57f0d98af75 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I59cbaf9b106eecde3385e8d646545284791f53e64fef5d89e72699fdf9d66786);
            Ie66d53b4bed43cf8037cd1937f7562e7bdd6cac54cfc8313572b853088528a0f    = Ie685d62aec7093c42c2c432f32fb1bca42a9af0ceff50f2ff2ffe57f0d98af75;

            I80b1e51f33d8c209746c92f8e1d059c87bff5b4f169bf9304bdd30f96c5b1d8d = I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 + ~Iac435cdd22e5425837ad24bd6141cb357c302af7ee7637e1cc2ac25474cf7506 + 1;
            Iaa2f1dc17d04b53a43d7435ff62012f950453b06af95243f1e1fae92885e9480 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I80b1e51f33d8c209746c92f8e1d059c87bff5b4f169bf9304bdd30f96c5b1d8d);
            Id812808edf2372138b1569ea1a2ae0583ef70eaad98a941b8394d5d9efeb44c5    = Iaa2f1dc17d04b53a43d7435ff62012f950453b06af95243f1e1fae92885e9480;

            Ic36894855099edb8618f29e72154ee32f3f130987bdcd435cde2f87ba39aaf0a = I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 + ~I886fbef883afc3146952de2fc934131aeb38bc2134c096497981d303594f1f37 + 1;
            Ie74bccfd27d7ef80fd7b51b8e57ade889188901b44e7236766861e8e9601fed5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic36894855099edb8618f29e72154ee32f3f130987bdcd435cde2f87ba39aaf0a);
            I6b9daca681053a70322aec979459e65099a78668854de86dd3f51ad58c5dced5    = Ie74bccfd27d7ef80fd7b51b8e57ade889188901b44e7236766861e8e9601fed5;

            I676598186f1a742ac68bd8a533c205b9b5cc6aa540b0519a995388d5db421574 = I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 + ~I3b3f53fca961a376010d1a5b0c49f91d58b351d0306b8433ac22a70f5a1f1673 + 1;
            I4d27f6db1cba68a36e75da65709b30702412affd297564d2b4e563e41db875f5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I676598186f1a742ac68bd8a533c205b9b5cc6aa540b0519a995388d5db421574);
            Ieafce3772abd32b8004981fe3f3d102d629075a15b6dfff65169984219911dd9    = I4d27f6db1cba68a36e75da65709b30702412affd297564d2b4e563e41db875f5;

            I2212dc39f8bda130c6782e104418cbfea3d2089b3d0fc700e8acbebf1fd9d296 = I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 + ~I58d3b6391c1720bf6ac7458ce499fe3b0573e8f7f324db1a796d1126e42e57a6 + 1;
            I0fd6ce3dc520f3fb4fc9a66c0abe0c05b943610bb0bd11b7f9dd10befd5c0b99 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2212dc39f8bda130c6782e104418cbfea3d2089b3d0fc700e8acbebf1fd9d296);
            I279bb276ee61f29e0c143251191c161862c9d95cf0bf3a3fdcb6b3d6acaee983    = I0fd6ce3dc520f3fb4fc9a66c0abe0c05b943610bb0bd11b7f9dd10befd5c0b99;

            I371e726b1f426a879388bc0d28dba55143a4674655374dd183793fa42b8bb67b = I026613966a447de48dcf9ed49a02404926befc89b67557a293b66303e737da28 + ~I3d71ea5bb4c4be8ea80abe59367519a071132c913eaa5c6538baa8c3faf243d4 + 1;
            Ic7a11ca0ad51e87c9eae3a026eaaf462f9f4757831277dccbd25881de07202e0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I371e726b1f426a879388bc0d28dba55143a4674655374dd183793fa42b8bb67b);
            Ife98dd3babdd2b2db4edbc673874d3f8f184f531c9d96b1a89b68ba60a9a57d1    = Ic7a11ca0ad51e87c9eae3a026eaaf462f9f4757831277dccbd25881de07202e0;

            Ie412b52497a49cb060e42e15db8793b4af98294d202c14543413a6e30de8fe09 = I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d + ~I0d6546f557347e1d72c176a40dcb077c9c4c78ed89975154f5bbb3875eb1131d + 1;
            I9abd971b53c2f6c0d24fd41004554d3175db4b8fd63b38c7667ff78272cb26ee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie412b52497a49cb060e42e15db8793b4af98294d202c14543413a6e30de8fe09);
            I038f11e434287c1e184cece6178f4ce26889bc2ea583aba8889b8953306e2e60    = I9abd971b53c2f6c0d24fd41004554d3175db4b8fd63b38c7667ff78272cb26ee;

            Ie3226e6cc2a926d44860fbdba32984e2c3a007c1dbc172c3765cecc6bf4efba6 = I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d + ~I88e5fe043e16a274d915245b02d2094d05fb7710f6078dd6b33c2a21676200c1 + 1;
            I24d9c2b238ea5964b3c4bb358f301815fa15836cade3b5ab5ceb0e81a6d3a6bb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie3226e6cc2a926d44860fbdba32984e2c3a007c1dbc172c3765cecc6bf4efba6);
            I25c61073e64c8149ae96f3157045d317349321841e21a3d69b3baf3bd70bbd03    = I24d9c2b238ea5964b3c4bb358f301815fa15836cade3b5ab5ceb0e81a6d3a6bb;

            I7be3e45435a982ec33d6b56aef2c5a81f233859f8312e4b328c0a9e8c11b5822 = I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d + ~Ia2343365eee39c9305def2bd744d3e44bf20b5bab8a48c6a2d95908f74f3cd18 + 1;
            Ia755a5da1132f62cc35903f93050e9743df11befaba728cfa055601606c0caa5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7be3e45435a982ec33d6b56aef2c5a81f233859f8312e4b328c0a9e8c11b5822);
            Id156956a3b93d6a741a81c5a94e057e054ad7d4467a54a691bbd147afb30ead7    = Ia755a5da1132f62cc35903f93050e9743df11befaba728cfa055601606c0caa5;

            I5363dc622b9c481283f71015f9fb2a340bf5f440344dcabd8adb4961a89bb36e = I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d + ~I1d5510ca99815d74f26804206bac7f1e7eec3727fa89d91b014becb49a815abc + 1;
            I4646084cb89b559ecb864051cae61dc568e6b9c6db4f1030904a572f7e58a22a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5363dc622b9c481283f71015f9fb2a340bf5f440344dcabd8adb4961a89bb36e);
            Ie4eea240addf4997dde0e268e6404bea936a04629cd4d244a101a6a38e6ec03e    = I4646084cb89b559ecb864051cae61dc568e6b9c6db4f1030904a572f7e58a22a;

            I194ca19f61c5d4e4df1e7cb9398ea02166bb2f231546f23d151370c7bd533425 = I808016dc266503fb14bac0c9ac1e7c8d4d9f1fe3da2a45d6d8c38099baee951d + ~I6adbf5489cbaa65213fe0804e7494a2b8be9db9132a6ab7058764a1a53480999 + 1;
            I58754d218860b8400d1e6ffc21c817a447bb64d182e74f0d162abd70e15c5db6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I194ca19f61c5d4e4df1e7cb9398ea02166bb2f231546f23d151370c7bd533425);
            I536f7bfebdfdbdfef2f9b530022a63e1a70a1ef0b344d7f34ef956bed72fc94b    = I58754d218860b8400d1e6ffc21c817a447bb64d182e74f0d162abd70e15c5db6;

            Iabf25360f3e96668f6ed500de6bde88342e176aa39205579d171adff86c5acf5 = I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 + ~Ifc4886636576352e5307fb1fefefded0d693fd059a3fcdd6b4c9dbab1b908114 + 1;
            Id3a8f1a1dfbdbc1705527f0e6f864ae594bdb100ee8b14a349147d98da860f09 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iabf25360f3e96668f6ed500de6bde88342e176aa39205579d171adff86c5acf5);
            I53a83ec9af418aeb6869bf9db2b0ce128564fcf62d2a16506906303025076ca3    = Id3a8f1a1dfbdbc1705527f0e6f864ae594bdb100ee8b14a349147d98da860f09;

            I67a8f91668c29b02c6638bc4cfb4d99364679a1e19ae54b6928adccda64333c0 = I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 + ~I2fbaaffcceb2dc6a4f6d9d34140997b18356dc3803bb0a6c6d5f1b3f980e18da + 1;
            If36c8f00155dc15627d5005ff98abb7a6eebcfa62de82fdfa50d86fc6e7cc166 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I67a8f91668c29b02c6638bc4cfb4d99364679a1e19ae54b6928adccda64333c0);
            I4644d5f1dfb72ca4669b26a415cb9aeb54051fe8d28a6461d696f00bdf6c930a    = If36c8f00155dc15627d5005ff98abb7a6eebcfa62de82fdfa50d86fc6e7cc166;

            Idd22bb99613e9b5b2120390d00fc41e25227523bc60e6d281f9ab3e0d9eae0a4 = I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 + ~Ic56053af1a36bedb5e1670282ac0a93d782faf76d25a25edab3dadb09a302de1 + 1;
            Id97692b9a9b0e7edbdf517b47ed0b87d007cca8fafa703956ffc2686b727ca9f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idd22bb99613e9b5b2120390d00fc41e25227523bc60e6d281f9ab3e0d9eae0a4);
            Ie02a7d9471f0915572b8db6797d0ea1f2fa380d96a4e02a5783e584800e6676b    = Id97692b9a9b0e7edbdf517b47ed0b87d007cca8fafa703956ffc2686b727ca9f;

            I3234917db6bb05ba543d97c095bcbf419df98d4fc7a64899f340864d7965708c = I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 + ~Ia3690db3bb1809f3df1fcc3a2dd5f807a0ef26c4cf61810b0f9bb590951f8e36 + 1;
            I3391de01ebddc6f92c31c74e3b3ce12ae2081b56b461ce9e890a0fef3d14fadc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3234917db6bb05ba543d97c095bcbf419df98d4fc7a64899f340864d7965708c);
            I0f39af323e102d03f5089838b2b6576c03169135defb533f54e57d8450f1130e    = I3391de01ebddc6f92c31c74e3b3ce12ae2081b56b461ce9e890a0fef3d14fadc;

            I111227fa4bd1705699775e2dab468800630a0faca805bac5a9bc6d39e3e0c721 = I3ea2934ff44f79e8b1f96680610cb65dc6993d926a5d30be6b4b699408a3f1b6 + ~Ib4e392b7b8f87358dd5cdefe7c272531bc6bb1f27bf1411c1a2f4331809a83c5 + 1;
            Ia5f3145a0720b745a384e157d352823fe10bb6436875a5c52ad6c81c882d9e9e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I111227fa4bd1705699775e2dab468800630a0faca805bac5a9bc6d39e3e0c721);
            Iaaee3c7078bf1bcda85bade0d66984c675177a0f1c66c58f47e3775916797a57    = Ia5f3145a0720b745a384e157d352823fe10bb6436875a5c52ad6c81c882d9e9e;

            I17f10c5cfeb0d1c9030ca3b64a6cccc65dc578fda6a627ac3d0d0c03aea66041 = If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee + ~Ib897fb3696e7d68b81ff3c1573f5cc234d32e10d066864ec203487a8e56f4ece + 1;
            I8f807b6151726e387854a9a6c778b3b069ed5ab61b41aef6541f3c2330b71673 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I17f10c5cfeb0d1c9030ca3b64a6cccc65dc578fda6a627ac3d0d0c03aea66041);
            Ifcc101725d905f243fff4a458ab8da67311d5563911d69daad960072e1927054    = I8f807b6151726e387854a9a6c778b3b069ed5ab61b41aef6541f3c2330b71673;

            I2d431ffdead0e5f6add0bec3d162c7045953e597d33fde53a111f929f278b8d6 = If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee + ~I15ba9fcccc2e3aaba7bb5967d35eeecfc3bfa7ce27f82435be6dee9d0a4af829 + 1;
            I6bb8ab1ec9d2824241e526c7aad88002dd83769fe53a79caed88f4f25929dc8e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2d431ffdead0e5f6add0bec3d162c7045953e597d33fde53a111f929f278b8d6);
            If5e789a890f931a53acd095741f7a5936f15da9e0007b159a3a3762ec13223f8    = I6bb8ab1ec9d2824241e526c7aad88002dd83769fe53a79caed88f4f25929dc8e;

            I57b332bb53fbdc45a8274e8a6838c2d3722677a6b560c2379ab92e225f4aa64a = If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee + ~I2cd11587dc2659cd92fb2c4f894bbd9d252affb93f75c3c691dbb02225b4e887 + 1;
            I5637f02c1a3f8b9ac950dd6a246e2721f9e4d30906ec3662975bb3528e3d7170 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I57b332bb53fbdc45a8274e8a6838c2d3722677a6b560c2379ab92e225f4aa64a);
            Ic7fa79c98c1eda80a19d8475857fb44ab41c53596b0b59806fa776d4c4ad02f4    = I5637f02c1a3f8b9ac950dd6a246e2721f9e4d30906ec3662975bb3528e3d7170;

            I3ae1dc3a3f40ad8a03dac4c2c2b657d83c3522992ba57052e238fbc8b836af26 = If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee + ~I241e6ca6efe96759bbb20d710c448c9c322aa3345fcdbedf625e297070af52e4 + 1;
            I2f381294ee877c6e693fc57e804a48a9efe7e3289f2967a006a7da1659cfaa3b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3ae1dc3a3f40ad8a03dac4c2c2b657d83c3522992ba57052e238fbc8b836af26);
            I6c1edf3d3971f7ab6f93e50a9500cd37fa3bb42d75c70d236f514e4c15a61f2b    = I2f381294ee877c6e693fc57e804a48a9efe7e3289f2967a006a7da1659cfaa3b;

            I0980470783afadbf12692805326a5b81079ba76f1c19e80bc7f0a30e73a5294b = If6b4c8f9f23ce5c85ede8598d77210c4cc284664dc46386f75a5e7fe3ad3bfee + ~I6b528ad76bac25170636a86ebaf7efd14ee7159ea2c83500021e39e968786428 + 1;
            Ib31ed62a3528251d6f00b4c346c776a8d5c3906b66e951288449677cc9865773 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0980470783afadbf12692805326a5b81079ba76f1c19e80bc7f0a30e73a5294b);
            Ic3234b24482f57a12d4db307382a5591bd66ceb0dd4bb120eadc7ab2770d003d    = Ib31ed62a3528251d6f00b4c346c776a8d5c3906b66e951288449677cc9865773;

            If55dc3c3f903107602154e84ff4739788ba44ad35a05bdd8e2987d02dbfb165a = Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 + ~I101eb18f34badddefbdefe0c2448e2a8a243e4803ef3244b25365881bf227145 + 1;
            If6073191b5a616ca29300286d02c0ea3f8eb57da345d41625650caac734bae9b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If55dc3c3f903107602154e84ff4739788ba44ad35a05bdd8e2987d02dbfb165a);
            Icaa9abc6adde275d5c5011fc8cf6ead11032cc1bfc286b3a392ec507e4ff0d4c    = If6073191b5a616ca29300286d02c0ea3f8eb57da345d41625650caac734bae9b;

            I6aee7f7827cffd92b9148e455718c252b04105a64b8d9c60ccab52ee1ec08e31 = Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 + ~I20ac47b3e52f25ce7858fb7952654107faed4cb5cf3abe1ba915710d1af4c933 + 1;
            I2ac115af593010e9556a2ce7fe8e479b1d1d15b34750a8084c442b1be7a181df = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6aee7f7827cffd92b9148e455718c252b04105a64b8d9c60ccab52ee1ec08e31);
            Ifc444a5134bbeeda6005a847d5ce4e180e6c809776e32d1ac709c3827d1d84b4    = I2ac115af593010e9556a2ce7fe8e479b1d1d15b34750a8084c442b1be7a181df;

            I619b017a1e80738f224764b9062ff6a3b9f2321eeb8fec5ec95573033d33a9af = Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 + ~I51abe903b403df434eba534a1102cabe0a0e976c047fc5cc97a6c8e73263c531 + 1;
            I306ef55d92e069bbb7dcaaa61fd648d31d246928bed83dd8b2764f94de45356d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I619b017a1e80738f224764b9062ff6a3b9f2321eeb8fec5ec95573033d33a9af);
            I41fff62fe024b1bc1071aae30dd931c1dabf2e12d0d1cdc295bbbbd946d63358    = I306ef55d92e069bbb7dcaaa61fd648d31d246928bed83dd8b2764f94de45356d;

            I812fbc992824cb1e29cc2c40421e63ca06fb97c9d9e40094473cacafea5f0e0c = Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 + ~Ic7abe3b0fe121e025ad7f7802b7800f4097111a1108ad088e869e81e5374c42c + 1;
            I915bb804d2926482383b55712d495d9d5a5df9ef4621a5ff8a2a4d5bfc882c09 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I812fbc992824cb1e29cc2c40421e63ca06fb97c9d9e40094473cacafea5f0e0c);
            I8ef6ca3a27d76c9635bc942fcfb21cae619dc5b7bc842952e2a29f7f2915e62b    = I915bb804d2926482383b55712d495d9d5a5df9ef4621a5ff8a2a4d5bfc882c09;

            I925edaebfbe72a77427ff9387ca2b955f2eaf2c3b6d76bc14f6acb37b4f98720 = Iecbf6b74e90a26b4aee9899a15ef638effd639adddac3e31b65c214ca0f644d4 + ~I294be7c0765f0d4209d4442136d706edb2080883d5c78a3c71d66b5946116bef + 1;
            I6cdb31ece4d35306b0d4aea87dff3b178f6664744c85f6307e1c1d6153d74c72 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I925edaebfbe72a77427ff9387ca2b955f2eaf2c3b6d76bc14f6acb37b4f98720);
            I1ec8e7e460c616e3d6459dd35f82ebcebdc1bd7f9680c38489e292be831ada10    = I6cdb31ece4d35306b0d4aea87dff3b178f6664744c85f6307e1c1d6153d74c72;

            I5842c1f6bd94143ce3217369de2df9d5f2035e55dbc619313375adc7bd97f727 = I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 + ~I82a2a0149ccdf627e13b7d422945e626fa268c22b3c30bbaadd0a8de14ddcf32 + 1;
            I4282e3203fc14bbe70311010f6132cef075c94dc8fe22dd1f115e58e560c2652 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5842c1f6bd94143ce3217369de2df9d5f2035e55dbc619313375adc7bd97f727);
            I3c396eafe78ef3a7c94cae71c86a808a9fc88960e7519256fb1c0b54bc865334    = I4282e3203fc14bbe70311010f6132cef075c94dc8fe22dd1f115e58e560c2652;

            I2af5890840cbc6f131cf8cca27929dc20330f4248a5d7b5071de85d941bdf2e2 = I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 + ~I0738f605ff9ccae9ae63f8e6fe7a9b537d97e13bf3f23c7b0daa4fc414eb7eb4 + 1;
            I98cf027b8e2ef347c03bcff057b551436e1b053e2439164297c60094d957f760 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2af5890840cbc6f131cf8cca27929dc20330f4248a5d7b5071de85d941bdf2e2);
            I78382168abd43ba48f24ad5e574782b47afeeffe0632ae5b4aeff07ebedabf4f    = I98cf027b8e2ef347c03bcff057b551436e1b053e2439164297c60094d957f760;

            I01542998e0af4239394cf341547e6dc36ea36f77aa1f2b371a6f915e99846f20 = I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 + ~Ibfb1cfcf89fe21ebca17ed6bd834fb8567cef4ccfb8f03fd5edaf59000ba0cae + 1;
            I8a156bf85802162d32801b45b639076f8ba98827cf96d3e1cb48a5a3b774b491 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I01542998e0af4239394cf341547e6dc36ea36f77aa1f2b371a6f915e99846f20);
            I55de212bade4801bfd54acbc885f19f7f43fc63874f6a531f8289cccb06c81a2    = I8a156bf85802162d32801b45b639076f8ba98827cf96d3e1cb48a5a3b774b491;

            I1ac783cfcbbcb2dd26bb3b2a766481a364b520ff970a1ae49f52048c0cbc228b = I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 + ~I55d5daa0c4cb89aac08ecbaaaec1d6afa2379b277051281d3c15abaa6af05edc + 1;
            Ia9058e9aec6d06a5fa6d715e681719f75ca9938f6fecbce752a4d166fb9f2bca = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1ac783cfcbbcb2dd26bb3b2a766481a364b520ff970a1ae49f52048c0cbc228b);
            Ia4c73e87649527da20616919420137fa4c1c8cfb4c85f4728a8441109168c6ad    = Ia9058e9aec6d06a5fa6d715e681719f75ca9938f6fecbce752a4d166fb9f2bca;

            I5ab65b455c544d54467f0a12db6ff74521cebe6cf47f583a02508f73674f5bca = I24c3922a2a3068b56be2370753404ae70f2a5f66b72bddbd7bff1086eb196116 + ~Id834a34ad825df7c595e3754b5a5638badf560cfb68ec8de2903e73e88b1a113 + 1;
            I2db4e765057361b39c8d20e87f89051b0016f067baa15cf01865623088a9b984 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5ab65b455c544d54467f0a12db6ff74521cebe6cf47f583a02508f73674f5bca);
            I04eb84d9339dab27e5615403aad9f09e40f6b123c73c8c8fd6c27f8e91ed4af6    = I2db4e765057361b39c8d20e87f89051b0016f067baa15cf01865623088a9b984;

            Id3731847bbab8d64f89de08c1fd5a8a089de6eafc93e0a079bb7e0a990d3a010 = I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347 + ~Icefdcbf9ca1f8e02b93f295ed8dbc43258b29cbc0cdf9c9ed5fa60117263d502 + 1;
            I4203cf0a99cde14acce3ce3c04a6405aef0edfda7026924b1491de1d42089051 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id3731847bbab8d64f89de08c1fd5a8a089de6eafc93e0a079bb7e0a990d3a010);
            I49fac311626d99832accfdbaf5db0e3da11e0d89693c843295ada1310a5d8f84    = I4203cf0a99cde14acce3ce3c04a6405aef0edfda7026924b1491de1d42089051;

            I519df6e33d8ef22d52e32b8119be2aaec1f50dbccc5d79dbae0f55ceb6cb8f18 = I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347 + ~I3f3cf1014fe01e02bb46b2e8a19716cfaecfec0e44fcc344107589dc409044b1 + 1;
            Ie8a61b138cd654efb72fb596046bc9d2b50c97e34d4a27a1d457261b4f8a9fc6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I519df6e33d8ef22d52e32b8119be2aaec1f50dbccc5d79dbae0f55ceb6cb8f18);
            Ic15cf2e839052d47aa87202bae190c69e5410914d9e00120099307d6f7a663c5    = Ie8a61b138cd654efb72fb596046bc9d2b50c97e34d4a27a1d457261b4f8a9fc6;

            I9b4f99332934a592b74d60329e811e336cbc4f6af94e1e7585e47c8096b05b3e = I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347 + ~I0c851ecaa50ea3e1769828a7f51da7a8c3b0c0a11eb9002b108693f09e60667f + 1;
            Ied33aea50e5d0112a854d4877d3bbcb4bc21b4ef75e4b120c0104770d83aeec1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9b4f99332934a592b74d60329e811e336cbc4f6af94e1e7585e47c8096b05b3e);
            I74677cda9719646b1c842acbed5d3b13462ef153d0a8907019b2553c808f84c6    = Ied33aea50e5d0112a854d4877d3bbcb4bc21b4ef75e4b120c0104770d83aeec1;

            I513af0998e26ce841c280947d55c670808280391fcd874412081722d9a9915c7 = I45c3294dcbfa1aeb134d8c83c176967fb10d518a3567e1816276650e72c5e347 + ~I09e3897931014e7bd9540023eb8fe1097e36eb5c51db24357b492a132c3a8805 + 1;
            Iac16fa27063df4a80f23e3757dd21e3116aa16f591d7e80e7079571e2f2ab6b7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I513af0998e26ce841c280947d55c670808280391fcd874412081722d9a9915c7);
            I4e0c405b4f7107ae7d9a35eff8fc48672c1ff35ede5dcbaa4340926c9d9e65d4    = Iac16fa27063df4a80f23e3757dd21e3116aa16f591d7e80e7079571e2f2ab6b7;

            Iea8434e90fef04642cfc1cbec886240547c066665e40258a1412ba69225faef5 = Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9 + ~Ic3ea8409cfacf50e41b97c65b0440348d06b8f196001ba1fda6348071b47dd23 + 1;
            Icd7c491a614817929db2d44117b8bdd384f7d9387d4bca021959efbc58fb7b3d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iea8434e90fef04642cfc1cbec886240547c066665e40258a1412ba69225faef5);
            I1db1a5d4e476af4fb7bbf80331760238438096833616b30904a4b6fbe0057e63    = Icd7c491a614817929db2d44117b8bdd384f7d9387d4bca021959efbc58fb7b3d;

            I4fbe4e6bbc2d22f919e4642a3f6e950358f3ad9c6ee0d7997ed355969a8023b0 = Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9 + ~I99c4a78ad7af699907cae52326915f18ac1a2a6f9d99b2aa71c34d10fa78fbce + 1;
            I9114e7211d58cd46c3e15d782c0822ef34b1436c74a1842a8af9abddb2117c7c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4fbe4e6bbc2d22f919e4642a3f6e950358f3ad9c6ee0d7997ed355969a8023b0);
            I083b6e833d8b3bda9d56f159a5e297305e44fad9f2024a3204c6e5b7afca9405    = I9114e7211d58cd46c3e15d782c0822ef34b1436c74a1842a8af9abddb2117c7c;

            I83d1b40ee8296b6a8bbf02a87c6f077c2230f2e8875c679642386b74c055dc49 = Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9 + ~I4878199f761be0332cf7d653cf1e73cd52f938bf9ca0f32724d499765f313d46 + 1;
            I8fb26cd47b8f0da1d89b9818685edf5f9c9776e0df5beab4ebddd0e3c616c7e2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I83d1b40ee8296b6a8bbf02a87c6f077c2230f2e8875c679642386b74c055dc49);
            I410bc8d9b13d79713c47cab785cae1ee4db55ba3e7a207519bdbc646dfa815dc    = I8fb26cd47b8f0da1d89b9818685edf5f9c9776e0df5beab4ebddd0e3c616c7e2;

            Ia70f5a20618894e74f792df1afb11ebd1e590400cae3cb09cd1754416a26bd07 = Ib07c5746b957e7a7dba26c45d06cd6e60f1bbf776a9a28142663bc1ed0f854e9 + ~I674ac3fcd5872491a3c412a02e367a9c29e4dac14a8ffe8b6382c60a29fde8aa + 1;
            I207e7042b2c0cdcf57378c651ebe265368b8b922f54a33e5b327d55548833526 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia70f5a20618894e74f792df1afb11ebd1e590400cae3cb09cd1754416a26bd07);
            Iab1ad3fda6ef48c15a116045600ab96f057c4e2769b1736742ece54e049a9884    = I207e7042b2c0cdcf57378c651ebe265368b8b922f54a33e5b327d55548833526;

            I8b2a2914ad57445d7e6409d706a2d5c9cdd01b8f7163d153c1647304ed71c1c4 = Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf + ~Ic9e13fe7c29048953ae3698eb5d214d6b71367a78bf1042dd6b58064a6cc596d + 1;
            Ic3a032b15228b0da60d25deecdfa1ec1898c483d70e6d08be8f89248292b2fb1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8b2a2914ad57445d7e6409d706a2d5c9cdd01b8f7163d153c1647304ed71c1c4);
            If01282d291c85bcab01b47104be9ed13915609c85c61d979b60b02847a685e4f    = Ic3a032b15228b0da60d25deecdfa1ec1898c483d70e6d08be8f89248292b2fb1;

            Ibdb714449c61293321fdff34d19ff92c2a66cd677739a387bfbbfeb482a17aa9 = Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf + ~I072f20811fc3b3515b7794a416e5ba39cca6a9579de36442fb39771729dffa8a + 1;
            Ida75a6cb83f408b8efb2b6a75c221c6d3ec50c673bad1265d400a39da9eadfee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibdb714449c61293321fdff34d19ff92c2a66cd677739a387bfbbfeb482a17aa9);
            I2c3551c0a960cbdcab2b802148c759ca7c8dc401d98b251d9ea21d6de16d3bf8    = Ida75a6cb83f408b8efb2b6a75c221c6d3ec50c673bad1265d400a39da9eadfee;

            I6640a4310bb1a9135eff3995cda6d740dfb307d44c62603190f7cbfbfe285718 = Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf + ~If4f8191d57bfd0311981d36c3836f8da526830c6fe2dae5933650b290075ef17 + 1;
            I9d246b2101b98789f6c8b328fb0184f6d02065d04c6935ef49dd5baf259c1e54 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6640a4310bb1a9135eff3995cda6d740dfb307d44c62603190f7cbfbfe285718);
            Ic7977549066f72a2e4c0d91c592a5d93a2a64fd1ac48cafd6f0f4600912f3fc1    = I9d246b2101b98789f6c8b328fb0184f6d02065d04c6935ef49dd5baf259c1e54;

            I13d152d9c14bf7e9d0d71bde2846f80bafd4553400bccebd37d850034d62514a = Ic347bdc15bb8fccc7f3953a9f323928c0bfb29e262b90ec48981e57c0aef3caf + ~I9ac796f1901c19aeab344ea2c785af3ce41bd23dffe88b1b5216f8f8c0b16e40 + 1;
            Ibf193fba82d63a518161b53b8a23b3fbd93fbdda529aa080fe932edbea6fc57c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I13d152d9c14bf7e9d0d71bde2846f80bafd4553400bccebd37d850034d62514a);
            I08c54adda4326fbc5985605f17f5b1c47ce821476ba25053aaa7449a571bf33c    = Ibf193fba82d63a518161b53b8a23b3fbd93fbdda529aa080fe932edbea6fc57c;

            I3c0e2c1dc0aee993679368343156a72f56d55c38911596cd28c13fdbc68ebe53 = Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2 + ~Idc5ae39b0c3c764ed6d9b7859b7627b97e24c2b4df7d97229a88cfc0c22ccd87 + 1;
            I351f23377572c7cc4bcab051aeda29360f51b89eb290bac8e484fe05adc29065 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3c0e2c1dc0aee993679368343156a72f56d55c38911596cd28c13fdbc68ebe53);
            I74a65dbb33c6088646be4339ced1e6167ed3c67fe3f520e10d4fb2c96358ce62    = I351f23377572c7cc4bcab051aeda29360f51b89eb290bac8e484fe05adc29065;

            I76208cd61a51a2330f9d46b67e0b036db6de794a34a380a75ca6f60439344546 = Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2 + ~I9e8877d4beab63d4bf103c07e1cd9330daccde2cdd266b2942f56b2a8e8a926c + 1;
            Id85a42323f6615cb44efeb003b9a3bf7309bc463bfe55bbab0aac732f99c975c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I76208cd61a51a2330f9d46b67e0b036db6de794a34a380a75ca6f60439344546);
            I378dc69acacc690da268354f08a9f1fd08b11a899cd2253c2cca3c979245a06b    = Id85a42323f6615cb44efeb003b9a3bf7309bc463bfe55bbab0aac732f99c975c;

            Ib95f8920a685d0da3fc07ac7ff3a19ee1fd5fc65dc4b6db141a709668c2d579a = Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2 + ~I6aaddd1a59b6e96dd8cdd4a57d8fc03132dde1c5b0bd06dd6f0a240c2a04f947 + 1;
            I77385a4a50aa8eead5b897d5c076357ef507c90dbfec7d442ff728bc20b90048 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib95f8920a685d0da3fc07ac7ff3a19ee1fd5fc65dc4b6db141a709668c2d579a);
            I8519733c2d4de3643ecf515bc788e665d7661c947a6532dcefce59b255fc05c5    = I77385a4a50aa8eead5b897d5c076357ef507c90dbfec7d442ff728bc20b90048;

            Ie5269d77c7963028196afc5b429c121674eb881ef85f0c30e06bf3e0b5b3a7cd = Ic6bb987782bbe2823102ba9a4c8f81aeeb59518b429448719adc9fd3fd6549c2 + ~I0d186e0127f200b704a4585b2fc43ff1a9ab19833a90ac881abde94b2da89376 + 1;
            I6ac9c9564bd70c4a8c9a6a76450dae9f55e8008338bb7d9f85f52e06b17ba7fa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie5269d77c7963028196afc5b429c121674eb881ef85f0c30e06bf3e0b5b3a7cd);
            I2b3f1cb9e25ac68c67abdee581e7dbb74b039b9f1f04459e3a4049769f27c474    = I6ac9c9564bd70c4a8c9a6a76450dae9f55e8008338bb7d9f85f52e06b17ba7fa;

            Ied5144deb00adc8fdbd1024c051f87a6725bd5211f5d24ed9d965ac7bf0dbdab = I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 + ~I18886d5e45fe8011ebcf9a20aebf875a01f1b793a54ccefdbe44a896e92cb0db + 1;
            I02325f467c1fa16e231a42dbb8e973427b2a4c081fdb336e3f3838d5f7a7061b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ied5144deb00adc8fdbd1024c051f87a6725bd5211f5d24ed9d965ac7bf0dbdab);
            Id79e7da27c2a195d433419bcc0481ffe12155390f0a10ac6be75723cf2ad53f2    = I02325f467c1fa16e231a42dbb8e973427b2a4c081fdb336e3f3838d5f7a7061b;

            I604e5b545ac6c440263889210560ae82bc9dc0f3717b456ea8844cdad1813c2a = I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 + ~I786cf639910ac9a90b1abf55f9e3b66d87c4bb98a2c8e38142969ee5aefcf6d4 + 1;
            I389ed2df5d3890d3c2f628edb1a043d51a972de9cb338f32389788f5acd90028 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I604e5b545ac6c440263889210560ae82bc9dc0f3717b456ea8844cdad1813c2a);
            I9aa3880979a20743da2aa753686d0ecaf0702008920d80af34d834ef1e2249be    = I389ed2df5d3890d3c2f628edb1a043d51a972de9cb338f32389788f5acd90028;

            Ie802b6bc444bb7d279d93b810491f7dd483ceaa3c122368578579700a1723669 = I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 + ~Ibee0b890887202cb33c8fb07639c7bc536951ce8e661d561d7e7a7355db5f9e1 + 1;
            Id9e38d40473faaf687741f97150071792a45a4926ec46762a3d1729e7b1d7111 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie802b6bc444bb7d279d93b810491f7dd483ceaa3c122368578579700a1723669);
            Ie591b9c2c777632b671f8aa86f6befb3d02e16c23329cbc7c07438588aea4c9b    = Id9e38d40473faaf687741f97150071792a45a4926ec46762a3d1729e7b1d7111;

            I17e1e63cdaf581226fb06f909c0c75f2ceeaf45e1ebe93127d22a0ee6ca7e8b9 = I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 + ~Ibf0c6b2fd7ba6e86f7cea34ea8434ec5353399651fae6f00cae29cfd32174563 + 1;
            I49092cce392bbf2662076c5d86322bf8c9c77a778ef3893fb58e9b08396f2d24 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I17e1e63cdaf581226fb06f909c0c75f2ceeaf45e1ebe93127d22a0ee6ca7e8b9);
            Ibaccfedeb751c2506a2342df2f75fe492accc5c68614fcb90b4f5c332c088808    = I49092cce392bbf2662076c5d86322bf8c9c77a778ef3893fb58e9b08396f2d24;

            Ib106ae5d2b37f2048bc3c493b80c76048d8b5c4e1ebedf0cdcc6bf20958f39e9 = I852dae977146864ac9ff8c1f2a25769808afb6c8b8a04924d8810c1d7aa400c3 + ~Iae8191d31be3785db5d8e5d328fb2d96b0b5d5ecc7f9d14f0bdd3f61a9bb6781 + 1;
            I5b1f9cbdb5bf4a096a6c8bcb4db57912d6cad99055ec47831516d612f7129dd2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib106ae5d2b37f2048bc3c493b80c76048d8b5c4e1ebedf0cdcc6bf20958f39e9);
            Ifa134df77ff670a0cb559c384c786af4de916cea66ca13147d43f4030d474d0f    = I5b1f9cbdb5bf4a096a6c8bcb4db57912d6cad99055ec47831516d612f7129dd2;

            I6da36192889d17f86e9b385d553a116e1315dd88657c56f92f4603cb75e6de4f = Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b + ~I5bb2c70350634acbcf64debae260225ea2ef5b67ce5d03f38d56d3db9de687f5 + 1;
            I81a866e481435399f8705efd8f264d7419c1acdc086298638158f4d75202b567 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6da36192889d17f86e9b385d553a116e1315dd88657c56f92f4603cb75e6de4f);
            Ib378be3532348ccba868d918209ee3f013c1844044c8a93467a93c3463f7a36c    = I81a866e481435399f8705efd8f264d7419c1acdc086298638158f4d75202b567;

            I48595b1f5633b6439ad79fc3c53fa5da509c15abaa66b7b6aae7fe56e8b560ac = Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b + ~Ide94701dd8ad54a630c6eadc44221ee5786180f247fcaec8a7787f25c4070968 + 1;
            I44c742e7ad2e3e18153ce9b645fc21efb4e3016f063b05a8bc1825b05a303374 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I48595b1f5633b6439ad79fc3c53fa5da509c15abaa66b7b6aae7fe56e8b560ac);
            Ib85e84ee2add613edb76e2321f7a5d6b4de3be9b1ab97905b5980277ed273dd1    = I44c742e7ad2e3e18153ce9b645fc21efb4e3016f063b05a8bc1825b05a303374;

            I7ff33f6abb8c5ed6800e5c1c58b974df6d1359987f819291202ff2413494aaaa = Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b + ~I31d4c202b8434aacebdaf5a60c34d7bf3864a5a7c4707efbd1cc3dd82a9ba59e + 1;
            Iff70805870814e2f1b8de2513c56a30b9e6194298cb863c87a6e75221c8ef1db = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7ff33f6abb8c5ed6800e5c1c58b974df6d1359987f819291202ff2413494aaaa);
            I10ee9fd16ea681268e4bcdcc30b515d990dc30d3fd41e059e9f1dcc80042ae1f    = Iff70805870814e2f1b8de2513c56a30b9e6194298cb863c87a6e75221c8ef1db;

            I914341a688ccdf40369a1abe1fe5bf72b3d5ddd306f81d3364e2ed4e03970149 = Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b + ~Ia7c03e6396e5145d0027d0963c1f8b7068636ee262fe31aa442a5512e0d4e99d + 1;
            I6188d9b90b4bb155ad464258b5d3ae28e757f4b3ca73453ac4ab3d6cfa8e6643 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I914341a688ccdf40369a1abe1fe5bf72b3d5ddd306f81d3364e2ed4e03970149);
            Ic33e33bdd936748553ff29221e983dc115121fc84bd1a2799a3da8120be82c04    = I6188d9b90b4bb155ad464258b5d3ae28e757f4b3ca73453ac4ab3d6cfa8e6643;

            I3e201da437cb62d4d6db5d7fbc655eb26c3a1d49dc3d7ec08b65b4979eaa76fb = Ic54ba117e42f2bc236913907b5727aec583ab5fdf1cb0926091f3cc098b8269b + ~I4694c593512d9d84542af4ca5b0f3022f9b1433d7d6435ffd4b1e53093bf4a58 + 1;
            Ie2603a3570f686ace17fc46e9c5190f79e2cb32b4e6d3c39c26265951b22dc00 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3e201da437cb62d4d6db5d7fbc655eb26c3a1d49dc3d7ec08b65b4979eaa76fb);
            I0705a3be469f22a69c0c4d2366fd0eaee02065685349db5abd81049530fbf842    = Ie2603a3570f686ace17fc46e9c5190f79e2cb32b4e6d3c39c26265951b22dc00;

            I59be2b7a5e95aa90e3d27275839badf750e2f713ff498aaf28bd202039ceb029 = Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 + ~Ia249a4e7b5c5f1f4458d969c346e560a28969f33c9b0371c6bb21776d319afcf + 1;
            I97a0471ea526aac1fb508c6cf38c387c6afd71b9089e63470279445f4ac8f7a0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I59be2b7a5e95aa90e3d27275839badf750e2f713ff498aaf28bd202039ceb029);
            Ic0edcffe7bf2caf311b42675297cde79af81c022f660757cdbed53dbf5c04eaf    = I97a0471ea526aac1fb508c6cf38c387c6afd71b9089e63470279445f4ac8f7a0;

            I634697ab8c90d12c2b2b2a65d6545a8de51ddf645111a26570ecbdafe71644f2 = Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 + ~Id4182b8f05992677e12502bcc058d967481d0dc2c9c4731b657f04696a5b5bbb + 1;
            Ia2ebfd7cea041d6ce3b26d85588f2113701cf7f6970206eb4ea2001c3ab0f52c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I634697ab8c90d12c2b2b2a65d6545a8de51ddf645111a26570ecbdafe71644f2);
            I600367d873f901e6b7f92a4f9c0ac92c9f8efa6da1d6e6945f83b863e8bb8519    = Ia2ebfd7cea041d6ce3b26d85588f2113701cf7f6970206eb4ea2001c3ab0f52c;

            I300f54df5ff39044592d1e17773b678120282a58df676eb35de5794a0fe9e562 = Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 + ~I9dd21c6b63d36e7dde6f3133ab04263a47559b648e8717de7065e7f140911d3d + 1;
            I41854c843f5042d94267a6b9d374dd0f5c46fcb45df0f40b587aca943f7bb396 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I300f54df5ff39044592d1e17773b678120282a58df676eb35de5794a0fe9e562);
            I8e30a7f3eb36b84c9df9d59f6164c757c8612fb12567ddfd03c32388af750bb6    = I41854c843f5042d94267a6b9d374dd0f5c46fcb45df0f40b587aca943f7bb396;

            Idf7a27915130178e3aff7acb7a945422a7955b81a491f1579d88f01797270738 = Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 + ~I9244711e562e8ea7e5e0de1921bdbbc5b64363d51d121922f441d8f36e949c69 + 1;
            I542e912b5cd0969a23f6d60abd1923cf0d333b3f20df92061570f156f395d756 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idf7a27915130178e3aff7acb7a945422a7955b81a491f1579d88f01797270738);
            I8d123ed314ee10c10f04151727cd5ce1e836c01f0f8143285b54425633591008    = I542e912b5cd0969a23f6d60abd1923cf0d333b3f20df92061570f156f395d756;

            Ida7fdf0874cf846834b903eac34741e8b445fec4ac30ed1451ad758a50d90aaf = Ib554d0a4108936aa437a8ef2150d3d6824d974e011edc1cd78fcbb7cd0bb2485 + ~I78c5059e528b7671e27f847d6042b3fa707258c664749d857004679c6ff96a73 + 1;
            Ib49bc31787442badfaedc737b3e1e4014bbd7818595fcf9cf42f23dafe03fa9c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ida7fdf0874cf846834b903eac34741e8b445fec4ac30ed1451ad758a50d90aaf);
            I0ae31ee6a1c597ec90ca13dd69a651079d801c279292523953428af55188ddea    = Ib49bc31787442badfaedc737b3e1e4014bbd7818595fcf9cf42f23dafe03fa9c;

            I6ecf3391cb1fa3dd5e19dee9f9d10088818c528a1feeea04869723baa4e0f2ca = I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 + ~I7efedd1a063df95cac921f7cea9ceea1ddd1afd3a70289c50ea2a4807310518b + 1;
            I3069d559ed47e3e17dfd391829deba4bec9932d5ceaee52ba24e585c3ca750c4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6ecf3391cb1fa3dd5e19dee9f9d10088818c528a1feeea04869723baa4e0f2ca);
            I7bbfdff59068ad7e527ada31d96fd47cb737e6b7ba56b1b2b9e522fe3a63a954    = I3069d559ed47e3e17dfd391829deba4bec9932d5ceaee52ba24e585c3ca750c4;

            I7a0182d704153bcdbc1bd5927e4a45326e90a16a9a962183407f29753db6a41f = I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 + ~I598f53ba5c7ffa41f21af94375843b0b7a911670719edc80705508ae32ac0ddc + 1;
            I74beac54df2553b0529872dab3dc06224f214ce3e1028033e9830a31dbc6b036 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a0182d704153bcdbc1bd5927e4a45326e90a16a9a962183407f29753db6a41f);
            I09001eb04237069c413098f07bb41538c6d39b0ac000f175d61ee3c0b47cfae2    = I74beac54df2553b0529872dab3dc06224f214ce3e1028033e9830a31dbc6b036;

            I044b0c28219d5422e97568291ba0de670fbeb09c83f1eb2943afe0a4be000651 = I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 + ~Icc14287e817338eea415b9f8dae2527d6e71853a49869ea829d1b51aa7013dab + 1;
            I2213f69a2b20b811c1ffe8ddc5b7a0c31df06430e2d02679663fe31305bb6c87 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I044b0c28219d5422e97568291ba0de670fbeb09c83f1eb2943afe0a4be000651);
            Iddcd6e6693d5f625ba82ec2cdb0a93ca1826dca4989d19221c8127513648eab2    = I2213f69a2b20b811c1ffe8ddc5b7a0c31df06430e2d02679663fe31305bb6c87;

            Ia82e0334a1b24c5ff4ee87a2d117c3c7301aae9a45e4704b36436f166435ac5c = I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 + ~I81c33c11a5d878aea61749e54e68c024fda21f27f7f4fcf45e5b042e8ca4c3fa + 1;
            I85dd7ff4d35dc1bfbca02c07a3f89560d8b9f8f10c9f28ed1709e4e00583b5d7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia82e0334a1b24c5ff4ee87a2d117c3c7301aae9a45e4704b36436f166435ac5c);
            I89df294963327dee66a931b858b05dddd97e3fe4d048ecbfaa9c15e28c57602e    = I85dd7ff4d35dc1bfbca02c07a3f89560d8b9f8f10c9f28ed1709e4e00583b5d7;

            I1cf673d7825554846ea143f7954ebee1453bd097d3051107dafefd72ff05ea29 = I15dc05c2cddd067ea8e5dc4fc53a918341888c1fd1beb5fdc6d8f77523942fb0 + ~Ic83ed3610853814d7c9d6932b644f9c924fec7d67e303160a3c5b99c625634c0 + 1;
            I385ea910caf7d0563d1214dbd983b37fd5cceeae24015a0b4cc253612b316c22 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1cf673d7825554846ea143f7954ebee1453bd097d3051107dafefd72ff05ea29);
            I1f0110f45df674628a1a02cf01dc58577628dd88049b93ebf02b5c4143781ade    = I385ea910caf7d0563d1214dbd983b37fd5cceeae24015a0b4cc253612b316c22;

            I3972965d0045633d150172c2debe5d89bc8aefb8473b1c697d26accceec1b2b0 = I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 + ~Ib91519b86b75cae1ba5b32dc531cae021a01350f4e184d39373bf5553f89a7f8 + 1;
            I5c1a4f9167a1ddf22a7642545eb95954fe17112c630b62d9e95f899783de734b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3972965d0045633d150172c2debe5d89bc8aefb8473b1c697d26accceec1b2b0);
            Ib0995588ac28564326a4dec88344ddd733075750fab9f4f8fec64cc91b3b48e2    = I5c1a4f9167a1ddf22a7642545eb95954fe17112c630b62d9e95f899783de734b;

            Ic4b7ca6006b1fc68a4e04414ba1c587cfef6136c1ce1702fd09cfc264ec96920 = I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 + ~I42295332275fc6fcb94c042fbe6b48d3d03038fc27c535c7e63674f58da60bf0 + 1;
            I231bdd513a7d05321aa7ee4d1bfc4b59edcc82ae92b1e27403f0773bdea92e92 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic4b7ca6006b1fc68a4e04414ba1c587cfef6136c1ce1702fd09cfc264ec96920);
            I3a2ddd5962242d66fa4b8bca39a81765dfbc6c0b6b012ee42329dcdfc12ae9b3    = I231bdd513a7d05321aa7ee4d1bfc4b59edcc82ae92b1e27403f0773bdea92e92;

            Ib4e8f9db85c1b658d5be48822318c0688eb41b8d011aa69d188be0680d53de8a = I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 + ~I3db60bf522be36d36bdcc35d1d5da9cff2db6e8f89b179726fabca1a7c67b255 + 1;
            Id0b5d2604bb5b289b82f24f9e91c4669cbbc04d0e3d79aa18ebe3dd27374837d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib4e8f9db85c1b658d5be48822318c0688eb41b8d011aa69d188be0680d53de8a);
            I83cd839beef638f212312a0093595ec3d71dc80e240aba892f6404de6d614bec    = Id0b5d2604bb5b289b82f24f9e91c4669cbbc04d0e3d79aa18ebe3dd27374837d;

            Ic95ac5beb10ecc57a9669b74ccc04b6d5327b39b5a085d6937c1ceebd9cb480e = I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 + ~Idfb0ecafd00955b66bbc43f1585659b2fd82fa239ab0274450da985354bc4c14 + 1;
            I44a2a1b5e4fefb27d702cad5d65609674fef85f845b8cc0da1c6122c867d9317 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic95ac5beb10ecc57a9669b74ccc04b6d5327b39b5a085d6937c1ceebd9cb480e);
            I3420837ce14103293c9ee75848088cd144ed5b975add2adfd479ad10eff552ca    = I44a2a1b5e4fefb27d702cad5d65609674fef85f845b8cc0da1c6122c867d9317;

            I32d8bf76f6a512a10f6231445299d254d8fb22c51f6edb2ffb1c69b44804cf47 = I044596abdbbf059c1c0685d99eaaf0162da286cfc2784c0c0697b73c17ffe4d5 + ~Ie33f8884c8fca47e2055b28f4398f3207f7ea20f8d0858d2a0699ef2da5a8f03 + 1;
            Ic3e639bd8b640b9a08515fb88cb35f8d263c8b4bba6612a800b303bb21974a4c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I32d8bf76f6a512a10f6231445299d254d8fb22c51f6edb2ffb1c69b44804cf47);
            I641204b71e0368d174adf904e08c12465fc7a18e1adf1372e1649efad206ba0a    = Ic3e639bd8b640b9a08515fb88cb35f8d263c8b4bba6612a800b303bb21974a4c;

            I100ae29be1331206365e7953c6d6faa026c8c4dd25311560d51afdf2db866849 = I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c + ~Iecd27d9347b5f52e83b7d0fbf7e51de4a3711cbece5ee265b12663b77b58914b + 1;
            I85f4e180cb842542efe4294bad76481afdab9af7982dbc049af943d3fb23787b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I100ae29be1331206365e7953c6d6faa026c8c4dd25311560d51afdf2db866849);
            I10bd3ad7827da7bbb0e1170d7e495b88ab6ac55e0421b4f208f5c1ccd722198d    = I85f4e180cb842542efe4294bad76481afdab9af7982dbc049af943d3fb23787b;

            Iab0de1945cb02c4493fb064c1efb72f4e5a0483452c5c29276c4c7e1deb5087d = I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c + ~I97f8487b89684c5c6952770b0468738f72682d6230be6a5a31a92fe50bfb239d + 1;
            I2d2a89c4664389a9d5615140b32a9a994b150385e23a1ba81bf0823ae34ff5b5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iab0de1945cb02c4493fb064c1efb72f4e5a0483452c5c29276c4c7e1deb5087d);
            Iee26e4077668d0e7329068693c4279480b26e4f16adb0161c8e7f87de802a14a    = I2d2a89c4664389a9d5615140b32a9a994b150385e23a1ba81bf0823ae34ff5b5;

            Ib13e8ac762b6740072f1415df276b0ef0703a282b8dd7268638bbdd370a05e90 = I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c + ~I42336bb9a452e51859fbc836c4294468aced58a32a221057096f5119d459edc9 + 1;
            Idff2c2e52bd3a5b88eb4da782cd2bfcf9621c26033b6643a8ab96749a80c9fe6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib13e8ac762b6740072f1415df276b0ef0703a282b8dd7268638bbdd370a05e90);
            Ia8e573753ddee4fe18b1f9fbafcd135efc7fb7e7eec52e45b5148b0dcf346050    = Idff2c2e52bd3a5b88eb4da782cd2bfcf9621c26033b6643a8ab96749a80c9fe6;

            I7b4e445b2a01b541d52ab461384c1bbb27cbd46e82cd7c401f4350a5e468d237 = I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c + ~Ia50c90193d9c7ee51018451884df0da92f138710bf95fc32e439b39bea3f3b01 + 1;
            I13ca4018c147e25a38463d2fa98d04240b46a846f1b8b13f69b99942a4b2539c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7b4e445b2a01b541d52ab461384c1bbb27cbd46e82cd7c401f4350a5e468d237);
            Ie8e89070910f06608a4df5951936faf465b4f235d92b3cf8a3820d03bcaa83ed    = I13ca4018c147e25a38463d2fa98d04240b46a846f1b8b13f69b99942a4b2539c;

            I70948947c6b4777cf695a6ac2097443bb59059da06704ae1f5c84b42144e4a54 = I3805fae004899b31e29b7d8122b5a1f3e9974502fbbdacd6b2d05754ae13013c + ~Id140833a04f0b4b903ad4e99046b17f76d4c405703fba227d36342b6f1fdbd08 + 1;
            I45e1276a5f5af744327fb6f85b50f8aa50bb442469cbda4ba869adf5a8d0fcbf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I70948947c6b4777cf695a6ac2097443bb59059da06704ae1f5c84b42144e4a54);
            I1a0b36a215887b4419ebcfbddb0ab8b4b9b21c4643051db135c9d9ee53c6bb3e    = I45e1276a5f5af744327fb6f85b50f8aa50bb442469cbda4ba869adf5a8d0fcbf;

            Ie5e4bdbeb1b832d35e7974194a251885c1bd525aa0c434055cf87fd540b224d5 = Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 + ~If81604260c143a45d248461563d4d94edd94bb71d791a637dcd30c5c0cbbb965 + 1;
            Ie63f997e6206a536a5e45901da6593c5c49645e6cef643846980c4e2070091b6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie5e4bdbeb1b832d35e7974194a251885c1bd525aa0c434055cf87fd540b224d5);
            I84694b26e240bcc3e7c9b224ce3c2f5891fb546a4fc11e4597819fd9827c3105    = Ie63f997e6206a536a5e45901da6593c5c49645e6cef643846980c4e2070091b6;

            Ie12a5b8c714d7783eb66355736714fac95237a0f821071b9b379359f5d6665f4 = Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 + ~I3e014fe75658214d8ffa60f966549b131bff6a16020d7858523ac829b0126838 + 1;
            I275a2a54f37e000edfcc6f35cbdf2ab6c2a28604ce2e6dc31d6430693c2ddd4a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie12a5b8c714d7783eb66355736714fac95237a0f821071b9b379359f5d6665f4);
            Ie69f3ad2e3dcb172e525302a533963ab9a2a08af8d1ec71e07d0946d393c056f    = I275a2a54f37e000edfcc6f35cbdf2ab6c2a28604ce2e6dc31d6430693c2ddd4a;

            I1b5dfb756878da24a1f7528fe4a866bb750e2dbede6da8548653167c555ea8b0 = Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 + ~I0a22f1dc32c83db6603459232e78078eac21f865aabe0b9a03923e63cea874ff + 1;
            I5848db5ea2fd0385e583946224dbe078419a4c9684d15157ec460537baa30d91 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1b5dfb756878da24a1f7528fe4a866bb750e2dbede6da8548653167c555ea8b0);
            I6e0e1c5361317aa91a6e54e23fe2585744a1ec47fcb2412ed152b660781c7832    = I5848db5ea2fd0385e583946224dbe078419a4c9684d15157ec460537baa30d91;

            Ib07212f6fae72454c08283293951d3fff4ff77cf5455f98c5a85218c07a897dd = Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 + ~I157157e9b85b39f2f22c57c4beae22472512ec83319dd9ac30075b4266761031 + 1;
            Ic0dbeca58e8f490493dc5672f4aeea9b98fb9aa4aedb922714f3aa21a4836223 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib07212f6fae72454c08283293951d3fff4ff77cf5455f98c5a85218c07a897dd);
            Ia338a53ab734049efb28655e209908f1fd2c5d19f8056463d711cc1e50dde602    = Ic0dbeca58e8f490493dc5672f4aeea9b98fb9aa4aedb922714f3aa21a4836223;

            I8af68a180894ba478298d5c06025d929869476ca01e3bee443254dc410fa10e4 = Id0e4a59852289b002e9d0758c2edcfb6d3ba145f40ac1b5b93b2143d5a0dd439 + ~I90d7a3c4ac0a18444eceec2569cae3d5dcb3d33d2e46c329068b0d35ad063971 + 1;
            If7363f53cc60b20a744ae33ca65adb0345b104fbedfc2ddb5bb00b1dd50bc13d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8af68a180894ba478298d5c06025d929869476ca01e3bee443254dc410fa10e4);
            If63dbf3e3c6000184af28e72b5f2960f6a376f509d5693a96d2ab9f92ae7b237    = If7363f53cc60b20a744ae33ca65adb0345b104fbedfc2ddb5bb00b1dd50bc13d;

            I9455f55f4c34a937845af7d359cc07d1976a1fb4f3a9e7a262316e137b241b6a = I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 + ~Ifd8d2fce7b2a1f0fa487e5be6c007a21b5af1d79da5447d461cd37c189e43561 + 1;
            Id8ae67d7680689c7007d27eb5af9c5bc1277025b9ca78c804632ce105d41fb08 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9455f55f4c34a937845af7d359cc07d1976a1fb4f3a9e7a262316e137b241b6a);
            Ib89d5800576f979f189d88e7976f8d49b8470bcbf6b365f7cc6031735e3adb4a    = Id8ae67d7680689c7007d27eb5af9c5bc1277025b9ca78c804632ce105d41fb08;

            Ifaa7c357c28b482e992040ba6eb62623f7ca590303fe66b20480f8eca1b79974 = I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 + ~Ibe646b6da0465c3fb411afc4e03d45f553cf91e67cbcd46674a0051ac1092e30 + 1;
            I7f21d46e9cf807c74d37e3d383186daf9288e68431e128ddf72f9f448f671ad5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifaa7c357c28b482e992040ba6eb62623f7ca590303fe66b20480f8eca1b79974);
            I622321198c6f868e554b595d1e1616dd63ad46a80c33bbe896df9b6558418ccc    = I7f21d46e9cf807c74d37e3d383186daf9288e68431e128ddf72f9f448f671ad5;

            I48fe5a4d8cc9de9df457625de0ccd81303342c2653cb9051ac93358c46aededb = I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 + ~Ia28734d68fd59a227094e3d5643b87d918753610e867c1d047d8878bd9a46be3 + 1;
            Ie9f2f5a180ba3e3b29c209d7e3c735224fab3c309f2dc627046d864a58f42897 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I48fe5a4d8cc9de9df457625de0ccd81303342c2653cb9051ac93358c46aededb);
            Iafcf26b8f2df7719a0b660b41de28c5a325e50d75382579e53aa9d065bd81cbf    = Ie9f2f5a180ba3e3b29c209d7e3c735224fab3c309f2dc627046d864a58f42897;

            I4a2a60be7efe872271b328a84bd0394ce67c2d59ca77082b5a4ff71b5b5f2707 = I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 + ~I7fed914efeb5727bba8c1dd0a5cab385a750a2cd9215923b596d1ae914639761 + 1;
            I6dfe9c7c9935ceb07f55d4fcf7feea54e13050347b5991fca21d79ad74608aa1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4a2a60be7efe872271b328a84bd0394ce67c2d59ca77082b5a4ff71b5b5f2707);
            I859639da611c77242efe899343358a650652277ea45277d9792b619196c66a1a    = I6dfe9c7c9935ceb07f55d4fcf7feea54e13050347b5991fca21d79ad74608aa1;

            I51a55a7f067596679dc3e69c0d0fe9c92b776f65ed24981709079891bb7d0edf = I1af7a70e18c25fc571a7f3542ccba9b01f0c402ed7df962a35c84d79727ab451 + ~I5c7c7df860c87ada06c17210746ef84d27aabaa26e9cad20397822629716d4a6 + 1;
            I65290aca857afa1ad9b6aa754dfaaa0671d173c7b3d9fab7cee9ebb973b32862 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I51a55a7f067596679dc3e69c0d0fe9c92b776f65ed24981709079891bb7d0edf);
            I2899ec4e420edc766050ec0042965f87c79455271a54ba7c947e94d37450a033    = I65290aca857afa1ad9b6aa754dfaaa0671d173c7b3d9fab7cee9ebb973b32862;

            I4afb194348fb5347cbed837090c3d94bf4a27f44202d58ddde64915fbf8c7bf3 = I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847 + ~Ia49277306313784711d5d8ff63e6a0a77d3fbae050dc1089c734c826be497dcc + 1;
            I8748f772ce4e677c9220c1fb10521d69acb830ffb623c0490c1410b515445dbc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4afb194348fb5347cbed837090c3d94bf4a27f44202d58ddde64915fbf8c7bf3);
            Ibb256fb3d4bbe6ddc65378ced36e01255d8164d29755891e06fbd4caf2a290cf    = I8748f772ce4e677c9220c1fb10521d69acb830ffb623c0490c1410b515445dbc;

            I7f468cc83b7f0da006d4b41ef40e5bc4e84e7ea6811d5d66b61690d80c82ffb4 = I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847 + ~Ic1034fe189ea09f2aa3b69428828a2b7dbfe9389dcf48dbdbe0f15b9157f7c49 + 1;
            Id6123d9000c37cf18ad9bee82fef91900b7ee165a1841b5a4d23af27bcd0fbbe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7f468cc83b7f0da006d4b41ef40e5bc4e84e7ea6811d5d66b61690d80c82ffb4);
            I60f4bae66121b814e2faa564c162bccbd2ef0a73bcaf10c3c78e30ff2edcde4a    = Id6123d9000c37cf18ad9bee82fef91900b7ee165a1841b5a4d23af27bcd0fbbe;

            I73fa2b0e761bf641629b61aa0508575039d5ce2efefb7dbb1d7b25da2b3553cb = I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847 + ~I06414f803df7c8e59f01524020e09627cb11f3809c3456a9a64655062b110885 + 1;
            I7e43798e3391bdb6c6a9a6ad85e51c960fe4bba982ae765cecfb287b0573e5ff = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I73fa2b0e761bf641629b61aa0508575039d5ce2efefb7dbb1d7b25da2b3553cb);
            Iac70da997560fcd3949fde686e6f8a3dc834a2ab7ff2beaeedf7614710bbfaff    = I7e43798e3391bdb6c6a9a6ad85e51c960fe4bba982ae765cecfb287b0573e5ff;

            I513c50e5893017204f1fd591753a0f5d29f4b4ffa8466c613a9d12d419ca8281 = I2416f8532fa923a4979b7153c048e71fb582124c5a9147bdade98438756f3847 + ~Ieef9e0d39f2e213f365af4a6a34d0d2c7d50155e8052e9b1944473641922e9eb + 1;
            If8b3199a20ef98c9f204d2a8686fa71d5094b2e701c6f84b7630ddcce89c77c2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I513c50e5893017204f1fd591753a0f5d29f4b4ffa8466c613a9d12d419ca8281);
            Ie32e4f67efcbea2f033a66104b3315b46a1c857781ac63283f4d955384bcdd4f    = If8b3199a20ef98c9f204d2a8686fa71d5094b2e701c6f84b7630ddcce89c77c2;

            Ib2deb611e086f8f21f132eae3b128b0b8dfa06caeab1cf2fe25f94801fc4e184 = Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1 + ~Icf9f5e717c65afd1b3bbc3d6c1bd960155773ec7790543f56c86637a891decd9 + 1;
            I916b56be359d608276fb2fe1be1c65df20d635e00211fdba107a1d6f9c0f0a36 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib2deb611e086f8f21f132eae3b128b0b8dfa06caeab1cf2fe25f94801fc4e184);
            I4720d84525310ad5428da40677f1cd99365d1467c29d214ab4ae300277322cbe    = I916b56be359d608276fb2fe1be1c65df20d635e00211fdba107a1d6f9c0f0a36;

            I427ad9ada9b609bf66d313618975a2a4702011b7ef9e55e40d37db31cf075173 = Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1 + ~I53a66c670d7345059cea712c026fe8c524e74b030af0de054cf6e053bb304248 + 1;
            Id0b3cca386cb4a6627354dc8fcb01c27aebb58435b78d7df234937d5aa2bc457 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I427ad9ada9b609bf66d313618975a2a4702011b7ef9e55e40d37db31cf075173);
            Ia1f10017528e76925426be916c558186f2196a0c4d7520e57e0895e14e7c1d53    = Id0b3cca386cb4a6627354dc8fcb01c27aebb58435b78d7df234937d5aa2bc457;

            I54c2c2be59b9e302a4527e1fe4136fa3c31561d04ac55f71fdc5bbf8b8488e39 = Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1 + ~I0734166e34887037bf713bdf1df0f7219241551cec455ed45881734727f90032 + 1;
            I72ad7a4f024406e89bfc87296a9c0456459b729b9e4adb046d703069cc9ed1fe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I54c2c2be59b9e302a4527e1fe4136fa3c31561d04ac55f71fdc5bbf8b8488e39);
            I46a3710c0e472a92b83354b668ac21c775b2c4e3dceadc49dc0cb712c08c319e    = I72ad7a4f024406e89bfc87296a9c0456459b729b9e4adb046d703069cc9ed1fe;

            I40cd513b6eb8a99d78aecb88ba332afcdd021ecdb00ee89d894853f642077211 = Ib289bf22265ed1f0e61f49515b4515bef7ac1e3a2af662c7720ceea89157cfd1 + ~I4771e59053fbd3e261c49e0be7e742e7cf9c5bdad030b67f1b955e13e9bcf083 + 1;
            I725f7893c803b548e668b87cdd368f2b26e58193cca109b618d87e949b8b0d25 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I40cd513b6eb8a99d78aecb88ba332afcdd021ecdb00ee89d894853f642077211);
            I594b73c43f22c1cc15daf1eb602be4366502100a0ad3a3bad7b7992c9839dbbb    = I725f7893c803b548e668b87cdd368f2b26e58193cca109b618d87e949b8b0d25;

            I2de25ddd85167a3af17c87c103f1d19ce367d6e020475b5440aadb42896091ac = I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333 + ~Ibf4bbd894f269bd6e6eaf9511141b91ac61b5dd3e77b4ffd07aa88474f251ddc + 1;
            I5d49190282814ee6220a4a003e2f4879a2e37459fb2c3a1e1ffecc35f57c26ac = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2de25ddd85167a3af17c87c103f1d19ce367d6e020475b5440aadb42896091ac);
            Id6264ccfced253e14f1f9be10f967d475695838c367808b97abbd7578447179a    = I5d49190282814ee6220a4a003e2f4879a2e37459fb2c3a1e1ffecc35f57c26ac;

            Icdeb4cc4b7cfd480c2fbeabb3f8e1ca72b7af731726a0ecde4c097dcf4d8f6a0 = I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333 + ~I7c10e2245efc27a4e2a96467eb4e3fd9c28be5f26f65c560653ff4742fa5143a + 1;
            Iebcafdf2cd96dc5a859f7087ad96383f07d57818696f1522555720021c3fa8c3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icdeb4cc4b7cfd480c2fbeabb3f8e1ca72b7af731726a0ecde4c097dcf4d8f6a0);
            Ied0e2037bbb2f2b7d0cef3d7d3f5b7123c006255cb7f2297df7e1a1eb03dee16    = Iebcafdf2cd96dc5a859f7087ad96383f07d57818696f1522555720021c3fa8c3;

            Ib6dc79711e470184d6cc3f360fbefc3c55c32f612d1743111dd6ca9b96c1a4e8 = I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333 + ~Ia7a158b91a24000cb6211d129d65e781a4e28b8333f897bb401042fbe17c37a1 + 1;
            Id8b5082d5099ba65d612d86118ba3489888d375a6d8dc1816ca6c4338150b98d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib6dc79711e470184d6cc3f360fbefc3c55c32f612d1743111dd6ca9b96c1a4e8);
            Ica6a39f57caae5761078aaf00587554f1acef5d9b2e1fb73931f5715ebc762dc    = Id8b5082d5099ba65d612d86118ba3489888d375a6d8dc1816ca6c4338150b98d;

            I2be6b0805c51599f698f3997780a6f81119106f870a679c00221c9d173040d5b = I754b572c6ce9d598bc275418d690728bf7b2020eda37f2829e8686a507e1d333 + ~Ic8c13812ba09457021ec6f39406b1106dc025551c62da4259930c361f19c3a2d + 1;
            Ia11ca5043541c5c51fba4205915afd0b4e97bc70d10317e9d3b952138dd15572 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2be6b0805c51599f698f3997780a6f81119106f870a679c00221c9d173040d5b);
            I0fe26cc77a5b117d82b8f0da27f4cc5e9465360eba32d35aeefc16ff600ad5f2    = Ia11ca5043541c5c51fba4205915afd0b4e97bc70d10317e9d3b952138dd15572;

            I09831b2bce6477d49a664abacd23b6be52c85544ebd549b0943f4218cc955bed = Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0 + ~Iba1a21e329197ff5e399aca440cec6d6bd3d9593c332cfcba84d52d541ff1ae0 + 1;
            Iefe655d513457dbbd05f22922accc5bebfc22843447254ee0d6eb4b48056884b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I09831b2bce6477d49a664abacd23b6be52c85544ebd549b0943f4218cc955bed);
            I8bfbee6346d016ff8cd0ef681e0efdf28d0f27b3e887397fa1aff647739e25a1    = Iefe655d513457dbbd05f22922accc5bebfc22843447254ee0d6eb4b48056884b;

            Ida6c7b0feb190489db3cdcd850ee5d64baa24ad7fc56b615ac1103f3c5311e06 = Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0 + ~I3c91639fa462a2a7e65410080b46408b692ca4639ed17637b1d465f38631734d + 1;
            I5e23dd0658534242ac135a6b401ee146d0ba48841d3464a8c58def92970d50aa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ida6c7b0feb190489db3cdcd850ee5d64baa24ad7fc56b615ac1103f3c5311e06);
            I57f07e2955da5218122f614720d5890af9d7b5ac4f033e9d1c10db08e7ad1882    = I5e23dd0658534242ac135a6b401ee146d0ba48841d3464a8c58def92970d50aa;

            I56189306e5774d3a224a89042fa23eaf4af107e2fd4fb1f6261943a46f8d8bfa = Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0 + ~Iee901b35683b34719c33d63d90b8ae11fbc338a170164aac943fb0b495c92b97 + 1;
            I4190e8ea4ed62c9f3512e102be78d80de31e05fdb31f39bbecec25c5fe4838c0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I56189306e5774d3a224a89042fa23eaf4af107e2fd4fb1f6261943a46f8d8bfa);
            I9c71f3f968f3265215ce730a5f922db81aa408218fc76de3b64ee4f9396d3f78    = I4190e8ea4ed62c9f3512e102be78d80de31e05fdb31f39bbecec25c5fe4838c0;

            Ife7eb04d87c4840ec5a25b0b50ac641fa8ae6ff206065248ad8ac718cbfe5272 = Ie59df8d18b771b60ec5922abe5bea2eccb547dc890fcd10f5cc444397b8e39d0 + ~Ic7aae8edebf83f3971440fd0e86e7700ac4cc0c087c9996d55cfecea8c489fa5 + 1;
            I22800d7bf254d48f28f9d0e56af31271b20bd989575a3ae510dc64f592b1e08a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ife7eb04d87c4840ec5a25b0b50ac641fa8ae6ff206065248ad8ac718cbfe5272);
            I3afdbbfca5c952e1800c1e15ca629173eac62810b6bf8097421addeae979ca81    = I22800d7bf254d48f28f9d0e56af31271b20bd989575a3ae510dc64f592b1e08a;

            I2ecbe2abd1b3ec06de80c5ba7b5f1ea7bc9484559a134199749c0eaefbc1f3c7 = I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114 + ~Ib5a93c88521f26a686316f032821a4e9540fdd8e93570ff35437df7522d34ab7 + 1;
            I4bfc7db23a7b268d945c751ac989718287b1730e8ec35d623ea7636b6946d554 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2ecbe2abd1b3ec06de80c5ba7b5f1ea7bc9484559a134199749c0eaefbc1f3c7);
            Ie9d906bda89623d793bc65968cd86bd0c63458c7a6b12fd38f7054069dfcd132    = I4bfc7db23a7b268d945c751ac989718287b1730e8ec35d623ea7636b6946d554;

            I1120c79480e003c87e8160381c89f4a6baddfc6927ae56952a233f96662a8a47 = I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114 + ~I0806d1e2ea1771b325ea80b71fe9223f495a3831a560f579401b4e94b6ed172a + 1;
            If4a3f6ad253dd104911b6d1a09ae4a3ece88afedd537e8f7fdfa8735aac88fc2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1120c79480e003c87e8160381c89f4a6baddfc6927ae56952a233f96662a8a47);
            I969b9fa05c651f6e2f2dc426e35c43864f9b5c6d4f6278b0f7ec4e7c5e872eec    = If4a3f6ad253dd104911b6d1a09ae4a3ece88afedd537e8f7fdfa8735aac88fc2;

            If0294554b2637dc70b079fff36543d68234f3f8e9d80ed67466ad3d8ab4e5f91 = I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114 + ~I7f1329fd762cf679c07aced91992aea071fe128bc24f06ce88bf49e876578a9c + 1;
            I2ec9f763c06f61ba0e1a2669b6ee19aa5be8a80a6ce04c0355956dabdad55e9b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If0294554b2637dc70b079fff36543d68234f3f8e9d80ed67466ad3d8ab4e5f91);
            I436c98ccee6d1a138f1c47ef4e5b7ac39db15122b2b134828b257dd629e310a5    = I2ec9f763c06f61ba0e1a2669b6ee19aa5be8a80a6ce04c0355956dabdad55e9b;

            I4c82e07db2a69392d528b47296fc3ce9bd342a9ddd3720f059ec38ea10b98efd = I2a6c4099aae304c169257f111ff3e350491908b5a8034d7a062f5869c3b86114 + ~I091bf548253a3b22f92aca6479b70ccb74a5f9eda8bd80e6bc1e059021f04b9f + 1;
            I280472596040e145f7bf9d23aac7c569dea951975e67e53b2677fca092dc4fa6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4c82e07db2a69392d528b47296fc3ce9bd342a9ddd3720f059ec38ea10b98efd);
            Ide4ad5678bce6a696f0c6cb163eaf670c47c2506acf7977c1031c6ec03e03a58    = I280472596040e145f7bf9d23aac7c569dea951975e67e53b2677fca092dc4fa6;

            I03b3c7c34463d46735abd1392e5bd16a783f79adc25f3471eaede71318ac5799 = I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a + ~I13f5f01dccbdf3df23c5bf603a9657e161c1e2368cb5cb48b212231d2fba7794 + 1;
            I593137c88d2dc13a0bf028b949e6ec556b7787557f6a5c72f0d1161db6b096fd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I03b3c7c34463d46735abd1392e5bd16a783f79adc25f3471eaede71318ac5799);
            I043258a364cd91821e9bb3e9c46441ac7d330c706e4b0b7e29c4b92f7c5ce562    = I593137c88d2dc13a0bf028b949e6ec556b7787557f6a5c72f0d1161db6b096fd;

            I8cf7dd68cf30611d1b03b4205f1a8dae3c8f8f943c04773e335a2ea90c555b3c = I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a + ~I840289556d82218416d7f8652d40586181f7b4ecedd132450594aac1bc47a081 + 1;
            I331fc2f98c551ea5b177eb3f3c1072371f7f7a02e45d4ae3fb41bdb96cf7426d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8cf7dd68cf30611d1b03b4205f1a8dae3c8f8f943c04773e335a2ea90c555b3c);
            I2f639b76b1afd86d9ba4d07d54f5b45df8cb99d7bc58cafd0c1a9a9001842260    = I331fc2f98c551ea5b177eb3f3c1072371f7f7a02e45d4ae3fb41bdb96cf7426d;

            Ic8dc799519d1df013b35ee5ba849490330504471458ece8164705be772acf907 = I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a + ~Iaf763109fb82e88c7ec019f7b9b668f88f84a5d4f760592d2dc9172c75be0aab + 1;
            Ic5a2e5d00e362ead90ecd9182e61b0e3a99a7756994cd358bfdecf8ffd957491 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic8dc799519d1df013b35ee5ba849490330504471458ece8164705be772acf907);
            I1dd0421d7e31a316541c339f8b4f1e3afbe37ce09254ed825c1b6086a0c0f3f2    = Ic5a2e5d00e362ead90ecd9182e61b0e3a99a7756994cd358bfdecf8ffd957491;

            Ib44073e6dac33e4dc0f497a79d4bdba9dfa398c9e95af1cd3c5406449505fcca = I0f9fe6d4d83a911056f4d0ccf7320ba3df1732cc3c956502d41636f17f0e834a + ~I5c1c30033bd61b271c765ba00b033a58c6389d4bd353ce68d1b193bc7138baf4 + 1;
            I15f2b29740b5d1a9a5412db4a0bf09bacbde963b08c243ebfbb4740dac56349f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib44073e6dac33e4dc0f497a79d4bdba9dfa398c9e95af1cd3c5406449505fcca);
            I50ccddac87e61ba10dd9410a224c74ca88b521dfed962bf601c38ae78299384f    = I15f2b29740b5d1a9a5412db4a0bf09bacbde963b08c243ebfbb4740dac56349f;

            I59b6dcd7306c00a99dad76ca16c9dd989f5dc46e7358a8c0943fae147da7b884 = I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210 + ~Ife767fdd58724398b336a58803ca328013f3a8228ede0cf108dcae054001de56 + 1;
            Iab45b41ab7c1056072ef64483afe800af63354919bd1a7ec95cd3d9219ab0301 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I59b6dcd7306c00a99dad76ca16c9dd989f5dc46e7358a8c0943fae147da7b884);
            I5fd9960aaa562ff70e5d0e913dd4d88aac1b73a95c41ba903c0b7fc4dd4d93b2    = Iab45b41ab7c1056072ef64483afe800af63354919bd1a7ec95cd3d9219ab0301;

            I385d65a11a7e793cb8b1cd9df81bb73d8ce3075e9eeb389c6b9665be6f3c5ce6 = I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210 + ~I58cee4a472b2fa2f17266cd6ab55d475f304bbee835aac31ac7879d77b8a23eb + 1;
            I96c8864be45f3a0501bcfbccd5bc984738c1e05cf6834d8aad47468465908abf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I385d65a11a7e793cb8b1cd9df81bb73d8ce3075e9eeb389c6b9665be6f3c5ce6);
            Icdff2336860758127c20c1d45d5723511fa42577417bf4f77d0c770abcbb175b    = I96c8864be45f3a0501bcfbccd5bc984738c1e05cf6834d8aad47468465908abf;

            I1ef957fc8b1559a10bf1f189ca736164c0e50b50786e31c70168fd2e0f65aaca = I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210 + ~I3724769b2a595469f910cfcf1f002009d9fc27808df7e59ce728af9a923726d5 + 1;
            Ic01034eb6c2ef07602777d1a6ce7195524d4d1e3093d15966e36f45fd58d5bb6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1ef957fc8b1559a10bf1f189ca736164c0e50b50786e31c70168fd2e0f65aaca);
            I9351e784be3825e94dcf67151cf38c9fddcf244bf5512db57dcc612882b449ce    = Ic01034eb6c2ef07602777d1a6ce7195524d4d1e3093d15966e36f45fd58d5bb6;

            I2ce557a4098587fafd3adf55d2195fa2b5c7da844d59ee5c4fd14d11374b58be = I02b15d57d48c99d9790f241e0a23b1ebe0e1510a842ee980a9ca3576fd7d8210 + ~Ia4370635785f2b904fb6ab3b8cdb86fba5445230a9d3d02cd908e04d92726f3c + 1;
            Iaabcf58807b565d00812cdda849cdc45a34b1e0019a539ddfcc9aa957814de19 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2ce557a4098587fafd3adf55d2195fa2b5c7da844d59ee5c4fd14d11374b58be);
            I23f7465a60acd0fb198e753834d30932ddab8939bb2df2172f54c7bdbe02e154    = Iaabcf58807b565d00812cdda849cdc45a34b1e0019a539ddfcc9aa957814de19;

            I384bff3d8617787aa577ea8607bf3f4ce49eb412b603810e854e8ee59ef3114f = If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48 + ~I26ad8ce808bb26201de4f63afd861583af9abc55c7623bf15bd1808c0b0c2be4 + 1;
            I5cac542afddc74aa26163f65fddc7689b04bc5f3bf1fda74a7557cb4dea506d6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I384bff3d8617787aa577ea8607bf3f4ce49eb412b603810e854e8ee59ef3114f);
            I40687a0e9fee803f38df7cf7dbc3d3107b859b4e80822bc59a157fdc606416b6    = I5cac542afddc74aa26163f65fddc7689b04bc5f3bf1fda74a7557cb4dea506d6;

            Ibcc6e1c0808d4a22bd66ca467b66a5d5fb1d60d5faef295c6abe67319e782ed5 = If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48 + ~I5246ce1dc41e20a5e4e3312a997e8c5be2d733f0cc95f74caa7e668f9ad2f1d6 + 1;
            I3fd692bcb65a1508f7a095a74ff2159e97a3c5c14ddd8b2c96a7a2bfe43d07e0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibcc6e1c0808d4a22bd66ca467b66a5d5fb1d60d5faef295c6abe67319e782ed5);
            I807d8cd303e5c8c8379a9a2954804c606d897fc06412c924a89f3dc9e29909bd    = I3fd692bcb65a1508f7a095a74ff2159e97a3c5c14ddd8b2c96a7a2bfe43d07e0;

            I26faf05df42ea98f85655adde1199ac6e46b738ff8a2e0b218e2457bac1fc3ea = If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48 + ~I1de9fe186e9fdadc6c62a9c6645dccfd3709778f3243d2a4155bdfa20d27a544 + 1;
            I0fdc11587841ff68e0606d5e9924388a5822c1f6f5c3dc2ef406e3af7ccf4e4c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I26faf05df42ea98f85655adde1199ac6e46b738ff8a2e0b218e2457bac1fc3ea);
            I1244d935c6db7b5441533aab87f518ea215aa6f5903b071f2ee8cb3359b3bcb2    = I0fdc11587841ff68e0606d5e9924388a5822c1f6f5c3dc2ef406e3af7ccf4e4c;

            Id337fd09c4d42ecaedff4e08ddd14fa65c5646caa08bd75d6c274bb9a48033a5 = If5df64d3ae3a434a9e58c75dcfa1c9cc827d428341fe8b1c781d0f36eb814c48 + ~Ie73ab4d16ef614a27522cdfd47f670a38ab58f89bc10c74975cf0b30400e198f + 1;
            I3245926b69b2db031c68574a86f56671d4dac371989b6670fd5cbf1106c85606 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id337fd09c4d42ecaedff4e08ddd14fa65c5646caa08bd75d6c274bb9a48033a5);
            Ia7cdab2a88c99d9780bb267234b2cb87946009484d21f4419c50e7570438e645    = I3245926b69b2db031c68574a86f56671d4dac371989b6670fd5cbf1106c85606;

            Ieb6923956eb85d8a6c65882d8673b841dad39fe763732488f568784d7f5d746d = I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab + ~Ic4e32c1234be0a530c66106794dc1114e4c88611be106ffde42a7ae486560ae5 + 1;
            If7e27c6552a8a17a2f1f9fa61cc6b4c478f1030f1ca44dcb98424d65cbf10f93 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ieb6923956eb85d8a6c65882d8673b841dad39fe763732488f568784d7f5d746d);
            Iacdbe6e2ae2cd5fa475cde0217452a14f05bc8d499b9ddeca568f6cd96ad6a2e    = If7e27c6552a8a17a2f1f9fa61cc6b4c478f1030f1ca44dcb98424d65cbf10f93;

            Ic1c0ecc66995dc98197e5e73789f8f644f15547d4b130262c526c636458d3712 = I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab + ~I42ba6c66d951bbe03a57fa7a4926d6323f30784fe87de73cce065cccaa9814b1 + 1;
            I37d8e18c384970e7a81bebcf85fe71c569fcc09b47de629e2258eee1c837ff31 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic1c0ecc66995dc98197e5e73789f8f644f15547d4b130262c526c636458d3712);
            I5aaf6ccf4cefc2732732ddd816c3eb7aea7146c6e7abf913a5193f6906fe9497    = I37d8e18c384970e7a81bebcf85fe71c569fcc09b47de629e2258eee1c837ff31;

            Iee6b04715421c83b0bd430ac4891dcf8a2df5f3fd80478d80de33d83f31d4fa5 = I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab + ~I735ec7a402f471520335d15ee3415e874f56381a2c0cab5c3a5b21f7d6f71474 + 1;
            I8d5e26d702af2d2b53b135bac7ec7097af7f878392c518c52571ead31ec485ce = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iee6b04715421c83b0bd430ac4891dcf8a2df5f3fd80478d80de33d83f31d4fa5);
            I96d8c1b67b028322f3d3e46d6306eac0333a8f3fe45073c08c5267157f73b71e    = I8d5e26d702af2d2b53b135bac7ec7097af7f878392c518c52571ead31ec485ce;

            I6751fa1b7cb41d853b4affcbfbda7f7f959e4a7e4caad11f988e00eec5acbcb2 = I8e7e3fb7bd9b4d93b72b9305ff8445d4a5f03cfe0bc0b440845696733ea7dbab + ~I76b8cfe5d3985f3c0f249680ed81aa3b21cd7af725925846e8875ef9e98a550e + 1;
            I1d7ba7c6a56849ae78cfb42345e7510951e81fc92ea2aeb04addc6d3962e2873 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6751fa1b7cb41d853b4affcbfbda7f7f959e4a7e4caad11f988e00eec5acbcb2);
            I600b1d1ff12460bfbaf32de67aff0e32087306628f0ba7db6736a81354309a41    = I1d7ba7c6a56849ae78cfb42345e7510951e81fc92ea2aeb04addc6d3962e2873;

            Ic3c16686cf48a3d8cd9abf2ee2c917a5dd071e8573454b02340f6e847302b029 = I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea + ~I668775bd016b2384bb3d1cb0a1e89a76d2af15b2307cc6a5d2e0d6c699b02544 + 1;
            Ib8248e176e10a6ee79f77bbd56fb4f86d032c600522b20afc7fca399010fdfee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic3c16686cf48a3d8cd9abf2ee2c917a5dd071e8573454b02340f6e847302b029);
            I225db641808b767d3f529e5ef2ac066e3abe953b8b434fd7bf4e02b57edc0f27    = Ib8248e176e10a6ee79f77bbd56fb4f86d032c600522b20afc7fca399010fdfee;

            I62722b1482f18c3ab03a94e845406bc30c1c47102fadc9b9642096ff3c504cf3 = I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea + ~Ic8108e830a58b12b8e3ef4897cee70758d1539ae6609d73b5455b94b0eee5510 + 1;
            Ic35e7904ec654dd5f5e382f1df5d76cd1e4cd0af95a57ed979a5b369ed8ebdb1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I62722b1482f18c3ab03a94e845406bc30c1c47102fadc9b9642096ff3c504cf3);
            I1b7380bca98b56ba1a2c2ad5d78fdadc1112b208e8d98b84c8d950f3f12f1658    = Ic35e7904ec654dd5f5e382f1df5d76cd1e4cd0af95a57ed979a5b369ed8ebdb1;

            I968319c4ca969a6396cc16b20098933dd8669213ba401ebefcc50670c0fac5e4 = I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea + ~Ic5921b5017385aa779a2016014d381a982c32c64d1643e79631a8ac842d5b584 + 1;
            I412c9dbea5975fe4fd5089a5d5b7e4270992142b7c2a5c4b59f2f6637215558d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I968319c4ca969a6396cc16b20098933dd8669213ba401ebefcc50670c0fac5e4);
            I651492ce35fed9d77d5167dd211125ace0af8d55b8aff148e760d8919d53b6b8    = I412c9dbea5975fe4fd5089a5d5b7e4270992142b7c2a5c4b59f2f6637215558d;

            Ibff476e387614c2089d64e400f457e70e4c8ff251bdaeb48e85c68f1756dadaa = I11265ee7f2bf2d1acf382814494fd0f2d19a317ed3941c1a9b792dcdee1bafea + ~I58919d58783467b7ad0108f86d6260f3c551692d00e6639260a68a7a512d8689 + 1;
            I480a5bbf4a2b6087f900087a2dc6c595ae36127a85d6551a9586443ca5c793c0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibff476e387614c2089d64e400f457e70e4c8ff251bdaeb48e85c68f1756dadaa);
            Id732b4b9de3f715537d32d6eb6eca4f6f9fa6d634bc283ceaef531bdef605537    = I480a5bbf4a2b6087f900087a2dc6c595ae36127a85d6551a9586443ca5c793c0;

            I16a9ad58728f11ad740c8517c5b084638388bf79ef9e4b8e845eccfa31479069 = I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4 + ~I9075819cc111daeabcc2ddedb4a4297b1a42ceac8b93213f7f76d0fe87c8c275 + 1;
            I2d42f8280d91ee6fed549f956ed81dcb31e70acdd0fb1fe4f63aa2bd3a7878f4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I16a9ad58728f11ad740c8517c5b084638388bf79ef9e4b8e845eccfa31479069);
            I78c5859a565a68329d5f75effa2fbe77e16d86bbfcaf79d5480374f8bb87039c    = I2d42f8280d91ee6fed549f956ed81dcb31e70acdd0fb1fe4f63aa2bd3a7878f4;

            Ie73acb967f41ab47a4828279172548c8a36b7b67a4129138f12f9715172047aa = I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4 + ~Ia187792bad45afcf25df25b18a076d255536e94db8d7bac4df79761df5f16050 + 1;
            Ia29c45f92e3672c1b0c186b711e5f0eba39186fccd95905a2bf9791609b8bccf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie73acb967f41ab47a4828279172548c8a36b7b67a4129138f12f9715172047aa);
            I411faecc88c5a9fcbc433d784eccf7024675c9b009564295eeb765079b8069c8    = Ia29c45f92e3672c1b0c186b711e5f0eba39186fccd95905a2bf9791609b8bccf;

            I769e3a9e63f6b86940c9136476d851dd2e123b17d42191d5fa078828c2ebbb6e = I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4 + ~I424c57a79fc220d56d1e499af6318dd2a2f4a4ebab1c83cc7762658b8c34479e + 1;
            I9572b18d2f9aa917168f389e7066eb543c9036fb55680d5dfda1e70b4d7a1193 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I769e3a9e63f6b86940c9136476d851dd2e123b17d42191d5fa078828c2ebbb6e);
            Ic429f74c6e97fa699700391c81e8a8ac449270476ebded49a8bcf8161a19260e    = I9572b18d2f9aa917168f389e7066eb543c9036fb55680d5dfda1e70b4d7a1193;

            Id8b5e6165cee66382652189754f7afb582423212885be9cda93c154f46942297 = I30e6985f1469cc76ab28cbce5065ff0545ab09e36ca173637030ff99306778c4 + ~I0d276f9604ec2b8621a86706ad1772058a29e94902e8eece60e3d07948e24cee + 1;
            I447026649273854452afc7335d4d52926fffb5950ed7a209f9f31e5aa95d6336 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id8b5e6165cee66382652189754f7afb582423212885be9cda93c154f46942297);
            I6efa3ca79fc64053e7e2744a4248a5c0df63ef15c66542967b53b2fcefe0d286    = I447026649273854452afc7335d4d52926fffb5950ed7a209f9f31e5aa95d6336;

            I104e372ee724bc6151a4854bcf5896bd1c49ff41214b0a48b3ab13f1b06d3fe3 = I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2 + ~I98ee0d4994c76a87aaef2967ab6cb88af05ab0a7972d2dedbf115ec19c426fa0 + 1;
            Icb1f8fa764a70745aecd528189909af5082393c7f4d69462d6c069a011df5c6a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I104e372ee724bc6151a4854bcf5896bd1c49ff41214b0a48b3ab13f1b06d3fe3);
            I00827962c46c637f5d74d450ff4eae848b4cb15add5bf1f607708b76c8551c21    = Icb1f8fa764a70745aecd528189909af5082393c7f4d69462d6c069a011df5c6a;

            Ia841ffbb8205a284e28cfd445b7b459f11034a0244d777b7136fe0a6009b53bc = I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2 + ~Id5eaf1d953b17df3896f9a30f37363d1a69fe3a956b97d307c895065ff32674e + 1;
            If7730750ecb044040333f33232026110e55becb8df689868897b76fb093b5bc8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia841ffbb8205a284e28cfd445b7b459f11034a0244d777b7136fe0a6009b53bc);
            I6cb1364420f9bdd072770a684de242f89990e3f144f160c2f5311bb00fe4daa0    = If7730750ecb044040333f33232026110e55becb8df689868897b76fb093b5bc8;

            Ia4613fe4f54fd9c2b61f4524bbc42c67307f872c50b5af9e9a836e9cbf8adf22 = I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2 + ~Ib5e2defed9b5fe67a6a551e253cf68006aca5e13092f7e9b53f8186c76a156dc + 1;
            Ie2ed41aedb52e82863b3dfd580f2d2b7aff367f1613d274ddd5a5114316f858a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia4613fe4f54fd9c2b61f4524bbc42c67307f872c50b5af9e9a836e9cbf8adf22);
            I41bc9fc093e9f311e6376edb8aa0640709fb3bd420ff8a7cb2092844fbe0e121    = Ie2ed41aedb52e82863b3dfd580f2d2b7aff367f1613d274ddd5a5114316f858a;

            Ic6c4976cc23f404b5b1d328f991e6ff7385f3bb0d61392626bfa621147866147 = I1c9ff360246e7966a599a29c14c8967751b529c3001a3d478594195ec41920c2 + ~I5463c05b1b55c142012470d627accadd8e34924e77ef6d139b3fbe1db1cb91e8 + 1;
            Idb92f51d1c0528dfafe1997ed4a9539f2f3d1b02900558ba6828e873a098789b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic6c4976cc23f404b5b1d328f991e6ff7385f3bb0d61392626bfa621147866147);
            I84519b5d45c05d737fb27ebd20ddbddfdaf7a22125df9eea17400856eed27992    = Idb92f51d1c0528dfafe1997ed4a9539f2f3d1b02900558ba6828e873a098789b;

            I59b0c136216dcc5613e45a5a841bde1c8243d06cea7caaeaabe614e968228d6a = Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597 + ~I7c6ea337917ea8eb0696c514db7ffb66719763162bdd0b7e0ac764c1ae63d24b + 1;
            I21742c373c52ea0c4872995841566c199318bf1f5849f05df796b79e171934b2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I59b0c136216dcc5613e45a5a841bde1c8243d06cea7caaeaabe614e968228d6a);
            I3af2de27ab7a899c5e55f150a53b7ef65e88309f4280269afb3eda2b1b408d05    = I21742c373c52ea0c4872995841566c199318bf1f5849f05df796b79e171934b2;

            I345aa1fe14f36a465f2bcb4de639be9f617e5d22257cf97f8eb35096383a8674 = Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597 + ~If2cfdc638b3cfc13d31615533cea59a4bf8123299239956479d3f1d702ef54d7 + 1;
            I541077747787cf13e4c324b089049dcda6ff46c252b180e3d2c8f5b422217533 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I345aa1fe14f36a465f2bcb4de639be9f617e5d22257cf97f8eb35096383a8674);
            I988d8e969e2a2ecac68a36a5f4eb0d6cb2c325e4be24c4716625070057ab9538    = I541077747787cf13e4c324b089049dcda6ff46c252b180e3d2c8f5b422217533;

            I1bea08777eb6009228b55fb534f502ea7deedeb705d33d4e56a7b5107a9a11e2 = Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597 + ~Iccb7ca5c2ab8a9a4e3776ef42997d1d645c5542c25ed35b161702ce450f90fd7 + 1;
            I1fa1de74e664f3ed0ac923d6bf1a11fd74a6337f2c8f983d8b3dfe0f6737dc4f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1bea08777eb6009228b55fb534f502ea7deedeb705d33d4e56a7b5107a9a11e2);
            I63ec7fce46bb02bd1662b19d58025abb479c4b57a0e4fd0642404ddf7f607077    = I1fa1de74e664f3ed0ac923d6bf1a11fd74a6337f2c8f983d8b3dfe0f6737dc4f;

            I5d6f4230452aaeb0bd33f7b39b467450b11175685cde0958391f4e7f5ce44847 = Ib31566c11aef2265f4b7161955923b1f9b6493671011842d39b2791d9835d597 + ~Ifca2987d8c7f1ca30013ddfcdb82a888ebbd7bc3dc421f7e3d6806f5f3a9aa2d + 1;
            I3846e68c708bbe037e97544fc1cd70e7ed94539ddcad0d21984791ad35556d88 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5d6f4230452aaeb0bd33f7b39b467450b11175685cde0958391f4e7f5ce44847);
            I086c1b2b7346139212d810647d98824eff245a9e24fa84006583fd56f1e76926    = I3846e68c708bbe037e97544fc1cd70e7ed94539ddcad0d21984791ad35556d88;

            I328d56833be24a38552b6110e2858dbbc3561a3783d9255efb5580d9f4071749 = I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0 + ~Ic55bde9a87033c380a5cfe5736d205c15099a2f2cf440f88472d7f6e65d360e1 + 1;
            I2b00e353fb14caee3c8e659e4c76b55ddaa6a17394c90f3fa53e52486059030c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I328d56833be24a38552b6110e2858dbbc3561a3783d9255efb5580d9f4071749);
            I401154446147692cdd273c1d6dbe5a225e466799d41dd00f9477c586add460a4    = I2b00e353fb14caee3c8e659e4c76b55ddaa6a17394c90f3fa53e52486059030c;

            Id835c902546b418343c3e52de8260db4304844475cbc1532389305577624e4cb = I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0 + ~Iaf14e804e3bb7cda8e67e39af906be2c966fbab4a6e73b8d60ee7ac5733669e4 + 1;
            Ifc3f186e24f214ba2d389536a913299116a402cb32c161f67fc854d73396e087 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id835c902546b418343c3e52de8260db4304844475cbc1532389305577624e4cb);
            If832820141ab4f3c34efb429966b47ce584cf58fd34d38a7ecd976235613c541    = Ifc3f186e24f214ba2d389536a913299116a402cb32c161f67fc854d73396e087;

            I8e604b3839cbca0e894ecdbb66a3c24f49a91c523f29e8984fff3e8bd1bb421c = I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0 + ~I5460bdaa1d2a7c1cb2e75baa2c211593afac76ce5160a620b385393217b4185a + 1;
            Ia86976aba4570aa0ae88d5ec887ea058cb4f7b49d7ec46b0ca215162564b1598 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8e604b3839cbca0e894ecdbb66a3c24f49a91c523f29e8984fff3e8bd1bb421c);
            If13409b9d8c65fe2127031b0e4f953f55c8a66c06811c6a5d261372aa2986511    = Ia86976aba4570aa0ae88d5ec887ea058cb4f7b49d7ec46b0ca215162564b1598;

            I402b028195ed3aa64305d0cbc85fa79e1f172c79704f8fbd86b74770352a2908 = I3f016cc0e914506de126e31ae0f59a066be52bc819007ee9707bbb55b79aeba0 + ~I5ff269ab544d2b74059a73d0ffe0492473b214d392d8c2ee760847e6c07a361a + 1;
            I5f93ff96a38e7ef38f5fe0f41333327e06adb0efc0ccc4c442058b75966ab5a5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I402b028195ed3aa64305d0cbc85fa79e1f172c79704f8fbd86b74770352a2908);
            Id2bc1d218fffb230a1505feb20cfb5229db9f3e2b0c7bb005bc8c59403fa35ad    = I5f93ff96a38e7ef38f5fe0f41333327e06adb0efc0ccc4c442058b75966ab5a5;

            I56ee0a1de27160410a2bc12cd4d550a3fcd4d560d81348cc36e94746f46f6341 = Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7 + ~Icbbddd7f07e1deff7aacc0e96a33556b62ba127dce877dea351b421ac8d00313 + 1;
            I9a2901c60b8a175d5462c32e4922a0bd931a186384b519b751929e551b477efb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I56ee0a1de27160410a2bc12cd4d550a3fcd4d560d81348cc36e94746f46f6341);
            Ia1846f3088723131b0fc158b2d942749466887bf940e29340846070ac9d5090b    = I9a2901c60b8a175d5462c32e4922a0bd931a186384b519b751929e551b477efb;

            I0c0d3684d621cac560ca9866f49e30d1f66c34c35b2e1112f078ddd15b79d826 = Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7 + ~Ica809c2eeaf6926552d9f811bf16c30146853674185c2315876fb5b2ea6d0769 + 1;
            Ifa5a98aa90cec881eabe5a6eee07f971778a40613c80891ff994d5a32d9ca6dc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0c0d3684d621cac560ca9866f49e30d1f66c34c35b2e1112f078ddd15b79d826);
            I5d5edfd68cef65681c36f4bcd770ec84a721eb515bc1d0fb7603ee0f5a63fabb    = Ifa5a98aa90cec881eabe5a6eee07f971778a40613c80891ff994d5a32d9ca6dc;

            I6f62f4f2fc06f1cb30147da56b8fc88874f748262e4308b0d794c057267d9ac1 = Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7 + ~I0583863d43273e6464e5e65a8714be627f867a0320302382d94ef661b21f73d0 + 1;
            If367e1e075614957d2fd83c76b45a3ebe11f58723f4ce4f310646680622de4fd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6f62f4f2fc06f1cb30147da56b8fc88874f748262e4308b0d794c057267d9ac1);
            I9efcedaa1cc036ad8613f9ba801ca4ff4afcd709f5e4aaadbcdcd130d1263fc8    = If367e1e075614957d2fd83c76b45a3ebe11f58723f4ce4f310646680622de4fd;

            I2054d562a308ba04e604931976e93c9c55bbbc95d01e5504ab55ca3d8394f40f = Ibf421edf3110427df6425b33acef568cf41d337beb282e7b5c8d8a79aaa7a3d7 + ~I26a6366fb57427f6a0d87d4cff8a293a0752887e71b829e747c27980a1a3dbbf + 1;
            If5001dd5906be258a2388828d2ea764df15f9efd4d2ed03ef3182e4ad7f3adba = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2054d562a308ba04e604931976e93c9c55bbbc95d01e5504ab55ca3d8394f40f);
            I26dc2d992b646fe215751740a4406ce2a30e06fa2251f0382248aed7a08071be    = If5001dd5906be258a2388828d2ea764df15f9efd4d2ed03ef3182e4ad7f3adba;

            I3d365702f31c0b491b205449d36828e3fc8ca71d1e5b3ff872f9eda67fb06e39 = I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566 + ~I91c159ee16a42dcacaebf8cdac4c59d45d2e93735cffd86620ffaf2b859c8795 + 1;
            I499268c16db9bdcaf38ee694fa0269ae0c5ac8bc01e49cdc813244d8dd10c3aa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3d365702f31c0b491b205449d36828e3fc8ca71d1e5b3ff872f9eda67fb06e39);
            If25d531f7d1101b94167fde8f48549338e9b003202bc68bcb851f94fccb01007    = I499268c16db9bdcaf38ee694fa0269ae0c5ac8bc01e49cdc813244d8dd10c3aa;

            I9cb1f43022cfd63f00fe801b2d938c16277eefc9dde55af7c332011f60180cb3 = I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566 + ~Iadaa0bd11c77d7ea8c8cfc4b0c805c5afe6b75f597b03729ef2cb704dfe48286 + 1;
            I3f4ce0299be5d6b63eecc05da273fd2626ee66b8344d7cac0519c35643c8f487 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9cb1f43022cfd63f00fe801b2d938c16277eefc9dde55af7c332011f60180cb3);
            I3e49103842dcd70cc7795bfb356ef7d178c1e87d94c08cbef0794b0956dff7b9    = I3f4ce0299be5d6b63eecc05da273fd2626ee66b8344d7cac0519c35643c8f487;

            I1deac6b91e43b89f481b4b593e33836db7cc46ab37edca0ff7eef8ad6b92789a = I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566 + ~If8ea1abf5aef298950b84058c5e76029f717309fa685556f09c32b72959f648a + 1;
            I1894f875406842fcd82bee8824917bd78a61df725b719ed831ca04d6ee0845ca = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1deac6b91e43b89f481b4b593e33836db7cc46ab37edca0ff7eef8ad6b92789a);
            I84b78cf1294735491099a4ece1a26f5a1bed53ffd09724d3383bc63756866721    = I1894f875406842fcd82bee8824917bd78a61df725b719ed831ca04d6ee0845ca;

            I6896936df9cb439a07c80302e95b21023dc476bd78f678e93c7ecf5e3a159216 = I71d8be0ba8a91c324d8aee936676fe9e3a16fd14e44e44de643aa74fdeb35566 + ~Ieb5560e3a4f6a9c4543d941ac57bd3805afa7fa17624e5739e8e639e8d0d0c5f + 1;
            I8f3d1beef9bff167f3b3e18f1121ad15059b6030ace5b42de03ffd20167678d7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6896936df9cb439a07c80302e95b21023dc476bd78f678e93c7ecf5e3a159216);
            I964fe2ac03da8dd1965fd87a79f3fb2adf8e1607b64404233c3a09867227531e    = I8f3d1beef9bff167f3b3e18f1121ad15059b6030ace5b42de03ffd20167678d7;

            I363b3334e1423f125eae3636a561c36eaa744a2c8c62718fbc648dac5ac407d7 = I8d320b2d799e480d78887d5a1483ff7fe5f1a986d75e808863a9085bfc3634fd + ~Id32cba1cfd5a10024378db5089213ad668054033f8614d1ae09b83fd483a25de + 1;
            I33e0fe9272640febb568aca8a4b79c740a030fbda58477f8c5314fe3dd6ffa97 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I363b3334e1423f125eae3636a561c36eaa744a2c8c62718fbc648dac5ac407d7);
            I58df6e4342bc054f0177b7c91a68a1afdac21b2d1d52434ef5d8272b92fef6d9    = I33e0fe9272640febb568aca8a4b79c740a030fbda58477f8c5314fe3dd6ffa97;

            I05044427a4868a31ef17917e7795eeb32270ef20859f5d3d4699fdd408c210a2 = I8d320b2d799e480d78887d5a1483ff7fe5f1a986d75e808863a9085bfc3634fd + ~Iecf240e8fe5f620bf43121455ba23a715b23f53e049d2a36f4bf52e2a061a8dc + 1;
            I9f8e0b3d76f589fcc9b17b95c68db92dbbe51ce063ef7ae57c527dae2bb92b50 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I05044427a4868a31ef17917e7795eeb32270ef20859f5d3d4699fdd408c210a2);
            Iac61de7786d6ba1a40fc62f7d70b3cb366469c6674ebc4ecdaa21346903a58ff    = I9f8e0b3d76f589fcc9b17b95c68db92dbbe51ce063ef7ae57c527dae2bb92b50;

            Iccd6dc287621f59bfd5a38c0a5f5a06e1195d0d5f465e7129b782ab12f8e01d2 = I8d320b2d799e480d78887d5a1483ff7fe5f1a986d75e808863a9085bfc3634fd + ~Id1b9b5118024dfae0e058f5418c9e988e0a5a598ef7553947de6f92cd7399201 + 1;
            Ib3c97690b15aeae251f2ecc0b59366eede5e54cc23f96c5f55a04866d540dabb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iccd6dc287621f59bfd5a38c0a5f5a06e1195d0d5f465e7129b782ab12f8e01d2);
            I3c94620659b19b26861b2f4dc674bd9b9ddd8a378f11b67d27bc0f7639e0842c    = Ib3c97690b15aeae251f2ecc0b59366eede5e54cc23f96c5f55a04866d540dabb;

            Ie388d32b93fe9ae25426208c96be3b8dc61e43e909c7d28facb3fae96dc366bb = I2de3b409715599c65489338e9218150f6c33cd987ece5fdd9c7b2ba5c06d3d60 + ~Iaad1ab5e7603d5441b228c5e899eea7781b6f486b836a7b662f38ea832c1b8fa + 1;
            Ia53a9dac8ef5ed6ca6e7d4a8e3ce09c23057963286442c6de8154990774e0c50 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie388d32b93fe9ae25426208c96be3b8dc61e43e909c7d28facb3fae96dc366bb);
            I4aeb03994ab1826b4bc249e1cdcbda394b864bcec0ca3bd6a0897fafa6d280f6    = Ia53a9dac8ef5ed6ca6e7d4a8e3ce09c23057963286442c6de8154990774e0c50;

            I076abe19140e558596312bb8ed87bfb0490feda6f1ef7c0ac1df979cbfec7c06 = I2de3b409715599c65489338e9218150f6c33cd987ece5fdd9c7b2ba5c06d3d60 + ~Iecf3e0156bbf76dff96948ab7bf67772773b6bd62bd0e0fbc86a6eea8b05d4e1 + 1;
            I8baa541fc5fd694b934bb04d8be6893f071225e454e095c6a69340d24c29abee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I076abe19140e558596312bb8ed87bfb0490feda6f1ef7c0ac1df979cbfec7c06);
            I4d24219bb14476929c0d4b4bbef3ecee057061ad24af5601a8de67871680ee10    = I8baa541fc5fd694b934bb04d8be6893f071225e454e095c6a69340d24c29abee;

            I7a738dfeb0fa39730802cd687a42613f8ca1967c0042bd54b092c2e36abd47f5 = I2de3b409715599c65489338e9218150f6c33cd987ece5fdd9c7b2ba5c06d3d60 + ~I50e1a6fdaffcdf8fa99074f4480dcc21971ba8f5747b24a33232f9152b07af1f + 1;
            I47904cac869d3172932ccef3ee79eb5e70fa1dedbf4887d2f23fc54456756d7c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a738dfeb0fa39730802cd687a42613f8ca1967c0042bd54b092c2e36abd47f5);
            I6729f7458757e512a921fff6abb9aa05fb498db59115c3b041bad959c15fad3f    = I47904cac869d3172932ccef3ee79eb5e70fa1dedbf4887d2f23fc54456756d7c;

            Ia3ab7d65dd9be4dc787c343b0e877e40ad8b5ce9299098e4f9cb86ed25fe1d1f = I56c293e90676ea7b55934e3064087e3a4ea95a1c6ee3bd4d606afabce05357af + ~I317bde7e15c3a4d1456e9653a45d4d574509cca539be5c064af2ea89db634f45 + 1;
            Idb2735bf9ba202c3ffb7d50c14e63bb88305bae465a10fd9df8e1a516569b257 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia3ab7d65dd9be4dc787c343b0e877e40ad8b5ce9299098e4f9cb86ed25fe1d1f);
            I543c9825f790b1e9264e3f6b5e66e64c773dd0866bda372b2eda0201910105e9    = Idb2735bf9ba202c3ffb7d50c14e63bb88305bae465a10fd9df8e1a516569b257;

            I20dcaab9d6a12d0b868ac37762ddbbf0199ab0aab46594b5775a27656ff61d80 = I56c293e90676ea7b55934e3064087e3a4ea95a1c6ee3bd4d606afabce05357af + ~I84cdf374f692a63dab22cd91edd4f71e1aff29b51b06f0bca914f92407bea09d + 1;
            I36abf86ea52d7dff510cd8b2223acc503829bf031477a5fb94f6cbeed88c1929 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I20dcaab9d6a12d0b868ac37762ddbbf0199ab0aab46594b5775a27656ff61d80);
            I8097cf47b760092e87e117165f17e1f66afbaa3ee78160fd0e2a597f613883ee    = I36abf86ea52d7dff510cd8b2223acc503829bf031477a5fb94f6cbeed88c1929;

            Ice4daffb593d295aaae1b2165bc2dc9612bf70ee6005a4200f764c76c430dc32 = I56c293e90676ea7b55934e3064087e3a4ea95a1c6ee3bd4d606afabce05357af + ~Ieb31a59d63544ea160d3934f0e38e6333f8571e77352bdbfd338d68c437f02b5 + 1;
            Icb48731efd9ce27f84725ef47b1e6733a95b4753274e4dbaef808d4764a470e6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ice4daffb593d295aaae1b2165bc2dc9612bf70ee6005a4200f764c76c430dc32);
            I4eb210e31e4ad434958f477b79dcf5b2694caf5c18f801a8d3b3b612eb0812af    = Icb48731efd9ce27f84725ef47b1e6733a95b4753274e4dbaef808d4764a470e6;

            I6740d7cf9a56e745fd86c9131b62b2dba6a7ae614338a59607a43f0b77d9bda0 = If32e43e89968b9f008cb77759dc7047519d200c512cb11c105b74c404603fc79 + ~I953a4a4cbd4e6c0ccf4880cec5c947f86d6542f9a7f125d7c8cd71f8665b9ddb + 1;
            Ib45b2ba433dbdf77fdf6bf72c9e7a1b60d7bd8977c20cc9ae07e7320c058252e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6740d7cf9a56e745fd86c9131b62b2dba6a7ae614338a59607a43f0b77d9bda0);
            I40b6ad89db699e7f672e55f672bfc979d85a462330e526aefd63b9724ff7de89    = Ib45b2ba433dbdf77fdf6bf72c9e7a1b60d7bd8977c20cc9ae07e7320c058252e;

            I10ad038fb26d337df3013912d38403548cb5e12d6e175518ac7e924e583e1fab = If32e43e89968b9f008cb77759dc7047519d200c512cb11c105b74c404603fc79 + ~I5b143cf694d99dabce0cb40d2d689fd7232531ab3a30888f811171b6aa2e024f + 1;
            I30cb24b52e864de98a09fc41e8719f6009e8642027c70850c80dd90844b08093 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I10ad038fb26d337df3013912d38403548cb5e12d6e175518ac7e924e583e1fab);
            I014e96c75acbbe2bf38e1c89b52e1a331eb3d31b984a67946eef2a5223b87855    = I30cb24b52e864de98a09fc41e8719f6009e8642027c70850c80dd90844b08093;

            Ie103edeedef5ea626306fe0162187acb812025558381c8ff0ca8bb006a2caa17 = If32e43e89968b9f008cb77759dc7047519d200c512cb11c105b74c404603fc79 + ~I81e45b654bee6c74edb5e034c89bed7151c60a69b554a35710d1b173fe45ea22 + 1;
            I62abc4525f5ddd159fd9af8e17f6b7a271d8aa70617eca684129eb9320ddefeb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie103edeedef5ea626306fe0162187acb812025558381c8ff0ca8bb006a2caa17);
            Ia3588e449670d7edbf99e52ccf0d7c8462b51e3d24ec5f0f7293290d47154f72    = I62abc4525f5ddd159fd9af8e17f6b7a271d8aa70617eca684129eb9320ddefeb;

            I082f12331831c80bb11a3660e45ab9fa6c122af71c82374eb645f01f89b03a15 = I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0 + ~If7fb04f8e3e8eaef8fcc0486d12d1e37a887bcdecb366c1e8b53a3e1cce0637f + 1;
            Ib5945692324b161750a7e5b6d9a2cba70565ddcb2f85ce9665da37e06c256ffb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I082f12331831c80bb11a3660e45ab9fa6c122af71c82374eb645f01f89b03a15);
            I6b3108db71d5eaffc5606fb88fe909a0462a77232258fd85cb6792954ad28c0b    = Ib5945692324b161750a7e5b6d9a2cba70565ddcb2f85ce9665da37e06c256ffb;

            Ie65f8e169c71198268320e9dea6a360718a61dfa0e33983344ab5070a97fe3c4 = I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0 + ~I8e95ffa3fdf70dc76c935f7d4dde6f39dfba8eb795f7ccc55510ab3caf678410 + 1;
            I3fc3cc1b4558877a3148d5567d5e5ef929459603af3c07214d2a05a5c9568e2c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie65f8e169c71198268320e9dea6a360718a61dfa0e33983344ab5070a97fe3c4);
            I55a1e3e076ea304ccd72b18524bfa076977a0f791806719d752ed020cb6c3e37    = I3fc3cc1b4558877a3148d5567d5e5ef929459603af3c07214d2a05a5c9568e2c;

            Ia1df41c6fad9069c1aab753a907bce8625c2d114c156b2e2c0429d7df6c30f17 = I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0 + ~I31734ccacbfeb8a5c0c30cfc84934f8d1636ce4ecae14fe7809d6aa8df35a9e8 + 1;
            Ie399b6c8ee179bfbefe764089dd280841d5e8bfa73941f40de3d7a293c4618fc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia1df41c6fad9069c1aab753a907bce8625c2d114c156b2e2c0429d7df6c30f17);
            I318f0ddae7fd42b63d856ad6923268574eb4f8f71cbdddcaa420e917a1d7ea51    = Ie399b6c8ee179bfbefe764089dd280841d5e8bfa73941f40de3d7a293c4618fc;

            I2eb3b47e1f13607457b31a324a263038853d4c7bb85f4c9c00c26c16403dfa7f = I45c764e8eca9bb32e03823ed07fc80d211842a86c1f6b1551def3864b79993b0 + ~I5144a2cef7d82b7a91f9d83ff8fdea356bb01db215bc167f0c498d55d1faa622 + 1;
            I0b0bec74dc25dc927944819c56c35d1df298227cb0fd804ca1b526db544b17f9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2eb3b47e1f13607457b31a324a263038853d4c7bb85f4c9c00c26c16403dfa7f);
            Iee19c6e30e6fb9258878db36251e2e15a071b41364b59473c9de2c0f0b8c9ce8    = I0b0bec74dc25dc927944819c56c35d1df298227cb0fd804ca1b526db544b17f9;

            Ia556763bb9b39f7ecdea64ef734cbbbc108070aabd560d87872fb475201ee4b3 = Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931 + ~I8fe688adfc161cafc0777f3c3ac9ae27372603ec55cb3865f90f38f9dbb59439 + 1;
            I8007db0cf24afff18bc9922f5b33406c49079a0374944211f7ca69ed7dd8b4f9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia556763bb9b39f7ecdea64ef734cbbbc108070aabd560d87872fb475201ee4b3);
            I4a9362c36b4a88ee5422688ee5550c97e8fe10b4cc23b6538ee81bfeef1472a9    = I8007db0cf24afff18bc9922f5b33406c49079a0374944211f7ca69ed7dd8b4f9;

            Ic0d0d1aa735e38d8af824759f30badc83db776ac7871d2f5d0c12594b25342f6 = Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931 + ~Id2dbd07db2080c14fd0026396339e31183fb5bb6a476999102300cf81f34b93a + 1;
            Ia79976d64cb4e1c9a542747c4a7ae62fe509cf1f8617cff283529b36e86464e4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic0d0d1aa735e38d8af824759f30badc83db776ac7871d2f5d0c12594b25342f6);
            I9dda3335af58c2daa92010ef90e217e0842b7740a65ce2a029ebde5b65e9fc86    = Ia79976d64cb4e1c9a542747c4a7ae62fe509cf1f8617cff283529b36e86464e4;

            I33ceeaee9a8251525af0cb5b6c1b9968c58696493f1a3ac45cc5c0e3b44fd5a6 = Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931 + ~I8a61ed94b6198131fccf4feb6be7327f59408e9de4def9c4a155167192c5f065 + 1;
            I5889799635ff332461bf6d25cf95f401edf86feb687d4013457a3298dd943c4a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I33ceeaee9a8251525af0cb5b6c1b9968c58696493f1a3ac45cc5c0e3b44fd5a6);
            I996cd6ee71fdd8f4b109acfd52bf495951439b9e49b87a6db4565bebbc7d1e1d    = I5889799635ff332461bf6d25cf95f401edf86feb687d4013457a3298dd943c4a;

            I7453e7476c16ded7f06fcc1f9c11a504545e00d1e15faf2f2d0cfb57b9f35c5c = Ie4f7f41dd4e9dd1ae42d79cf0d2ac38d3101511a703635579a6910d6e1e56931 + ~I67484837f2e585fbb85de404cad8f08ba58bd1faa81b9931f88473d7f4a9a06e + 1;
            Id3f8872c22051e28cc6cb6beed2ec233c7d8b79ed058acc23d862b30f0104715 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7453e7476c16ded7f06fcc1f9c11a504545e00d1e15faf2f2d0cfb57b9f35c5c);
            I705cf789e535bcc9523034b7f4743daa8f66f1dfa3d15c77b87e9f1845563690    = Id3f8872c22051e28cc6cb6beed2ec233c7d8b79ed058acc23d862b30f0104715;

            Ibdd02bba3f13be2c6f23b969be65c45c5a1b1d42b06a5189c10b452af7b1e055 = I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164 + ~I3af3a7e6138910d118e49b29a6de8bb8e6fbd1cfe13549eb0feea6cd07e6865c + 1;
            Ic620c07652badc1f7831a4e487498f6f875cc1d9c29604b1991dc89620485abf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibdd02bba3f13be2c6f23b969be65c45c5a1b1d42b06a5189c10b452af7b1e055);
            I4345f323dbf4da279580851ea1d0b7a2e5109f518ca914c88b6ac91e9ce8625c    = Ic620c07652badc1f7831a4e487498f6f875cc1d9c29604b1991dc89620485abf;

            Ic438ad9f1da18eb848fb486bdc7fef62f7a3ce12e948699f5aade5c2922e572c = I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164 + ~I7e12dde03af7a5ae0d05cdc9b29f31ef726c7bc51a7f07e374bfbc0846a24f0b + 1;
            I88787a9b8cae593784a9ffa45bb675bae477cadd18e0cbce021ecc9b4461dcea = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic438ad9f1da18eb848fb486bdc7fef62f7a3ce12e948699f5aade5c2922e572c);
            I8a484469fd2c86173f27a68b9ae6c15c3813761e5dc1035c2f9fe04b24a6d73d    = I88787a9b8cae593784a9ffa45bb675bae477cadd18e0cbce021ecc9b4461dcea;

            I7abea0145d10af48608127e2828ea265ca8883f1c43474ec82b2e24da693c566 = I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164 + ~I445cf6fbf071cc76e6fc981d7f2f201d0e09d3f47c1227feaac47fb57a14e85d + 1;
            Id093cb8cc2ca70696c70703a5a623de87427b286fe83fecbbe236110c68a8e8b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7abea0145d10af48608127e2828ea265ca8883f1c43474ec82b2e24da693c566);
            Ic6518d2e4de9b3feb98b24f5ff4fd43edb699fad33847f2e67ff731825f15177    = Id093cb8cc2ca70696c70703a5a623de87427b286fe83fecbbe236110c68a8e8b;

            I9aafd88945bf07d0d9b361fecf903a4c1b14db6dede3d95677ae0d01d0e36894 = I391c1ba9f97df92bd62c5f691e551697a2581de00ab8dbfadf28a270481ac164 + ~I4404bf7e923ee1bc0230835c00684d298572238aa8b9602dc48e177464224a53 + 1;
            I789fc42a39562699279fd510c6fe748b90314b0586a7e051058bad4b84370347 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9aafd88945bf07d0d9b361fecf903a4c1b14db6dede3d95677ae0d01d0e36894);
            Ie147f013af77ffb57ecdf0bac185fd60648505960bec48f3f18094b1b7e319ca    = I789fc42a39562699279fd510c6fe748b90314b0586a7e051058bad4b84370347;

            Ib7bfebc508c949b2dec0ac81a1029eac23947dd8b78872b238f1ff1bd0e19676 = Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e + ~Ib87cc4d1070a195aa8118b92d29d7c836685de2e44ba1b21388677c8e8a5fb25 + 1;
            Iae8a2a117b9f71a954b7368532a41c443d18950b56dcc9d12a7809dd4b6f9033 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib7bfebc508c949b2dec0ac81a1029eac23947dd8b78872b238f1ff1bd0e19676);
            I0a51859ca31f0b470011ae2b3bcbd11fd2c79f03c854103f016b54af79028ba1    = Iae8a2a117b9f71a954b7368532a41c443d18950b56dcc9d12a7809dd4b6f9033;

            Ibcfce28ff0415dd2da98a7ec1b48f013c33edb8b6224ee7637478da2889b6b16 = Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e + ~I39249b7f0d22c6116a7dfd0c0748123ebb6a9b7f931a492a534702157ab28c3c + 1;
            I386d1bd1bbf4aa7d9ccbe2cb4a9dbd9cf9bdc1fbccbac9039b32d0082f2442ee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibcfce28ff0415dd2da98a7ec1b48f013c33edb8b6224ee7637478da2889b6b16);
            I1f5d36144836b1c2e41164adaa02934f77b47f317c3f6e7452ea483c756b4ba3    = I386d1bd1bbf4aa7d9ccbe2cb4a9dbd9cf9bdc1fbccbac9039b32d0082f2442ee;

            Ie2c653cb0d05e3e9f884f7e78efe071774cebd49008f86c8106fb180e8196fff = Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e + ~Ibca42a442c971d363e4f848d203d2782af05ddbaad93e8cbf334328d94a8a499 + 1;
            I588bd9ed21e23969799b7c1ec15350266ba52e0eeacb1bc20803f8aefcacab6d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie2c653cb0d05e3e9f884f7e78efe071774cebd49008f86c8106fb180e8196fff);
            Ie1c46630d4cd6028c341687f4df0c2220054b63f8263fab4a11d3ad89f6518cd    = I588bd9ed21e23969799b7c1ec15350266ba52e0eeacb1bc20803f8aefcacab6d;

            Ia709de664b32e0acc613ab7448eac9837c7cb75de3469262a56bf32086894ab6 = Ib97e33c792a31c802cfd7dfde8e716d3084b7ef8b98b83e085cb6d8c3a56955e + ~Ied796eff44d61681c5d5de05933e785d387a97b2430fee26d96b0b24a1a54c12 + 1;
            I7045e20c9bb1e7137b3c996fe61c7aad0323741b7b5dd70d8fe2ad840a816000 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia709de664b32e0acc613ab7448eac9837c7cb75de3469262a56bf32086894ab6);
            Iedab2e8aa599a943abe7d0d1dabb0f7a5a7d4b97f36e982d5f548a4acccfe2c2    = I7045e20c9bb1e7137b3c996fe61c7aad0323741b7b5dd70d8fe2ad840a816000;

            I3feefae60ec0eb2602217fb4db5cb7bb3d4af0e5d6656f09c286220f83c14e95 = Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a + ~Ib0978aef78ec9b21853831a81aac1d87a2410594c7839432302eb5fa99a4c0ca + 1;
            Id056954ad6043df8f15fdd039c5180035a585020638d2e39e1e1392e283942a5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3feefae60ec0eb2602217fb4db5cb7bb3d4af0e5d6656f09c286220f83c14e95);
            Ic7ecf5c9528425bf54c120398b0e5f75dcd4acd18b3088fd8a16fe8207a592bf    = Id056954ad6043df8f15fdd039c5180035a585020638d2e39e1e1392e283942a5;

            I588d1fefd4585f5eccaea213e11f8d74f1308c3bb15bd7e88dd5275ef62e236b = Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a + ~I7958c747e1ef37e2995c52178d143af6a5f3acdf7c6d1cae518c82653ec18716 + 1;
            I213da828cb42a5d0f9025d51b36ddb92a677c7878c1f99496cf0c921bb8674c5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I588d1fefd4585f5eccaea213e11f8d74f1308c3bb15bd7e88dd5275ef62e236b);
            I355cc82d012dbfaa00529a9197d4fe0b654fc609360a0775d398ae0b3e95f2cd    = I213da828cb42a5d0f9025d51b36ddb92a677c7878c1f99496cf0c921bb8674c5;

            I211af75e159531ef945adcb8f51b79d5b1f27ee3835f2cc2f79124b235c10a72 = Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a + ~If4927b8f31777ef2940c413336113e906e0e3556c31b9b3233107b88b1d71999 + 1;
            I74a97e7cb539a14631bfc8532c9903e23e1889323443903126eefa3bc5e5be05 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I211af75e159531ef945adcb8f51b79d5b1f27ee3835f2cc2f79124b235c10a72);
            Ic0c2a03a257040df478653886a3a2400777322b4d4333c0da94211227433697f    = I74a97e7cb539a14631bfc8532c9903e23e1889323443903126eefa3bc5e5be05;

            Ibd0e4e5d04591535c937a5389e0763279d4c267e0d0d7f1256a9271d49892307 = Iaf74d4f6fb5e4caba7329211ab0e6186a7c5ce32892caaa7accfc7f5af2ba81a + ~Icd8838ebb43dad19fa96e741b32851dbaf5c469e0591a1231898a7aeb6ecc788 + 1;
            Ie31f193f6b43563eb5a1cc4fac89514b8e972743354f7a28c0b6c8c8e70f1799 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibd0e4e5d04591535c937a5389e0763279d4c267e0d0d7f1256a9271d49892307);
            Ic09079bc0fb0e140e7285e2e5af8caa802db98a774db8ce0bc5158e08becb4c1    = Ie31f193f6b43563eb5a1cc4fac89514b8e972743354f7a28c0b6c8c8e70f1799;

            I1857bbf85d1336737426b53588e78aa34ec0664ec1f3c4bc351040782a0c1719 = I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980 + ~I9d56c14b3465733b5c5fbff528a7a7d85c918a857257ba8e302ae84a0f4734de + 1;
            I3a3a48d2c08ae2a07dc1e291c0d51c6e30be91af52aa6a439849005a958540d6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1857bbf85d1336737426b53588e78aa34ec0664ec1f3c4bc351040782a0c1719);
            Ia7d33f990e505c818a46c2a54c13bd6680e3a34847708d89ee6f38999242e0b4    = I3a3a48d2c08ae2a07dc1e291c0d51c6e30be91af52aa6a439849005a958540d6;

            Ib5b72b3ca0b1aa00d12330c72c5435ad4ca90d598d05e7790f1da65af2f8c3c8 = I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980 + ~I80c4eccc6e6be84f8936ed3e9a9457a862eca015298ba2db70745f25a65a6571 + 1;
            Ib93a5b2f4b149124dc2bdc6a90438a5bddd75a83c0717b52fdb47de0cbfdf8b7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib5b72b3ca0b1aa00d12330c72c5435ad4ca90d598d05e7790f1da65af2f8c3c8);
            I0c87558b4bcfed105da91186dbea82b0f8d38c2473b578fb874ebd3e844edf51    = Ib93a5b2f4b149124dc2bdc6a90438a5bddd75a83c0717b52fdb47de0cbfdf8b7;

            I24f30205c1eac80e3a167d5b52d1328285db573a6671ad7e635e47f49646d05c = I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980 + ~I18eefcf5075eee79120ffa0e5875cbe7632d1db84b1c498107413f14b72820f1 + 1;
            I76e90676f89b877e33f8c96e6fd6d2f1c2da1fa8602fb65bf8c1aa18d8b6269a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I24f30205c1eac80e3a167d5b52d1328285db573a6671ad7e635e47f49646d05c);
            I5a7f5ab868cc2f4e823808a238df41f5e29c98d896557abab5eb1b5ac4231eeb    = I76e90676f89b877e33f8c96e6fd6d2f1c2da1fa8602fb65bf8c1aa18d8b6269a;

            I26ce0fefb116238e66b72d526766ce8f9b9d1de0df15d835668d928384e44827 = I4fd1c7608cf05c2a4343174d4aabc9b585e70dbcee50916aa2f9df88b8224980 + ~Ic6d60bc06b0eb51b5ff4b8cc0d0ccf55fd8e5c53aab23b3994ca8d094920d619 + 1;
            I7d7cad2d595d0e7c85112d240714aa5ccb684bac4b8fb57f4e8118890ae82063 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I26ce0fefb116238e66b72d526766ce8f9b9d1de0df15d835668d928384e44827);
            If3574e7d834ff9a2b7247d3262dcd4265a5aa04a73495afc4e8098f7da4cd0ce    = I7d7cad2d595d0e7c85112d240714aa5ccb684bac4b8fb57f4e8118890ae82063;

            Ibada8912d6b4053809b28c28b01acb109cd1c80309a62b9b5b8ae3b5a0ecc44d = I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7 + ~Ice9dcc5d9ccd6caf90dda22be9ce113c53c7eb492cfd5e0b237da4f92aac2d7f + 1;
            Ia153e17a2ae12333c7982319dad7b3d57721e5e6075d2ee89f61dd6c8b06f73f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibada8912d6b4053809b28c28b01acb109cd1c80309a62b9b5b8ae3b5a0ecc44d);
            I5187aa2268c0345b27861b3f411a57adfe94104cd1a48c7573407a0f79e345d6    = Ia153e17a2ae12333c7982319dad7b3d57721e5e6075d2ee89f61dd6c8b06f73f;

            I698dbb248637786ce7fde5591c80178aa213872056e5fbcb46cf7a23484143ed = I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7 + ~Ia2aece9bdb39e997b99e491171667091adbee475ea9b1c372ebbec109f9f714f + 1;
            Ief4ea9c80ee182d2353b1a258190c80085fcd78a2379cd59968ade8f12695d20 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I698dbb248637786ce7fde5591c80178aa213872056e5fbcb46cf7a23484143ed);
            If54927516082a9fec583e3cdeaf09539203d2f351771381d6c29c7961dc6f98a    = Ief4ea9c80ee182d2353b1a258190c80085fcd78a2379cd59968ade8f12695d20;

            I0d5b3b10a05b9ad2d2df1d67a669cf252f9dad522d241643ad3ed51b610a32eb = I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7 + ~Id059fc689baea934a9f278b1066a92d6aff850608c0797dd7257693cbfa40102 + 1;
            Icacb23d3c6ca588b3fbe8371627f9c6de649dc63ec23db2a94d3b532660a8a8f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0d5b3b10a05b9ad2d2df1d67a669cf252f9dad522d241643ad3ed51b610a32eb);
            I8e63aa98e26c7163ac7e004f9b363177513859fd81ce1d6be355e187166ee55a    = Icacb23d3c6ca588b3fbe8371627f9c6de649dc63ec23db2a94d3b532660a8a8f;

            Ifa2c9985b7daec8d06c292ca451d71e14a32aece2e26dd6d5ce3f102d70ed54f = I8453673fc6dbbdf92d73e5b2c333ac1c28f24a4ecc097e559e555c59d3b0bca7 + ~Ia0feb2870e46760bd3c58e5af56a40a73fcc6c9611766c77c4784f88c35f440e + 1;
            I5902d24b66bb202f53e54816fccd38cf887dcd18bdf15dc6893dc55bcb6ad9d8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifa2c9985b7daec8d06c292ca451d71e14a32aece2e26dd6d5ce3f102d70ed54f);
            I6e3f1705d8ba2b2cbd6b7749bf249716ede50edeca032e277396a885c69399ef    = I5902d24b66bb202f53e54816fccd38cf887dcd18bdf15dc6893dc55bcb6ad9d8;

            I6f84b4bab9b97d15495d515da0fa036b9ebc5a7193c2544274b3121dc23b8ae3 = I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6 + ~I908d977677aa9b15536027b54cf497ddb8741b339748986180944418fd848448 + 1;
            Ife31d9500920174f7dda41fc67b6e54774505ed3c35a04eea45ca45b8be20457 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6f84b4bab9b97d15495d515da0fa036b9ebc5a7193c2544274b3121dc23b8ae3);
            Idc29a95902384ae5ae3858cc3583cfc2fb39d4634b67c3c9858b9b6b9468fc87    = Ife31d9500920174f7dda41fc67b6e54774505ed3c35a04eea45ca45b8be20457;

            I922ca03f57cae28107251c50af6bc0b96a46be661f758e93f2b80d0c23bcb02b = I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6 + ~I050437a5474ba60337593b28d17e2bec5c76d26ea8afeac61be93e8ba0ada42a + 1;
            I658eeaa8e533a4e2fff6e0c78b3d12aae697a38c0ae02a835e4c62eebe7d946a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I922ca03f57cae28107251c50af6bc0b96a46be661f758e93f2b80d0c23bcb02b);
            I3ee26418f368f28b1dbc386529fe4d0034170fceeaa1cf5f4edd2132db250ab6    = I658eeaa8e533a4e2fff6e0c78b3d12aae697a38c0ae02a835e4c62eebe7d946a;

            I60dfd53c9dda263ede70e2debced85d2e29fb7f897347d5fb6bbe068b5d42b6a = I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6 + ~I4c5882b979d1f315e20e4a8fc06c794c0217b97de2613e193cb7a213c2119c97 + 1;
            I77cfd243c2c2f87ba6a4f19612488bb84593524abb103ab9808275bb0a3f3c09 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I60dfd53c9dda263ede70e2debced85d2e29fb7f897347d5fb6bbe068b5d42b6a);
            I82393d9631be548b7d2f25eff102ffad6a2a1b7a683c82d8046dfd07b66e26a3    = I77cfd243c2c2f87ba6a4f19612488bb84593524abb103ab9808275bb0a3f3c09;

            I4b915b467967001eb1ea2c496d782c2fa9506073cc4441ca6cc42f67e57ae822 = I9b402ad8da7585113ba25bb83542391c4bc0a631e32247daa578dd9c4966e2a6 + ~I60b4f2cd3f513ded6891a6506d0ec74357660440c94e62f4f7e2f886c1233204 + 1;
            I2fc93ebc02fddfbbe5a6cf5bb7aca44f0a664be4a2c8273ac638ff7f94c3b896 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4b915b467967001eb1ea2c496d782c2fa9506073cc4441ca6cc42f67e57ae822);
            I61291a36d4d546d1cb7c79a8a8c9ccbb4da2bf3fe853e05a56296804d5fde212    = I2fc93ebc02fddfbbe5a6cf5bb7aca44f0a664be4a2c8273ac638ff7f94c3b896;

            Ia556ece4fd10276fd9d7e0b3bd79ab15221b0891dfdcaa8a3d3f0988a356b78c = I1ee241dd9ec346bf09b25ccd2f1669be719a1411914d367372a46c8d60cb0f44 + ~If7c696b260799e0ccd86bb377086dd1be59c9d94754dc52605d659391439d3d5 + 1;
            If8fd28316f1fd0fb493c897bdf978233c0a1bec3cf2136146e8471b86e0c0f67 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia556ece4fd10276fd9d7e0b3bd79ab15221b0891dfdcaa8a3d3f0988a356b78c);
            I454cdecfffd5c06b833e81e8990b07a9b326eec23f31a7b6589b969f610d8ed6    = If8fd28316f1fd0fb493c897bdf978233c0a1bec3cf2136146e8471b86e0c0f67;

            I9dae8c584ed5197edc44374d711497fb81a91de44e3cc12d23de36f3269fdb65 = I1ee241dd9ec346bf09b25ccd2f1669be719a1411914d367372a46c8d60cb0f44 + ~I96ace764b2f8db5049595445104a408a641999152f2a6c63d22bc6946c27322b + 1;
            I2452b31eb1cfee03ef6f6c00ed42126b741fbdbfd43b74377a675383e146ca22 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9dae8c584ed5197edc44374d711497fb81a91de44e3cc12d23de36f3269fdb65);
            I0d0472e7c0ef483f8cb46ed393b7bcd5ea93f12dc2885368d5bf587c24198980    = I2452b31eb1cfee03ef6f6c00ed42126b741fbdbfd43b74377a675383e146ca22;

            Iaab44235fea66a54e56d75bf5d2732a95042c033defaa2a906b2390bdafec03e = I1ee241dd9ec346bf09b25ccd2f1669be719a1411914d367372a46c8d60cb0f44 + ~I90b9d06240e2a49693ac4ebe37203439a157a38d068e630c45341d7d677b816a + 1;
            I2117d5fe8b672b3eaa3c257a2a7df3819e54d86ca29f980dac153f8a9da37607 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaab44235fea66a54e56d75bf5d2732a95042c033defaa2a906b2390bdafec03e);
            I33dc9b3b4f5aac0a30c5ab73b222441f5fbeedb26b7b8749a0ab253f239598d4    = I2117d5fe8b672b3eaa3c257a2a7df3819e54d86ca29f980dac153f8a9da37607;

            I0a2d4121a3aa27634d62a6eab291465d8c2ac688a263dfa0d3fa9e007d825aca = Ia34cf7cdac966a47b902c17ef799ca34f3c17e4f5a410b97d7f07933b977db3d + ~I55e293b2d9539b16ee0f135097b8ec02fc9af54fc96ec3a3058af417b0d04e48 + 1;
            I90c54ee94f70ae9ae84529f1c52175bf663de85a58c8ee420146322ee9faf1a1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0a2d4121a3aa27634d62a6eab291465d8c2ac688a263dfa0d3fa9e007d825aca);
            I70ea317892671f95b146604245efea2c83830d5e6b03a1dd19f2ecb28b47a9a1    = I90c54ee94f70ae9ae84529f1c52175bf663de85a58c8ee420146322ee9faf1a1;

            I4643ca0b8bb8f9d58565dac92705b1e6ef755a8edd307a0105482001c06eea13 = Ia34cf7cdac966a47b902c17ef799ca34f3c17e4f5a410b97d7f07933b977db3d + ~I84744085fa951f13f4fef6c44fb0180e543fa6793e89f4dcb14c3da6b27105b0 + 1;
            Ifdd6eaefa7e96076232a2d0f399e537f2eae4cf57a837693be785373eeb8f160 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4643ca0b8bb8f9d58565dac92705b1e6ef755a8edd307a0105482001c06eea13);
            Idf920a1de857f846c8ab2646a68ee3a6053d935968cdc3d6b46308a473be4099    = Ifdd6eaefa7e96076232a2d0f399e537f2eae4cf57a837693be785373eeb8f160;

            Ib13dadfd1a4c8b6664863bff922da75c848e4e114e53ca32d4b93537cffe3fc6 = Ia34cf7cdac966a47b902c17ef799ca34f3c17e4f5a410b97d7f07933b977db3d + ~Icc84144f0fef09379e456de5410487e7882d373874a686f1b61db92511a91e2a + 1;
            I939c9cc4a14510cd9b1d69ec5f5649e80399a13c355e0f8bb8a5cda6df224e8d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib13dadfd1a4c8b6664863bff922da75c848e4e114e53ca32d4b93537cffe3fc6);
            Ifade018f22d237bddeb6fd8736ba424241846d20f2f32d2bb7fe779462ed7261    = I939c9cc4a14510cd9b1d69ec5f5649e80399a13c355e0f8bb8a5cda6df224e8d;

            Iba4a2105d76cbbbbba7cd474dff95136225ada8b4e62e607962200b0caddacef = If017b6342521fac4000803837465d5793375e9f4b8c2d9fda18843ec7b9e0752 + ~I8dc734304648fe3fba1dc7108e8697cb88b61a2ffa704491b2b9df8cc8354825 + 1;
            I8292477c74597003a879f491614abc033a2366dc024d96a5b38edc6517561f4c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iba4a2105d76cbbbbba7cd474dff95136225ada8b4e62e607962200b0caddacef);
            I9318e8402c23072dcc49ace45bb9814c535167574af63bc61463059dbcb0067e    = I8292477c74597003a879f491614abc033a2366dc024d96a5b38edc6517561f4c;

            I0a34efae03321f53acc6f183e7c3f22df19d0a0add67ceb5edcc38046ec33748 = If017b6342521fac4000803837465d5793375e9f4b8c2d9fda18843ec7b9e0752 + ~I701aa61e04d2787a36f529185ddcc94c832834d38ff92b37456b64ce46c69b2e + 1;
            I0e9f54539d4a95d17f80a316734c90dbf2799dd8311c6bdf7cb06d100d576254 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0a34efae03321f53acc6f183e7c3f22df19d0a0add67ceb5edcc38046ec33748);
            Ic0071db5dbcb92ea14e4b31a24b9f9febc208bf86bb0634f07d9cd3763461055    = I0e9f54539d4a95d17f80a316734c90dbf2799dd8311c6bdf7cb06d100d576254;

            Ia3189d8c7911fc25a6079d7e30557a3b7721d0ac84c03b38366c1db55c1d3f95 = If017b6342521fac4000803837465d5793375e9f4b8c2d9fda18843ec7b9e0752 + ~Ib5ba52b9ecafcedb064e66c38273f7833d0b6d0239a7fff9ef3a0e30d0f77dc8 + 1;
            If475d646e4baffa57990168021c33001ce2c5d28c7f22a83d42e35b6fcf1bd22 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia3189d8c7911fc25a6079d7e30557a3b7721d0ac84c03b38366c1db55c1d3f95);
            I64cc4cfd27023e75e5cb557e7bac31506d466107aa2cfe7809e148d8977f8393    = If475d646e4baffa57990168021c33001ce2c5d28c7f22a83d42e35b6fcf1bd22;

            I98c91ea87b40d44f2e5830fa4e4b285baa5cfadd6d5419e88936592f664d8340 = I8bc9b50c83facba8db598d0c5c71cf811e181fd16038a08f5aa04f00ff2bed87 + ~I6dd215113f113a81bfa59464b587ae7c95f02c1461664fdb818ce751c240b96e + 1;
            I0122a25f242d23f81bd7c99bb094666594eb9c2ba1ebbfca379b384411257045 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I98c91ea87b40d44f2e5830fa4e4b285baa5cfadd6d5419e88936592f664d8340);
            I560502a76e2a6f15d91f55a12133213d8896b50299e0a7ed30c5c5958d5f5ec5    = I0122a25f242d23f81bd7c99bb094666594eb9c2ba1ebbfca379b384411257045;

            Ic458bce5868967b65093883a779b50f1d51fd9fb924eb6bdb9933db186240445 = I8bc9b50c83facba8db598d0c5c71cf811e181fd16038a08f5aa04f00ff2bed87 + ~Ia57f6e4dd9ce4389f90c78df4fca73a681df346f58a85f61a74e842427848347 + 1;
            Id0e600a5ace87e9d404d63fcecff3d7a6b212ae81456381885943b78b98aa2aa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic458bce5868967b65093883a779b50f1d51fd9fb924eb6bdb9933db186240445);
            I7813b9f4f76a24bbf99a0f2d9cfe1d3a53eb0ec0fa5c72e06f1f86fdd1801c56    = Id0e600a5ace87e9d404d63fcecff3d7a6b212ae81456381885943b78b98aa2aa;

            I20382630b2daac9cb982d267670777192b41ca7e729303eb524e38603f056031 = I8bc9b50c83facba8db598d0c5c71cf811e181fd16038a08f5aa04f00ff2bed87 + ~I38a6e64d23e0dc1a449445bf10e786777e978aeab68b3a99dc5335b93c67da45 + 1;
            If1febcbc92a43732fd85592bd9013cf0e14fd0e3926826badba0e53cbcdec1fe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I20382630b2daac9cb982d267670777192b41ca7e729303eb524e38603f056031);
            Ia81295e4b9400e1737a8a8d335ed9765fbb59b817f0251f1f032ba3e48c6bdf3    = If1febcbc92a43732fd85592bd9013cf0e14fd0e3926826badba0e53cbcdec1fe;

            I8663595964ca4eb094c6cb80c0eb4ad319673883a254ccc35cc4be73ea5bb00a = I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c + ~Iabfa5de761b3413904b919f913ed73bf27f5249b7dc6bf8471a23f06a30431e1 + 1;
            Id88407a8f20b0589f462959accb7d6737ae4c244083469d5207033ff09f7eb89 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8663595964ca4eb094c6cb80c0eb4ad319673883a254ccc35cc4be73ea5bb00a);
            I0b7c06b48a33586be508f2334fc3eac5befd9ff87751db1859c5f01cc6d44b15    = Id88407a8f20b0589f462959accb7d6737ae4c244083469d5207033ff09f7eb89;

            I8192c0915a9b5e00cb68ec0dd1c26b26640f3f9c6e17e3de938b91fba44e3782 = I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c + ~I9f08c1a4053ac65909c96d240c83e15017c81fa41f351b0a707fb7882e49f4c7 + 1;
            I0b7fce50c3bb3677721cd1cd0867a43bc7e7d172db559dd6e92617f65eb3184a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8192c0915a9b5e00cb68ec0dd1c26b26640f3f9c6e17e3de938b91fba44e3782);
            I63860f7f2cc2e0814f98ead1e90694f745ef7a70e90f0af487d002ca46bf2c57    = I0b7fce50c3bb3677721cd1cd0867a43bc7e7d172db559dd6e92617f65eb3184a;

            I886c2494bdc82c917ee66135ce52c761c347c8fe42ccd63d769cf315b338f2da = I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c + ~I6a5f07e66bbd7e05ab9c5adc7bdc99f269386519a6212431d5793e766239e862 + 1;
            Idba8e69c73d0fb1bd1aeff84e1c6d06234801f1b37b84ce20a98d29b69e98915 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I886c2494bdc82c917ee66135ce52c761c347c8fe42ccd63d769cf315b338f2da);
            I48e0ff7c513e9892c552947f3bb0a96d7b00d0ccfa3d7fbcf067d996b3d58dc6    = Idba8e69c73d0fb1bd1aeff84e1c6d06234801f1b37b84ce20a98d29b69e98915;

            I24f0d7d25ccdb1594c03394c4cfccf9327de3684e2376c8f06e56077931820de = I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c + ~Icd7ce463860bc6f62da8d62b71970658ed2c5d5872a56b8429d9223197ef0ad5 + 1;
            I204e9aa975645dee8af1ae12716c4c3a3a6f3884a24fcb113308d16a718f5f74 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I24f0d7d25ccdb1594c03394c4cfccf9327de3684e2376c8f06e56077931820de);
            I904078f4d964b6f66502423cb801a285f9cf21964df0a9fc1b8fdb9e35090265    = I204e9aa975645dee8af1ae12716c4c3a3a6f3884a24fcb113308d16a718f5f74;

            Ibedce4b737f7d1af34a1abb100d92a4a680c939dfc6cc74ea55aaf139e0b9bf0 = I40e83b140f2431f6ecef22d0c8d3ce94b39fac706b8c2a1ed57aa0809900d35c + ~I83b2a186b150fb7290623bd1cbab9d044e9b5c760ed36ae218fb775354e46fd2 + 1;
            I21423b347d172e9152d4a76123a9fb34cceae15bb211e99de5a3f25dd54b3d92 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibedce4b737f7d1af34a1abb100d92a4a680c939dfc6cc74ea55aaf139e0b9bf0);
            Iaed17e55ab4220ad1c1485ce0b5e5518cfc682531407f36561bfff3ed5026ff6    = I21423b347d172e9152d4a76123a9fb34cceae15bb211e99de5a3f25dd54b3d92;

            I217ef743b51672b0333da788f3206b6ca50dd43195a27a9d1aa1b542b7f3c77b = If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 + ~I0442e99f7519b58fb576a898b41563a174beef69bb6a525712224f5d767a5867 + 1;
            I5c1ab87b7496ac411fe34c8295734d2eb6e3dce0c3770f06c2e61f1e9817f3e0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I217ef743b51672b0333da788f3206b6ca50dd43195a27a9d1aa1b542b7f3c77b);
            I101c35283ea20516f74f90cdf4ea7f1ac3a008d80dcb4b80235a17483b1f5211    = I5c1ab87b7496ac411fe34c8295734d2eb6e3dce0c3770f06c2e61f1e9817f3e0;

            I8863222d9076063d0d2c673dfc8fa35d8fdb87a6b37ef7f98988e5c780d556e1 = If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 + ~I698aa30e42ad4f250363d29dfc5117677b19f2da0afa75a013718ac5b9731d6e + 1;
            Ia0a6c602c6591f708fc304b12d671520ec5327d8e45f7f066d24195464f454f0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8863222d9076063d0d2c673dfc8fa35d8fdb87a6b37ef7f98988e5c780d556e1);
            I1184b619aa3fb52506bcb002a57a421ae2f9d3a85502d2ae8132f38092c38fb5    = Ia0a6c602c6591f708fc304b12d671520ec5327d8e45f7f066d24195464f454f0;

            I1a45983bc2d6c4bb8453ee08cc254497e08c85ca326de079180eda79e4a64b55 = If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 + ~Ie81fcb1c1ed576d911918860ec73a2b7823bb2d435a0477ef407393052729326 + 1;
            Ia440e9ed203fb96d0b71bec0c8c3f8aa3ae0cceba15ab536fb4704dcb62e27e4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1a45983bc2d6c4bb8453ee08cc254497e08c85ca326de079180eda79e4a64b55);
            I08fc2b9a844e2c482e2bf89714e92b5baa0ff2b9bc456c523d6360e5b5bbe2d0    = Ia440e9ed203fb96d0b71bec0c8c3f8aa3ae0cceba15ab536fb4704dcb62e27e4;

            I6e02998651462a264077c956dce9fffe5b787e53970bb3c192ab8ca4041e7ad9 = If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 + ~Iba39b0599ed448a7fdb07f6042ef972612b54c7251b256373b30788f64f616e6 + 1;
            I7f640efd56c0cd13cd6a2f7cebd9483076cc85b4668036f2739503dea91bea34 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6e02998651462a264077c956dce9fffe5b787e53970bb3c192ab8ca4041e7ad9);
            I5617f2c448f426aa20d4dc124625b298648c40b73307feddaa9806bf571a71f4    = I7f640efd56c0cd13cd6a2f7cebd9483076cc85b4668036f2739503dea91bea34;

            I72195f5a2c9e92ab9f5534742a45619c0c1840ca7e3955e24b7af70807d5a4b6 = If70840317a05550d95d44a56f59c64c1d42a90f0c170b9457e6268db9f5cbc29 + ~I507512179a289ecb7d9ddf5e853bb42798df8129655c06e568e0a4a1d880ef71 + 1;
            If34c9fd9dd42116ff47c3db0a0a293a36fc2af3d8b66c4342c75e3c98bc969e9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I72195f5a2c9e92ab9f5534742a45619c0c1840ca7e3955e24b7af70807d5a4b6);
            Ic9219b1b4792455d5f1c104798cfb3ace66806e030172b83b652747280a3ea8f    = If34c9fd9dd42116ff47c3db0a0a293a36fc2af3d8b66c4342c75e3c98bc969e9;

            I1cf05db080e64680bb79c5be7fb32bf5c038ff3ab7396d893b90914ad5472bf9 = If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 + ~I697a55c4cb2dd56ce91465bb6750d05200607607d7eaa0b27accbf7f20ba97c4 + 1;
            If5076cad6c2fedcd5c8e31e38043edbf8800ece300917426b42b72eb475bce88 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1cf05db080e64680bb79c5be7fb32bf5c038ff3ab7396d893b90914ad5472bf9);
            Ia1e3983b6aaba9149d835f0e79d761b34c608f894259979b9e02f9891b0e04be    = If5076cad6c2fedcd5c8e31e38043edbf8800ece300917426b42b72eb475bce88;

            I5249daa78d99d33112b5384478d38b33a088d48e042e4b0820c40fd027c0223f = If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 + ~I4d316d60bd6537dcf09dd9b7eecd93c86af11ddecc1ee65e4b9d65c136527e0d + 1;
            I5c344f207e2150409498a524af2c7238e06c755329a5f2bdc5c298c2ad34d4cf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5249daa78d99d33112b5384478d38b33a088d48e042e4b0820c40fd027c0223f);
            Ibd87e183657088945b5a8789b001bbe566368ecbc0a773fb784a3d26cb6886e1    = I5c344f207e2150409498a524af2c7238e06c755329a5f2bdc5c298c2ad34d4cf;

            I7f768fb70d35694f0691521b3989c85e7ce64041868b4f611ce7020ca3bbc1d4 = If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 + ~I0162ff342347e70b1361d5f3ea70c6f872d9b95ede7f80a0a18a69c84b5ebc8a + 1;
            I85328b4628dee41ae779fa1ca104a03dfdf089ad3ea8d7eede9a0869b1ddac71 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7f768fb70d35694f0691521b3989c85e7ce64041868b4f611ce7020ca3bbc1d4);
            Ic67c3bded52308b7875b1fe59eac4e253898565ad36a0f3cb39051d5a1a0289d    = I85328b4628dee41ae779fa1ca104a03dfdf089ad3ea8d7eede9a0869b1ddac71;

            I0dcfa4dc673b57614cd3760b4c618e128809db705602e53f5bdc6f6030b54a50 = If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 + ~I47d2361b09dd6690b6b0a7827348e9e420d8b97c4b620a4e4928c8cbd84c321b + 1;
            I9d0a71f3a423efa567a3a55121fb24edaab598e2f36e51d7d2375c99e0554472 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0dcfa4dc673b57614cd3760b4c618e128809db705602e53f5bdc6f6030b54a50);
            I496a0976329e8a4f6d29dbe1b1e9319f3f99afc9f4d3c645f264f4675b7ebf7b    = I9d0a71f3a423efa567a3a55121fb24edaab598e2f36e51d7d2375c99e0554472;

            I64ae510b10cfc41dc62dc76faa1932a4f159c6e2f4b1aa5e618bec62a190315d = If03c67e8b3cd9a2d215f2dece7fba0d102875369ac16b92af568545b2ee2c5c5 + ~I6182a01d42a30ec5e8883e7d4f5d8f1d657f78052fa4c8ca2c160aecffda456c + 1;
            I830837e25b025c27a2e2957d7d0e12ac498d8eebb18bdea627b46c57ea61bf2d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I64ae510b10cfc41dc62dc76faa1932a4f159c6e2f4b1aa5e618bec62a190315d);
            I93889e1f0f60b124844920662add026c1da1fa6650f347a6a616da18e8b96c02    = I830837e25b025c27a2e2957d7d0e12ac498d8eebb18bdea627b46c57ea61bf2d;

            I9cd6f2580a6f194817cbe4874192fab4f22fc58228a6deaafad44e14f2c27311 = If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a + ~I7355df30b826dd16e0f1fe3be878df80c2ca672dfd1392e2a81ac34fa3df69ab + 1;
            I802acbe8cfa680520493b84328e86b0cc0f5834df73ee11b2b35ed9997890e77 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9cd6f2580a6f194817cbe4874192fab4f22fc58228a6deaafad44e14f2c27311);
            I9bea46de6ec248c77242ae2154d5c6e1dc17ff892dc903bd685badcbaf62291e    = I802acbe8cfa680520493b84328e86b0cc0f5834df73ee11b2b35ed9997890e77;

            Ie5f920e3e83787bd026f94181b522cf7f247cc0863da71e59f8291dcc4c43de6 = If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a + ~I4eb359966514f007fea3e135207ab27fc596987f985b8a3ec6bf51dde2ff9e38 + 1;
            Ib29fb4c64cf1af8604b28c3cc158c13665bc570089df0e6ece0139f858aeada1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie5f920e3e83787bd026f94181b522cf7f247cc0863da71e59f8291dcc4c43de6);
            I88a966d14bd155320f8f49d164cf93516a3822b9098c6417bcdb8a64f9eb1a38    = Ib29fb4c64cf1af8604b28c3cc158c13665bc570089df0e6ece0139f858aeada1;

            I8eed9a916e362776814cdab4ead58e68fca91b54a6648993b57e919c07e132f7 = If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a + ~I0cdb70836bdb3237ff43b23b1676a274cc0dfcffb214799b78ea02c2b59049fd + 1;
            If5ee0d8bd36fdba065830db60c4511892d5e360e74ad676ce84ac82ba47d3e6f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8eed9a916e362776814cdab4ead58e68fca91b54a6648993b57e919c07e132f7);
            I23c475c49d2504d72c81fcf2a1ca3122e6dfbc9f1e9faa0253d0d36c27881126    = If5ee0d8bd36fdba065830db60c4511892d5e360e74ad676ce84ac82ba47d3e6f;

            I859eda2ded7b867c15e420278c996c195f0217d795b6d53acbfc10d218279f02 = If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a + ~I4eb03f5790e18ea72980b8c37b602469d6dba5f850ca3721f49279b4e14cb7c1 + 1;
            I3e2780681adfda07b74c32d8a680f36823f2019a5f63c879113a2b258a339a24 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I859eda2ded7b867c15e420278c996c195f0217d795b6d53acbfc10d218279f02);
            Ib19a40aaae7bc965afa2506ee77fab296894319861766d0f6ede0e69e01ad17a    = I3e2780681adfda07b74c32d8a680f36823f2019a5f63c879113a2b258a339a24;

            Ifa68deabe5c470e4f9f865f60e32710252f5f104571ba859388fd37ff0ef320c = If0deb5dc2afeaf739060bf86beac8013dd92983765107d8cb4460ac86727632a + ~Id645d98c8a2ba63ba9060280b1810d0ab7120f007f3f174e1a501a1f487190a0 + 1;
            I90657433c04f6300a3caf3c7aa1ea345ff62a9a5fd422d7326fe435a0236cb48 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifa68deabe5c470e4f9f865f60e32710252f5f104571ba859388fd37ff0ef320c);
            Ie10eac9c8e0f2526d443d3c8d9c007e29481ae4fd9bed2afac5a0861f80705c0    = I90657433c04f6300a3caf3c7aa1ea345ff62a9a5fd422d7326fe435a0236cb48;

            I1848915027beaf897f1fede8fb30fe33c1f7e5a565022bcae733a9462c9c8447 = If15a6d2660b407d89dda6c113578519092d37491671c47feae8a7a68565a9184 + ~I16ef3abe43350c9096f6c7e597c48fc86ed26a073055b7bcd696c34676529372 + 1;
            I7e6b7e7d088f47fdb77cd0972877c65678f1d1e84f865a4f6a2dc3530ae75e8a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1848915027beaf897f1fede8fb30fe33c1f7e5a565022bcae733a9462c9c8447);
            I873fa9e73fcb148c0eab3dfc8d6163714e0a0dd5889d5d5dd73244c4f700f3bf    = I7e6b7e7d088f47fdb77cd0972877c65678f1d1e84f865a4f6a2dc3530ae75e8a;

            I318c86cd2c86410c5bb1decc6f5df2d544973c518750df70527d2c1fc0b2947a = If15a6d2660b407d89dda6c113578519092d37491671c47feae8a7a68565a9184 + ~I034d52d03f918c91bfc6236c72b0d40b688e2bd353f9ca1f03f4c61449bf128d + 1;
            If50d96b50d6b829bdd534f141f7fd453812eab2373e6780f811dc8e43f61c9e8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I318c86cd2c86410c5bb1decc6f5df2d544973c518750df70527d2c1fc0b2947a);
            I2d891a9027bcd15bb7deaddca0e282e872204770ad4e90ffcd4826beb3c492cf    = If50d96b50d6b829bdd534f141f7fd453812eab2373e6780f811dc8e43f61c9e8;

            Id69048c2098191e826ad522a678bc79cf72544621a8d1d2ce28f0c5797251fbb = If15a6d2660b407d89dda6c113578519092d37491671c47feae8a7a68565a9184 + ~I6822880688515ff8108fe78fadc5d22b953ce5face9928836f824aad9355a713 + 1;
            I80f0dd7462a99f7863728dc9f513999e8df4d944672470fb4f614f0ab36b1bd7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id69048c2098191e826ad522a678bc79cf72544621a8d1d2ce28f0c5797251fbb);
            Ieae87e6a29536e19a2589665b2af980e34700c9a614fe1b7c4704a7a538a8f8c    = I80f0dd7462a99f7863728dc9f513999e8df4d944672470fb4f614f0ab36b1bd7;

            I54fb2b89dce635f5e04010aa85747b0fc135cbc6f58f5b1a92414b2b82fa9e3b = Ibc0fdfece0d7aab4a85b2874a047e1bd390aa826df0d979166e8721339410c39 + ~I3088ff7517eebe83fe5804308d22b8c6190077f576f2e680848092e21116b94a + 1;
            I9ad57caee3254be43c193b522b06af8f1b0603259b4c61f9db942f7d21afdb19 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I54fb2b89dce635f5e04010aa85747b0fc135cbc6f58f5b1a92414b2b82fa9e3b);
            Ia30f6d6396acef716d7383513ac1f4caface96330dcacfdc5302bbb0408697cb    = I9ad57caee3254be43c193b522b06af8f1b0603259b4c61f9db942f7d21afdb19;

            Ifdde108a572ae924a2890624cb24fd7f4beb70c6c8942886fceac443de8633ae = Ibc0fdfece0d7aab4a85b2874a047e1bd390aa826df0d979166e8721339410c39 + ~I00e08c73bb2036cde2d53598b9977dd2504934b9ba8b58bfccdd21adc2fd223f + 1;
            I97a181e9f8555a1bf3d9e9e1876e0ce599fa7c1fff5d905fdd14787e5b92956a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifdde108a572ae924a2890624cb24fd7f4beb70c6c8942886fceac443de8633ae);
            I794ed9d1df776d692b623e89b6d6ade5d265c9869957ddd8e256061bb513d7ea    = I97a181e9f8555a1bf3d9e9e1876e0ce599fa7c1fff5d905fdd14787e5b92956a;

            I0af9db61e66fad28ef275cd396214b69dd646a4b79c44e1673c4ad61458d98b3 = Ibc0fdfece0d7aab4a85b2874a047e1bd390aa826df0d979166e8721339410c39 + ~I694ec7b5bec025b308c4cb56eefedc2be0842202dfb047b5a94dc749c757bdde + 1;
            Ie9fe82e8e7d32f0c47e6b0f9514a270018114d60c63841f864daed7f586a1732 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0af9db61e66fad28ef275cd396214b69dd646a4b79c44e1673c4ad61458d98b3);
            Iaaffc28ce6e25495dfad668af2f560c988f5a5abb76db94b71563231400c28b1    = Ie9fe82e8e7d32f0c47e6b0f9514a270018114d60c63841f864daed7f586a1732;

            Ib6c59e6ecf314597ab396dbceb18037c0d32f40a9022055628288855ec99fe95 = I09301323ed69c3f202b9693f2db743880d6e7618dd91405aaef90c34e61d1caf + ~I830406b0cd2e64515811ab932e9ce01d413f0a68ab7939a2fa14e4eee7d04a5b + 1;
            I28db4525c76b4ffd978720f47196c17b188839e095de0fce72cfaca9754cf2ca = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib6c59e6ecf314597ab396dbceb18037c0d32f40a9022055628288855ec99fe95);
            I45324df36dd601c219634e39418995a9ab1bd58be03cb5dee89ac2d01bec1dde    = I28db4525c76b4ffd978720f47196c17b188839e095de0fce72cfaca9754cf2ca;

            I1eea8e0dc933632ff46ad76cc672689ea6fb253ee0c6168d915353d14fef838b = I09301323ed69c3f202b9693f2db743880d6e7618dd91405aaef90c34e61d1caf + ~I3adad3708bb709ccb06c77ab54c92b6c6629853f740147fd958e6200aeee81bf + 1;
            I41ad0bce74c3d43c94ef9f055ff34fbcfadc63b49f45c24e3480735e706842be = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1eea8e0dc933632ff46ad76cc672689ea6fb253ee0c6168d915353d14fef838b);
            Idc26ae0a7d9ab347f3c75ed2ac7c48f6937f9cc035d46be065fb4b15699cc989    = I41ad0bce74c3d43c94ef9f055ff34fbcfadc63b49f45c24e3480735e706842be;

            I6bd5ddd44f3524fc7691c1957820f067009d145a484faf5edd0d2e527836e12a = I09301323ed69c3f202b9693f2db743880d6e7618dd91405aaef90c34e61d1caf + ~I99a4bc7f129030d12eeef0507cf52503af3df70717d1ba9c38b5dd3a5ffcb616 + 1;
            Ied3eba558946ec39b989955200539b5593fddf4102f7811dbdc1fa0ee35d94d5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6bd5ddd44f3524fc7691c1957820f067009d145a484faf5edd0d2e527836e12a);
            I8e22237e0bc0b24825cc53a9b88f0ad973a825d25aee1abcfddcbb6ddc14ea48    = Ied3eba558946ec39b989955200539b5593fddf4102f7811dbdc1fa0ee35d94d5;

            I193b91d093965a3b2d7ce6cf215348724929cc0c1a3851f9885f822cbcf9ccc6 = Icb4397b9bafcf2461e592a0050cf42f2832d3497c940f82fbe98e855a1153129 + ~I08384d6ff32b692ca710ac4170d45cb5d2e2df509bbc473af140dc50f51fe46f + 1;
            I0a0b709e36be096f2b7a9882b1de9c86a46b08e7693be36bd4e70082d5a7e1a7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I193b91d093965a3b2d7ce6cf215348724929cc0c1a3851f9885f822cbcf9ccc6);
            Ieff55ba27500b6d175abdc30224d7d4c703ff1ce6a3b5d86475b739903839b52    = I0a0b709e36be096f2b7a9882b1de9c86a46b08e7693be36bd4e70082d5a7e1a7;

            Ib31c2929d1523de377924c1f54c6a251313afcbd3c1958aa3e9c0e097c391485 = Icb4397b9bafcf2461e592a0050cf42f2832d3497c940f82fbe98e855a1153129 + ~I8a3c94278b7c901702cf1b70e89c1832afee395077555d27badd4e2b6fde0b7a + 1;
            I788b4acf11f5bbb2ad13fb9d931f593b149f2e9c252773e5044d8a9268cc818a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib31c2929d1523de377924c1f54c6a251313afcbd3c1958aa3e9c0e097c391485);
            I79948c8c3800c594e6e33eff537e1b38872775f3674ce78ad963f09de0091486    = I788b4acf11f5bbb2ad13fb9d931f593b149f2e9c252773e5044d8a9268cc818a;

            I60d9fc72ce19f1ab5a6385844f0660250ee06d76e80845945bb345754280418a = Icb4397b9bafcf2461e592a0050cf42f2832d3497c940f82fbe98e855a1153129 + ~I668aff5da6360f719a2467c5189f3e53e8eeb310f4c4e26f55f8c39e9dcc4be7 + 1;
            I674adba378ccde904a1bd264c3b6dc3f85faabaa01831cda8320aab4561fca87 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I60d9fc72ce19f1ab5a6385844f0660250ee06d76e80845945bb345754280418a);
            Icf4362e74e763b339d2ba9634282b8441d0c293aacbc2879f95a53ef1a2122e6    = I674adba378ccde904a1bd264c3b6dc3f85faabaa01831cda8320aab4561fca87;

            Ia5a27c8c5d46b95fc3ca75cf9e499c6cf406d7320e97b8e0daffe069322e6466 = I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae + ~I257c396883faa57c509e7257bed0829f9ca51f30a1004ce730d48e1e5b40c0ff + 1;
            I6039c5bf499421e601aa8290ecfe5a0e32552869e3222d6a881938886ee0e50b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia5a27c8c5d46b95fc3ca75cf9e499c6cf406d7320e97b8e0daffe069322e6466);
            Id6a3fad936fae13ba6503265a6a9a2bd1c54dc3fcb3d196623bf8aad32225687    = I6039c5bf499421e601aa8290ecfe5a0e32552869e3222d6a881938886ee0e50b;

            I9bb7b61602527be7313761f2a4d22ca145be6a35d06702f60aa9c6c05e9e951e = I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae + ~Icf6fe11d7e6948c0bdb9cd50a0135c3b0fac213aef728b8a6555b7601c51cb7e + 1;
            I823e547aea1e595b2a0345fc0866815d5195979bd55744098366f536832a36da = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9bb7b61602527be7313761f2a4d22ca145be6a35d06702f60aa9c6c05e9e951e);
            Ic26999f764390a0c1461876b7687ee02acb7586ae1e24d171988084ca9d4aa82    = I823e547aea1e595b2a0345fc0866815d5195979bd55744098366f536832a36da;

            Ic3229f0918087445c3b245f3b6a66fcf9d241cf8c9b7a22ff7cc3f127bea4dad = I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae + ~I3d284d86f6c46162d3e0f913a5a6b0e1f2e34fc7ced6a0c226d5e78da81a0633 + 1;
            Ie728139df8a2d5d2cab83b4b4be5c462dd69107d1641666f7de5170c7e83d6dd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic3229f0918087445c3b245f3b6a66fcf9d241cf8c9b7a22ff7cc3f127bea4dad);
            Ic77bba83655ba517bc6313df02ee80ace5ba5e383e3794f971225d42bdf82690    = Ie728139df8a2d5d2cab83b4b4be5c462dd69107d1641666f7de5170c7e83d6dd;

            Iac6d1591feda87bfe1caec1ba6e2a272327d77aff99c6f47f8907caad520100f = I60d1d04834bb93883c91b0c12d003aa1fc9959033fe41930fa49b268ea78d5ae + ~I4583579034ed3bcee2ef0ea2b32a4adf0467f78a2770a84da9948e8d366c1f4f + 1;
            I5e202ec46a29f008d78db131cfe4015f74fdf5a888f7dc1a700a94c5c18375c2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iac6d1591feda87bfe1caec1ba6e2a272327d77aff99c6f47f8907caad520100f);
            I01ac098466c350975d0ecff2227564446e39a21fd133aab22628a9cf3a866b90    = I5e202ec46a29f008d78db131cfe4015f74fdf5a888f7dc1a700a94c5c18375c2;

            I389c3b8f8caab2e397e5f1368db3c31b6c9d81578e1c6ff3c77614bb3fa283af = I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e + ~I7ac4d72123feb2b9af1a6c3da5adba445042363194ef471c8761e289178d0253 + 1;
            If8df36cd42c3c76dd956f677770fc7b64fea6708efc711d8010a976ea719331d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I389c3b8f8caab2e397e5f1368db3c31b6c9d81578e1c6ff3c77614bb3fa283af);
            I97389ae6e03b0e2bee0e882909d2adf1aa34eecf73084ceab73088e850c24e87    = If8df36cd42c3c76dd956f677770fc7b64fea6708efc711d8010a976ea719331d;

            I261d8c9755317b6e7d448fed52871b8996ee8b2966c2cd1c0d9c8c4fff09c1ed = I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e + ~I4bed271962970c26ab72de275bea4b2fb0565d7e44f15b2a1df631bba9e5d4e2 + 1;
            I020d4065b6ac016b70540fa3ec5d128c4c095e5b2f0bd807223b03aaeb730aac = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I261d8c9755317b6e7d448fed52871b8996ee8b2966c2cd1c0d9c8c4fff09c1ed);
            I059c355ce17871c1a494b1a39b4ad3408ab5d28b886b143e04c71a29731f4651    = I020d4065b6ac016b70540fa3ec5d128c4c095e5b2f0bd807223b03aaeb730aac;

            I8802f7a26c9a45d00b3c92f9d62988533adc832b43fc024798ead3130d41af9c = I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e + ~I8741cd8af2f9c3a548c5c39709d7a186f0953de5af6d09d88901e0083a539096 + 1;
            Ie79dee20ce2f12658f63bf8f47e8435a7993e0185c8c6a9aaf81a2f7951bc1fc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8802f7a26c9a45d00b3c92f9d62988533adc832b43fc024798ead3130d41af9c);
            Ie5a7256fb2ee0e45b0cc306c46856bd7cc606efccd221b75d515f608ad567603    = Ie79dee20ce2f12658f63bf8f47e8435a7993e0185c8c6a9aaf81a2f7951bc1fc;

            I2955c07f64b9d8ca9a7a1ea0ff4fcc472588cf5046e22d529a9a674e264bec1f = I8aa6a5fa70a6421907e19d21a85f31542fc4e33178c2d9f05e71e2edfd501a8e + ~I86729a880fe730068d538da490087a1ab6789327f964722c9c14bd9b1c2af35b + 1;
            If8c5f6c0f6af8b9c18c00ab1116cb2cf9a93ec2f992be305dc553a7e858fca87 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2955c07f64b9d8ca9a7a1ea0ff4fcc472588cf5046e22d529a9a674e264bec1f);
            Ib419bb101d14a1958ca5b3a7c6a72d8fc15ca6e217fcac0f7eb84c776f3b0826    = If8c5f6c0f6af8b9c18c00ab1116cb2cf9a93ec2f992be305dc553a7e858fca87;

            I8e2591213eddf0e31054520ebf62ecfa31656b0b4d8cc948e2f0ad6705f72967 = I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f + ~I54b0290e037c2111cfef49e6b33d9a3fbe3e85f8fa8a5c707832cb5477f5c0f1 + 1;
            I7036a280bf3fb8f4d5ce054b2a19cc759ebf28fbfbeed38e6885b95899e1e4a9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8e2591213eddf0e31054520ebf62ecfa31656b0b4d8cc948e2f0ad6705f72967);
            Ie5a479b36bb003e0b2d92a68e955c1906c3969ee52a96b4aef5a84bc275f3f9f    = I7036a280bf3fb8f4d5ce054b2a19cc759ebf28fbfbeed38e6885b95899e1e4a9;

            I3ee55f4d76c10bda1e1ff4074e72e0c0e51486a3659df6c99998dd58f48ac2cf = I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f + ~I2785beda1166504e0b7ea979dbf6c2c5574159cfe36c60fced2dc64ebd05a9bb + 1;
            Ifa80df411d8316c4d2acf8c1a094ba67ae97da2e64e440745984aff2f7a6061b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3ee55f4d76c10bda1e1ff4074e72e0c0e51486a3659df6c99998dd58f48ac2cf);
            I380a702cee9dcf67af75101568b0a417c567c5ebc9e777dd1fd2d297c2455e90    = Ifa80df411d8316c4d2acf8c1a094ba67ae97da2e64e440745984aff2f7a6061b;

            Iaf6b2159a554a3e4e02eed8fac29e769a0ed0b4023fc888e72167c90055b82bc = I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f + ~Ibc54f1c4736e5a4608208441ce8d81831a0b6c7448083d6e6976981f8a38d1c9 + 1;
            I4d5d4c0a9031c2d7b9be5be76b42d25709e833098352ba533ad05dcb34571942 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaf6b2159a554a3e4e02eed8fac29e769a0ed0b4023fc888e72167c90055b82bc);
            I44aed07314ea5c6ed70e468558116a9b956c9a2d67e52229ac85b62c1b511d36    = I4d5d4c0a9031c2d7b9be5be76b42d25709e833098352ba533ad05dcb34571942;

            Ia11f0a7c148064962721b3b128e05210fab5edf48970dd483ba21c75d7076ae0 = I348e6ae792184b176d2eae27d1e7532a8be7d4733052a4c63990725045ebf55f + ~I0f8046b4f96acee2bfb4719bbff91b4b1b81c78ac36ec6e95008a3d9cb5ea6ff + 1;
            Iaeb27fc85e957ef3ea1cdd8db5ebfb513394c5f1680bd98e53b09552b554f80f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia11f0a7c148064962721b3b128e05210fab5edf48970dd483ba21c75d7076ae0);
            I7f63700c8702ba858d076a1901ee015cd80dd29b33e109b7ce64aa14493461af    = Iaeb27fc85e957ef3ea1cdd8db5ebfb513394c5f1680bd98e53b09552b554f80f;

            Ibcd8c95e386f314abf1373ef45a9e95ce079f6eeaea2beeed3118823f184bfe7 = I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce + ~Ic0fd25473d5639721dddea090dc037e39e4a0c08776c0a343408dfcfc402fa99 + 1;
            Ia109c552edbb715f4515acb56e6ce5edbc0bd73fe58165ed7cce5a35867f6332 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibcd8c95e386f314abf1373ef45a9e95ce079f6eeaea2beeed3118823f184bfe7);
            If8bbc0d7554b094c7dbd8b4a06c4ef791cd6e66621e4c3b97464052276957603    = Ia109c552edbb715f4515acb56e6ce5edbc0bd73fe58165ed7cce5a35867f6332;

            I8cde7e5629b3ca36c06d61c7836e7944e7fe1f12ee5bb6722ba97f125eaa5d54 = I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce + ~I8f671fbd5e9e240cc2f3a9c60c1340fb4bea46c25cda7ea5e42c7ca0c2360bb5 + 1;
            Ie22b4331ce03a83f7b77b0ae01cf869497d506d764f6295831de5522518bfffb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8cde7e5629b3ca36c06d61c7836e7944e7fe1f12ee5bb6722ba97f125eaa5d54);
            Ib65f0444b24cc43c4ebe5dc5fb7a2e0aad7c8d125bf92c527ba5dabd52d8f98a    = Ie22b4331ce03a83f7b77b0ae01cf869497d506d764f6295831de5522518bfffb;

            I9f8966a82409d3b30ee1cd52c7e0b4976cd317c1ec6bfd7c6c23e4157a556d9f = I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce + ~I4b9dd5299690e88d870ceb4939b7f8fdffc8419431458851a3691de4f78f9f15 + 1;
            Icd8816eeae15f7d5422c702821ce9d5fe0e272f5165cd7c6f100156f9cccca72 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9f8966a82409d3b30ee1cd52c7e0b4976cd317c1ec6bfd7c6c23e4157a556d9f);
            I088890dd5f7391be17333396dc9b8cba40ddef39e657378c312707e1ea43bb56    = Icd8816eeae15f7d5422c702821ce9d5fe0e272f5165cd7c6f100156f9cccca72;

            Id1cb12cdb0a13b705c9450d25160d92c2ce8624a1fdd447cc4db14c29512be59 = I77864bcb0c57c3e10a88e4c97b91d33264cbc3a2a9722a64ec548355f70a3cce + ~If08c85e70828c39162bc16d65747d3d3d0a6176e8db106b262bbadd651f745b7 + 1;
            Id2f34f393c20f24e86ee88f74da7085cae9c4df6d25b805f32adb16cb2bfc69b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id1cb12cdb0a13b705c9450d25160d92c2ce8624a1fdd447cc4db14c29512be59);
            I64fcddc23b1b1d72f4a5cd8707f8ec3dfb77bd105d279d01a99750b9ec4894d6    = Id2f34f393c20f24e86ee88f74da7085cae9c4df6d25b805f32adb16cb2bfc69b;

            I281aff7f22feb2745825babc1e61ce1ee1bcafbbe54bb01b19ff94ac6ad162c3 = If999edef9d50e83e5c53e4715e8f0ae2699c9ad1960e7e16ec5049a8ce0068e8 + ~I113d1ff61779dda7e1209787ba652b8b332fc5811cdc0aae65a304aa89d56766 + 1;
            I541091c82a0e29abaf2bb1c586f5c44501e90f7ac691f250690ff6fc4f186307 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I281aff7f22feb2745825babc1e61ce1ee1bcafbbe54bb01b19ff94ac6ad162c3);
            I323a7ad384b7514bf52fc27d18b29da7effc88c35471be18c85d0b61ece11db3    = I541091c82a0e29abaf2bb1c586f5c44501e90f7ac691f250690ff6fc4f186307;

            I0834faba181b93b43416922703257ebf7f2d35bcd63746ca52c83e57dd801731 = If999edef9d50e83e5c53e4715e8f0ae2699c9ad1960e7e16ec5049a8ce0068e8 + ~Idcb8d71f1ea9d314ae8f26e9f4b9e25ed245bad319b9af2f71b035aca6d8fa6a + 1;
            If809f343f9007d972db4bafabd3a2c1f1a5d8a7a965cc6924aa965005763fcd5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0834faba181b93b43416922703257ebf7f2d35bcd63746ca52c83e57dd801731);
            Iede33454e4e4f5856e3700d92d14d4b4ee573de70aa6715525cb1164348e6561    = If809f343f9007d972db4bafabd3a2c1f1a5d8a7a965cc6924aa965005763fcd5;

            Ia61ae97a6d0793a9e542fbebdea72393e93d4e1cd4bd260432bec83e5503116c = If999edef9d50e83e5c53e4715e8f0ae2699c9ad1960e7e16ec5049a8ce0068e8 + ~Ia0ee127b17b441cc11d664edf15d370368494e31b52c4865c97a065ef8bc43b8 + 1;
            I75b60c610ccc4ecb84b7616f74cf1cc68e4312dec53d71e99911cfc9f69ec69c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia61ae97a6d0793a9e542fbebdea72393e93d4e1cd4bd260432bec83e5503116c);
            I6254bd01448c9d8e8b348c9cf6f62da72b3e66c76cfc692be2250a30039c48db    = I75b60c610ccc4ecb84b7616f74cf1cc68e4312dec53d71e99911cfc9f69ec69c;

            Icede982a125cdcc6a88aab18ffc06e98ca57e02601729b20fdafef5236a03ca4 = I17d1cca0614280eb976be22c9779a9238712e3fd3d27b84bc092911227433180 + ~I6159ddc580c73acd6e2391f4c6cd9989ebaa8947db61972e4fb97f1e12efd17b + 1;
            Ifbb0c6db7e47972ee1ef163f0f3b0e8346b27ad9fe17801df9f1c4f9a79c6ed8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icede982a125cdcc6a88aab18ffc06e98ca57e02601729b20fdafef5236a03ca4);
            Ib50a67b0b1f097d85a05aefb1686e6d51cbbda0406226d20772af68de6e6d139    = Ifbb0c6db7e47972ee1ef163f0f3b0e8346b27ad9fe17801df9f1c4f9a79c6ed8;

            I365aeac8393552a9c42403a734816538b26d9c1429d9dcee2ac6d312fbcd917b = I17d1cca0614280eb976be22c9779a9238712e3fd3d27b84bc092911227433180 + ~Iac102173e8323a836c8f86d266f551fc24ccd14aaf39c7d9ef26c465d38706ac + 1;
            Ied45ebda32de8ab6f352042b494f0350315f9a86a12bcd18991d3dc774876ce0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I365aeac8393552a9c42403a734816538b26d9c1429d9dcee2ac6d312fbcd917b);
            Ib0809c22530a4fef601b75ff7573a7e9606b2da1938ed0918b43a958b9c2ddb9    = Ied45ebda32de8ab6f352042b494f0350315f9a86a12bcd18991d3dc774876ce0;

            Ic7aa7756d5779803ef1deba260ec7a2dfbd59071f84e0e73118751dbd57b2737 = I17d1cca0614280eb976be22c9779a9238712e3fd3d27b84bc092911227433180 + ~I8c494bcba3ff73ff29d9d388708fa34caa73b883730349aef6c2648a2f5a1409 + 1;
            I63bc47a8fa8e183d1451318367b43a76386d269e4ec267b71169127ad5c5a46e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic7aa7756d5779803ef1deba260ec7a2dfbd59071f84e0e73118751dbd57b2737);
            Ia0febef423616e7d4ab3957eea2ba1de8a8bba8b027652658ac2ab5aab11b9bf    = I63bc47a8fa8e183d1451318367b43a76386d269e4ec267b71169127ad5c5a46e;

            Ia771e5a1a22d051469c95101abb12e406a5aa0518905b1c475fd4fa0b7fa520a = I20665258f942651538aba58d63ca7f531a375ce0ad65c83a1aad4cda0815b334 + ~I2f4a0e474435a97fa5d2d056d9de566288c0624cb094d71685934475b58572f1 + 1;
            I6a82ec3534f3eacf85d6fb59ea0a6d640df62089427d83d5a9f494661e44e942 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia771e5a1a22d051469c95101abb12e406a5aa0518905b1c475fd4fa0b7fa520a);
            I8cdc972ad763857aa9a0cf1145ac106bedcf7897da19e06cdac06cbbc52e0141    = I6a82ec3534f3eacf85d6fb59ea0a6d640df62089427d83d5a9f494661e44e942;

            I9af1d3493b4b64704551be835abaf50ac8b247571a802846076fcca1f5f8fc6b = I20665258f942651538aba58d63ca7f531a375ce0ad65c83a1aad4cda0815b334 + ~Ic96ea379edce04b88c524fd17a2b6fb2283e45735640aa3d8ffc7f1bca77c78c + 1;
            I63f3c451c1d8566df035f6ebeccdf248343fabcea08423509f9caab46bb7a75c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9af1d3493b4b64704551be835abaf50ac8b247571a802846076fcca1f5f8fc6b);
            I10d197005aafecec4bf8c18547bda5a551dac520da311ee42db394ac67f413f1    = I63f3c451c1d8566df035f6ebeccdf248343fabcea08423509f9caab46bb7a75c;

            Icc0a08bd18253bf9fad9b320fb7462c70107db49b1c8f67126a9bcf2734f54c2 = I20665258f942651538aba58d63ca7f531a375ce0ad65c83a1aad4cda0815b334 + ~I7ea6f607967e7d251d71b4c4b3dd545a4a9ae8298c3ee2356bbc16ebef06cb2e + 1;
            I955d2b4663596b343e2ceab53a3bb73447741d4f3c8c935f35d72cf9b44249e9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icc0a08bd18253bf9fad9b320fb7462c70107db49b1c8f67126a9bcf2734f54c2);
            Idb166c946a1916a593a1931a1651288e452553572b5b4e272aaa917a4afbc42e    = I955d2b4663596b343e2ceab53a3bb73447741d4f3c8c935f35d72cf9b44249e9;

            I75bb712b6207e8af8c090db486b02880a7c3f82ca47a48929c52e898e36967fc = I5337e70d66d8fb81df05813fd3a172c8337b5d2ca39976efd9dcaeda77844be7 + ~I8de3f6aec12696eef7d069510ff25e6e620fc4fdde5f92923a707116da636284 + 1;
            Ibf7b181b75b6f0fca207af49cfb93611fb71c31c28a5604de13112e8d521d008 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I75bb712b6207e8af8c090db486b02880a7c3f82ca47a48929c52e898e36967fc);
            I3ca7faf1b6e8e04fdab54e1a4b313720f91992013d31b492f9aa49e54676aea4    = Ibf7b181b75b6f0fca207af49cfb93611fb71c31c28a5604de13112e8d521d008;

            I05e3db1dd36c0de58cd3d6d5c692cadb9ac76c905af96474615ac491db900051 = I5337e70d66d8fb81df05813fd3a172c8337b5d2ca39976efd9dcaeda77844be7 + ~I9c0a341c77ecbc1b3c44afee03ccc5a8f34b1275db9c439eedca9ff61a1a1eac + 1;
            Ia6198ea973d8346b504b6da6f2fe193b989253fa47992f709c17ecf344f3572b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I05e3db1dd36c0de58cd3d6d5c692cadb9ac76c905af96474615ac491db900051);
            I77a2d0c0f26725cfe51712e4d1fd8663cdcd4668405e3fabd33e72bf7d008343    = Ia6198ea973d8346b504b6da6f2fe193b989253fa47992f709c17ecf344f3572b;

            I7a6454c2bea6d09f07fe94c2c000ebf70ae11e4552e7e6e2e1d53e09bc529e5e = I5337e70d66d8fb81df05813fd3a172c8337b5d2ca39976efd9dcaeda77844be7 + ~I215148c89dc37a59b3eaf2f38679554281379dc6c8e57718e1c22c091f4d76cf + 1;
            I2dda176f6e7f4c75b5cb93278b95ba9bd30bda61c0d44c103e5092e71d4db7ee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7a6454c2bea6d09f07fe94c2c000ebf70ae11e4552e7e6e2e1d53e09bc529e5e);
            I3c9445224e3dc806a499c5a5faae2cd5691cfb5497852d3aced39ec164d9a5ce    = I2dda176f6e7f4c75b5cb93278b95ba9bd30bda61c0d44c103e5092e71d4db7ee;

            Ibc7f54032db8aeb207641aefc8926732096c74282c740ed04545ea01d1375d62 = I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 + ~I0b60295163435ae3d3b31e9613d753e7e41fd66c11fdf2e7248d7864e11d9d84 + 1;
            I8578eac4c908240f9cd21d004858326a5c6d88ba020a8b0f27955896bd227e30 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibc7f54032db8aeb207641aefc8926732096c74282c740ed04545ea01d1375d62);
            If86de9d134174799b06582013809be1a492e36de3aeae4cab7bdd6a827223976    = I8578eac4c908240f9cd21d004858326a5c6d88ba020a8b0f27955896bd227e30;

            Iaa2a9a1fce1a32dd04ceb055eabc32fe90fc765c2246d2a29f0e847a8ab49f1d = I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 + ~I97a73864c1c919943cec586befbb524fa6d6da6a60e1503bcef8116c646b71a0 + 1;
            I6ce58155e37948ec0a5842ed20258c382c0fd9889e697912d1ee1018a5e25d74 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaa2a9a1fce1a32dd04ceb055eabc32fe90fc765c2246d2a29f0e847a8ab49f1d);
            I6c7e61c506c8d841d4747e5963d49e0237b106ba6cb15a0fc9e4680ccab02c5e    = I6ce58155e37948ec0a5842ed20258c382c0fd9889e697912d1ee1018a5e25d74;

            I3bb50ccd25f72ca813c999533e808c0dfbe3747a6dbe023a303d64e0cd571423 = I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 + ~Ica10d27b8c94c1e740a2287ef28e5d3fedab4221b391b0a3a1da3a472f094039 + 1;
            I13016deb611dec6abdc3b14008afeb343ae5cafa44375dcbb1d09da08c80cdbe = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3bb50ccd25f72ca813c999533e808c0dfbe3747a6dbe023a303d64e0cd571423);
            I9c17caab5e5aed3ddf7a867cf514cdb5f65c3591789f1058a756265f97aabea9    = I13016deb611dec6abdc3b14008afeb343ae5cafa44375dcbb1d09da08c80cdbe;

            I32f852a9a6c5c496bfbecddda78b07f0cff10e6f360c3938827fbe389bbb1d64 = I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 + ~Ibf57f9e63049a49e05739966f1ec2fe4520b2959db6fee3a18ead9ca03aac230 + 1;
            I046da9b39f69a49ca827ae6c66c4164d2c64cb390dc8ccc238a70c68f00e29c4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I32f852a9a6c5c496bfbecddda78b07f0cff10e6f360c3938827fbe389bbb1d64);
            Ic818ff3260f1543c8d940d36c72d644a7a3a243220548792289117ca6a793c02    = I046da9b39f69a49ca827ae6c66c4164d2c64cb390dc8ccc238a70c68f00e29c4;

            I79162ac11cabd67e684b36c8633d4a001a7f794c60468829974f8ad972e9b6d2 = I628613502e3141086348f62966f8db49e3dd9488fd3e65416cee777b52eae0d0 + ~Ief3b5e8fee2d099a90990de9303f34d600235d989d25a30b5a7e2654c18b5c3c + 1;
            Ic7d0c1eb012c5cf07f8df74a28a53ebfb026d43c9161bd7cb0de0fdf8bf6a9cb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I79162ac11cabd67e684b36c8633d4a001a7f794c60468829974f8ad972e9b6d2);
            Ief965ff00c0da0a12a68cadf50622567e99dd688e9bb810dd46f69e3eacb7285    = Ic7d0c1eb012c5cf07f8df74a28a53ebfb026d43c9161bd7cb0de0fdf8bf6a9cb;

            I44868fdadaf261c99a76756dbc2feb061aa5795b84be4aaaaf2b2f14580d85cb = Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 + ~Ie3806d0fc4177d813aade41ad46537a9a335516135161cb2ef18ce822cb301aa + 1;
            I7f53d47b7607b32c4f7401fd9fb07a28d9dee9a3119dbcd0b6f09292a910107b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I44868fdadaf261c99a76756dbc2feb061aa5795b84be4aaaaf2b2f14580d85cb);
            Ib4d1942b7949b0a4e79441e13e3b6b7b36bbb136c2bed6ad1adba30a840f4b55    = I7f53d47b7607b32c4f7401fd9fb07a28d9dee9a3119dbcd0b6f09292a910107b;

            I0e0b35e726d873d7a4d436a763ba90d981031d080d8030d7d1e11907bb246f06 = Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 + ~I211a150dd66153a3c2c72be4c24145e4c9f0b2f9a3032fee9233985ca9d2c4ae + 1;
            I46c1d6509155e8a243b0d4fca0c08cc86e520b8142ff55887efd0b27fc9ec619 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0e0b35e726d873d7a4d436a763ba90d981031d080d8030d7d1e11907bb246f06);
            Idc7991125ae81f1c0d5f221c7fccd90e5aaf92e72e0421aa687e6c1e0f8afa9d    = I46c1d6509155e8a243b0d4fca0c08cc86e520b8142ff55887efd0b27fc9ec619;

            I35bb67b450432187151294ded11a662620636aed3ca3ce1396869fa2b60ed816 = Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 + ~I60f3a2c7d8e3935c04abc8aa09b0a2ef540f13bc98beefc600fd70aa25421191 + 1;
            I8a41819311f3c31efd56be044479263c2afbb88f7c90ebb8ad570237506878b3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I35bb67b450432187151294ded11a662620636aed3ca3ce1396869fa2b60ed816);
            Ic1e2fa322b42a15a886ec6ba9f67656a39c8bd6a13af883081336da43d9d0406    = I8a41819311f3c31efd56be044479263c2afbb88f7c90ebb8ad570237506878b3;

            I90bb979f2ef58854b3b2a7d6b0a574774403e9766c60b1888f1ac97ccf4b9889 = Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 + ~I7cd31013bf73ff7f7aafbf06eba3fe8110dc5490a280c2d79ce53c77896f564f + 1;
            I6c2b8dce255f31b35ddec9776805ae6b3dd2d4d843a755375f49d28a7f7f6d8d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I90bb979f2ef58854b3b2a7d6b0a574774403e9766c60b1888f1ac97ccf4b9889);
            Ibdbd014d7bbe12aa223eaa43939e3459f35b9970ed075d4733932cb66042d281    = I6c2b8dce255f31b35ddec9776805ae6b3dd2d4d843a755375f49d28a7f7f6d8d;

            Ieace5fcde163f3e9bc1be0f05b04d00432343111a05c7195e0999a3cbb3d95d9 = Ic1fcbcc74f9525bf6ef310c35328cb885084c3b442d705030e3d56f3188630c0 + ~Ia2233f4704a9724ec75efe5e31af6807f8f1529f641ec05d053d6a12308f485b + 1;
            Ibe35c53955eeba706ea61cb7d516b391278b1e27ae1eb5f796d45dca20a11928 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ieace5fcde163f3e9bc1be0f05b04d00432343111a05c7195e0999a3cbb3d95d9);
            I4dcdb2c22db70cdfa468f9249fea4262e91120e0d995981b34919e26c9b5bc5b    = Ibe35c53955eeba706ea61cb7d516b391278b1e27ae1eb5f796d45dca20a11928;

            I8dffb8fb698239dca36a5371fe756164e127a33e709084a74d3d2f548edbe1b0 = I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 + ~Idf57b2bf209c68bfc70fe2759595334fabe3d50dcfc4fef8637586c6623c9c29 + 1;
            I4df41d0da488a9cf1999eb318b6654e68637641f78ce9be4636203d6dcab3285 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8dffb8fb698239dca36a5371fe756164e127a33e709084a74d3d2f548edbe1b0);
            I2f6966ba5ca0aea5cb187d9d90bb6b743b80bbc7fc4547396dac13a22603e7d4    = I4df41d0da488a9cf1999eb318b6654e68637641f78ce9be4636203d6dcab3285;

            I7d8b7acb9dfc4a40ecb4156435977770c6a8f6713d612777664eb4c545208943 = I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 + ~I81b8212f2e15845be4d129b192895f659d31a061a3a033bc3ac9ebecc75f73fe + 1;
            I79c3d77c250619b76005964a5d8b3dc5480c395f1b541d7234d846955213a0e0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7d8b7acb9dfc4a40ecb4156435977770c6a8f6713d612777664eb4c545208943);
            Ibec37c7599a7f7cad52a48cb44ea0ffe117ac5ea206590a3eb8a2c661913c9ad    = I79c3d77c250619b76005964a5d8b3dc5480c395f1b541d7234d846955213a0e0;

            Icac43b0373871bc847869a8c5a86a423b2bf8378da0d3f1753a42ac604f5785c = I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 + ~I3af491b2352720f2bd378052706f4ce571453d59b0fc78b3cb0bce2d51ce5700 + 1;
            I0997b7b9813944c111e41c7f375c0925dab34b604959dfdcc8dfcaeb701d6d62 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icac43b0373871bc847869a8c5a86a423b2bf8378da0d3f1753a42ac604f5785c);
            Ieea63392582d451f7570a458bd235afaec2d11a7427d4e706bc1d73128993792    = I0997b7b9813944c111e41c7f375c0925dab34b604959dfdcc8dfcaeb701d6d62;

            I309283aa468ebadbc72fb7bdb48e76697f5222c1e527837ada3ba12084ceda60 = I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 + ~Ic6d228f83da7a1c9a71d8fe70d5adbbab8856e5fd3640d805c4076f5f7d53553 + 1;
            Ie6e358691e81a9c1ca0a585b69352779f083e4f3e26d03152194b1a9238f0f0b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I309283aa468ebadbc72fb7bdb48e76697f5222c1e527837ada3ba12084ceda60);
            I2fc14612ec75b59c28fa90d7a5bfd1bce6d5d1fe0c46ba45f77ee2f9aa9e481a    = Ie6e358691e81a9c1ca0a585b69352779f083e4f3e26d03152194b1a9238f0f0b;

            I055caf108b4457e691ec20569b48a56478f8b0cbb9211271c3a7cb2836605749 = I4ea96ffa1be73b4159bc9e7d00fa716e32d244c87d3ba58e3e504313c7794093 + ~I6754b9c9cc470509e67ba88c2669e1f70666489af9ca14de9fd4e4328d18e245 + 1;
            Ie3480800eed0a0bdd9a7131caf3ce773b28d952484926c279b3a5e6244925a6d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I055caf108b4457e691ec20569b48a56478f8b0cbb9211271c3a7cb2836605749);
            I876dccf88204e4113c5f80bdf348624dfbd5a1439638577670da4c6afe1d5f70    = Ie3480800eed0a0bdd9a7131caf3ce773b28d952484926c279b3a5e6244925a6d;

            Id0bf924bbc09ce9d0e83a26d569bca939f3bd410a63fa3b1ad631798a9171102 = I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 + ~Iaf95e616f53a061a7bf59bf1128d2cf6a5ef64d24b292671a3124a6e010d964c + 1;
            I1ddb5092da74c5ef9553f80099ceb2798e717d25b24053400181825ba303c5da = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id0bf924bbc09ce9d0e83a26d569bca939f3bd410a63fa3b1ad631798a9171102);
            If0c1eced668b91b966c13a44ef09ca1209f96723c7e3d030a757d45d0b61141f    = I1ddb5092da74c5ef9553f80099ceb2798e717d25b24053400181825ba303c5da;

            I3896b59b701e291956a090ff59ca6867a6267fb825629de82c88309ade2dc8a8 = I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 + ~Ib07af5e0c881985b1aa0698382702f78d3ec7ac69cd0deae7496bc63e519a738 + 1;
            I552b1b2def8af8685711597e1db1da516b0766591b757ea9f33c666f9e243ff8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3896b59b701e291956a090ff59ca6867a6267fb825629de82c88309ade2dc8a8);
            I5f3fc42a6dc35a49dba82814b80238d6a9f6e9c8cfddd4d72749a3197115b969    = I552b1b2def8af8685711597e1db1da516b0766591b757ea9f33c666f9e243ff8;

            I1112f35be1ed8725b875aec8350b0843ebff9231fd3d3a49914003c23192822b = I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 + ~I144fae9c9898630fa027b3237ed3434c76965eef2eb015effa7c8677b19c91a3 + 1;
            Ia5703a4566bd7f99d071749104ecbd4712bda3f156cec8a1c4d4d40303e37fc2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1112f35be1ed8725b875aec8350b0843ebff9231fd3d3a49914003c23192822b);
            I677e11f6dcc443a45cc24e28c955adce7dc006e6b26e0ade792740c59d91ed6d    = Ia5703a4566bd7f99d071749104ecbd4712bda3f156cec8a1c4d4d40303e37fc2;

            Ic953289eb284e6e85659eff600c7b373dfd72773441baab0ae1ac4585370d79d = I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 + ~I5b480e9176a1bb70ebc65f73af78889d266a8efa7414cb97cc5255a5ca5f01ec + 1;
            Id5f32d64dc52d3fa4da97ed5a432d520af0cbc1e4714d57788e668a7bf3fb310 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic953289eb284e6e85659eff600c7b373dfd72773441baab0ae1ac4585370d79d);
            I703d9bd8f5b9435c814d93ae7e2327a45e0febce37b67b770c2b93f30ba39972    = Id5f32d64dc52d3fa4da97ed5a432d520af0cbc1e4714d57788e668a7bf3fb310;

            If07db5ea1a4431d5d3e3040559bf352e46983992fe80c37e84468e7f798caacf = I7f4752e40cd4b568e4e457afb93fff14604c53c76de129cbeac0542b65e3a781 + ~I133d5432ba2f64f1ad612b2505fb95ce91962b6ac761dcd0e92f75d1b663d7b6 + 1;
            I9977445235192d6416fdf5221fac29c4586af4f83efa91e128a0cc18cf648281 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If07db5ea1a4431d5d3e3040559bf352e46983992fe80c37e84468e7f798caacf);
            I4d518a62a0a46b493ab538e6ccaec00b9b2cd08aba9695482997b884ae7b006e    = I9977445235192d6416fdf5221fac29c4586af4f83efa91e128a0cc18cf648281;

            Id66a032ba386ed0856ac30d1393b9bcbdd32f34a514b18903c95fc66b287c7e0 = I7214b0ea3f1135ee6e703c8e873696254a514ff1e88c32d42757c8ed40a5b907 + ~Idaa2e762bb01a89e36234967b22cc76cf290937df9295939bb4c4ad08cb8413f + 1;
            I5fbd149fabfe16474e75301b3ec4e0ecf4c70537882f00d8c8fc630e7656b368 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id66a032ba386ed0856ac30d1393b9bcbdd32f34a514b18903c95fc66b287c7e0);
            I67fa42eadbdacb43b464b7246fbecac6c261d3cc37d501efdc1e83b9b1ff6055    = I5fbd149fabfe16474e75301b3ec4e0ecf4c70537882f00d8c8fc630e7656b368;

            I41dadde0137c88dc8b0e9d86734803a46461074a08c6f61e73c8cce898ce64c3 = I7214b0ea3f1135ee6e703c8e873696254a514ff1e88c32d42757c8ed40a5b907 + ~If4c7abf17850a5fcd64bb4ebaef1dc806938542a3bb2b9eee643fdfcfeec23b8 + 1;
            Iceb61d5ca2b0e3fa972b66d7215d7e24047180d638846c80cba9b4e84e147d49 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I41dadde0137c88dc8b0e9d86734803a46461074a08c6f61e73c8cce898ce64c3);
            Idb5ffff327b8edefda5ee44436f5f31deac21a01781b65e2429b1e1a025c997c    = Iceb61d5ca2b0e3fa972b66d7215d7e24047180d638846c80cba9b4e84e147d49;

            I55543ecec7c46f5fae535eca894545a441edeebb10f1b2bfef7c7fae234cedd9 = I7214b0ea3f1135ee6e703c8e873696254a514ff1e88c32d42757c8ed40a5b907 + ~Ifb664074b1a8bb954cb940a11ae4e7de1278edf3614b861ccd83dfaef95319c2 + 1;
            Iac3ec84d526a71f93a304493831b4f9597b2ba176aea1b62dce09eebb9dd0e4f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I55543ecec7c46f5fae535eca894545a441edeebb10f1b2bfef7c7fae234cedd9);
            I0384038afb05788ee28f773a244ec49cd78da115f5d864f8497df2b36f37ae54    = Iac3ec84d526a71f93a304493831b4f9597b2ba176aea1b62dce09eebb9dd0e4f;

            If7778495e794f7ec0ace1408db22f95ed302e9f124858dd6e119eb3c91520821 = Ib9f05dc23ded7e25eec5344da5ea617060c2cb525c22aff7dfc41f86026b864c + ~I7addf7487638274202ddfd183ba052556f89f82da9e873224c5dddf27d2d5a66 + 1;
            Ib6afefc545bb77d065a44983762a6b83fafb326b323fec8946ac2f7b11865d26 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If7778495e794f7ec0ace1408db22f95ed302e9f124858dd6e119eb3c91520821);
            Ibee29fffd6b844b0fc4666fbb35c295ccc5a7b99dbedce125b370508cf6b0b90    = Ib6afefc545bb77d065a44983762a6b83fafb326b323fec8946ac2f7b11865d26;

            I047343beda3ba4373e81c19c51ea3ccd5320a6ba2a595860f87ea9e041afbece = Ib9f05dc23ded7e25eec5344da5ea617060c2cb525c22aff7dfc41f86026b864c + ~I8952c026089661f4ddd0720f6ab16e46334fc934e6775e7163aad8cf5dec6b68 + 1;
            I9781f084a762fe71955603c76c6d57791f2a642ab73c8393d5ed79b42dca7b66 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I047343beda3ba4373e81c19c51ea3ccd5320a6ba2a595860f87ea9e041afbece);
            Ia8f9f47f8cf0ac244089271b1cb952cac9d90aa94b91eef48733afbbcd992952    = I9781f084a762fe71955603c76c6d57791f2a642ab73c8393d5ed79b42dca7b66;

            I9138132d9e54b759171955a69beb971d2b73d6cef41137e9219277fd7627d6da = Ib9f05dc23ded7e25eec5344da5ea617060c2cb525c22aff7dfc41f86026b864c + ~I76ca3c17438c05fc53f6f7075ff7404c0838f62472ffebd41a61afb1f3ea5dbe + 1;
            Iff4386a737586e5cd21336fe2f577e54c5c8bebdca0c7fb944923f8a9ef09d2e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9138132d9e54b759171955a69beb971d2b73d6cef41137e9219277fd7627d6da);
            Ie80058ecf96cf544095e34ccc9662fb679b8da3cf6f10797805cbcaddfd63804    = Iff4386a737586e5cd21336fe2f577e54c5c8bebdca0c7fb944923f8a9ef09d2e;

            I5a11b582e017795d316b18512d5f7809300e13a89ee878deccdc3e4ee9556e3d = I4d36f91f636848b5418807d5da024cbeb73a4b63a9b55c2b9bf48f22f2196857 + ~I7925970ac367f8374fe02f6e4c8c339c58808928696f0acaf85d96fb3f202f00 + 1;
            I1ebcad455793356bccaa94bc33207b868ed70c398881b3ff78c8eab610605708 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5a11b582e017795d316b18512d5f7809300e13a89ee878deccdc3e4ee9556e3d);
            I680b7384eb5b44faf98980956603d7db164a819fe394beff4e94872edcbece0b    = I1ebcad455793356bccaa94bc33207b868ed70c398881b3ff78c8eab610605708;

            I0f690c5588c55c55f7e38c94b4b0678f65ea3214eb2b3923e6888f15ad2e632a = I4d36f91f636848b5418807d5da024cbeb73a4b63a9b55c2b9bf48f22f2196857 + ~I58db55229ca30218227b598184e85d57a0e3a8b61308f8114cd709232573e566 + 1;
            I068c9d5ac9f999a475341bd2e8328de90021df28cbe517e182ad5de16d1a0f51 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0f690c5588c55c55f7e38c94b4b0678f65ea3214eb2b3923e6888f15ad2e632a);
            I7bdb6b57635075a7bb8408a878d4ef7f2ff136804287cfbacddb40bb20dd053a    = I068c9d5ac9f999a475341bd2e8328de90021df28cbe517e182ad5de16d1a0f51;

            I36e15452cc41552f83da26036b7b94a2ad425d1441a3de1d4e226851a8bcb3fa = I4d36f91f636848b5418807d5da024cbeb73a4b63a9b55c2b9bf48f22f2196857 + ~I27ed900fc3d84c4ab4570c3bb88b5e9a7077389e5fa169cc4e1d606f09c9c755 + 1;
            I1524d287bf11b9e8bd9c37a61011f3d9a6d18bc1dc48aa254cf288134bbef748 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I36e15452cc41552f83da26036b7b94a2ad425d1441a3de1d4e226851a8bcb3fa);
            I27f0b66e246c474ca71e1ae20503843b31921b5552092c5ae6eb872e76808395    = I1524d287bf11b9e8bd9c37a61011f3d9a6d18bc1dc48aa254cf288134bbef748;

            Iac99102c92e103b1b841f87f7c024aead79f11f036aff50058281258beecf469 = I55699a1c81182c259ac531c5587702742eb60c998c424e33a62849441a5a94fe + ~I46777db6f6f68d76ef34c4a9c585ac04e8a978663fecf72d2dbaea3287dfea2d + 1;
            I2e88cba4b7ba164003b35e7b7266a2d22b85b731144db715c2675eb9011bf01e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iac99102c92e103b1b841f87f7c024aead79f11f036aff50058281258beecf469);
            Id81f3fed6908e777951bdff6448776a9a80348c44058ba0f9450999a26f6155f    = I2e88cba4b7ba164003b35e7b7266a2d22b85b731144db715c2675eb9011bf01e;

            Ib74288457c278f35939cc8e326fa0db500d368d628b4e60af7921c79991a45d5 = I55699a1c81182c259ac531c5587702742eb60c998c424e33a62849441a5a94fe + ~I6f71faa84bc155810576a85be759d7c06d84dd53b5e2dbc74ab0175e5d64d3fa + 1;
            I18edf674979e3ba4398115ff3e5912b2a41737a1641df1ab7c7539e10cd53785 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib74288457c278f35939cc8e326fa0db500d368d628b4e60af7921c79991a45d5);
            Ie4655a76ed253aad70f2340070cd7b6f2041e6782a87be16ea66ee0fa2e2ad74    = I18edf674979e3ba4398115ff3e5912b2a41737a1641df1ab7c7539e10cd53785;

            Icca50300b717929fbd20809910f35bd0b6fdeb04585be02a41a9aeb2b23e0041 = I55699a1c81182c259ac531c5587702742eb60c998c424e33a62849441a5a94fe + ~I3ef4c55a4a3281a468daa3233ccdbe660c46a930220b5c9bd3caf6041008bdad + 1;
            Ib8387757c67a87e7a37c530022a9539aab577c140512fc5481f00fc9ef52a140 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icca50300b717929fbd20809910f35bd0b6fdeb04585be02a41a9aeb2b23e0041);
            I8acc445f4b9f01af1a8f4f34ab10028472b79a2c1d1d3b8aed7d040f5ff4cff9    = Ib8387757c67a87e7a37c530022a9539aab577c140512fc5481f00fc9ef52a140;

            I0f6953fe9ab3a2018fcdf430ea420ccae2fd35b2acd637cb083370cc86155cc8 = I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f + ~If50a43f14a383995b16d784cc119d01749fd30928019bea1b7aba0039c4c350c + 1;
            I4d2bf12a647b50d4ab9b14ca939986eb9960c3019be93049f9086529acdfee39 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0f6953fe9ab3a2018fcdf430ea420ccae2fd35b2acd637cb083370cc86155cc8);
            I11f1c07733856926d4d980234959cd48f8b0247270d6485cc57dc3456ba7adbf    = I4d2bf12a647b50d4ab9b14ca939986eb9960c3019be93049f9086529acdfee39;

            I0ed51fa81db29c53a4033d2a60ceccacaba9e1abdc340f1226e4951b8af1d49a = I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f + ~I0e4ad715cc833c775ed97e88f28c4196d28bcee4370205307f4266e1fc572cb1 + 1;
            I6648e8e7f5ebb09e748ceaf1dff7eb3cb073b8d035948f93b25c45bb10b2589f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0ed51fa81db29c53a4033d2a60ceccacaba9e1abdc340f1226e4951b8af1d49a);
            I26f2f2938065d9336a83a2edcb5595f6976c5c434c76d4c44e771cb8a0c685c4    = I6648e8e7f5ebb09e748ceaf1dff7eb3cb073b8d035948f93b25c45bb10b2589f;

            I15f92f05ad628c0f786341269ec6b7aa37408eecb1415a026b776fe4b1ea167d = I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f + ~I1f9214a0b2b730fd678664ec457d15dcc243ba1d68ea198ef2792ac2440608ee + 1;
            I248153dbc85025b19e54dbce1436968e1467457e71047a73fd6b1365aa362259 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I15f92f05ad628c0f786341269ec6b7aa37408eecb1415a026b776fe4b1ea167d);
            I059b4a33ad6774feb79158ff05ecb4287420d94dc0c57650fb90f11fb7fb83ec    = I248153dbc85025b19e54dbce1436968e1467457e71047a73fd6b1365aa362259;

            Id182102124b3765c410c79e6b7560532537d8ce5d243f64cab3c4a73ac894292 = I265fd10cb36e7a3c607cdf96cfd87086b85db27c6103bffaf2cac333af05975f + ~I9d323aa17bffd7ea7a66ef99d4d004ce664a0e7e5388ed24a4d45c69a4d9b396 + 1;
            Iebae6187f539cafedc0df54b1428bc9b57c6aeb3320a5bdc212d444a9a4fbcf9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id182102124b3765c410c79e6b7560532537d8ce5d243f64cab3c4a73ac894292);
            I9a9e162c226e402630bd217ff502dc5aa823ee7c089801803c5ee091b5ea4026    = Iebae6187f539cafedc0df54b1428bc9b57c6aeb3320a5bdc212d444a9a4fbcf9;

            I92c3d579813e542874bc16d04e9aa52c9f79b1b55fab5f166c74f6ab61bb195d = I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7 + ~I88f1c4536adedb4ffea1b595f5fa753329c4aa2187a3245269734a18a122e189 + 1;
            I9b9bf6eb31652e7b62bb383e61221c03099b628ce1f87617b7c90805088c161e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I92c3d579813e542874bc16d04e9aa52c9f79b1b55fab5f166c74f6ab61bb195d);
            If30f29822c81c32a3f153165fbdd82ff6cd9527a6a065627852ca8d5d1a0b122    = I9b9bf6eb31652e7b62bb383e61221c03099b628ce1f87617b7c90805088c161e;

            I552bcbb774b1f6cbc437d0e597e9f85a058a1c86dc9327c0ac420c6cd272adfa = I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7 + ~Id9a38b1906060dc5739f9446bb2dd1a6b6603924d4b7889c931988fb52cfafff + 1;
            Id8b61d2b7d04b31046b959b2e56f86603abcd13532e8c5d7496b769f872bd6fd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I552bcbb774b1f6cbc437d0e597e9f85a058a1c86dc9327c0ac420c6cd272adfa);
            Iec9d3d3ad44a5c22fbedf1fc73a01cf348f8c4b16c5f3f0cf55c85f8d92ca22b    = Id8b61d2b7d04b31046b959b2e56f86603abcd13532e8c5d7496b769f872bd6fd;

            Icc1b7731fd55becb0c39c2ad581762a4053fa931b7944cfbf14ee41929363b6a = I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7 + ~I5502a12455fae3619e0c2297d5e4a8062415aa3ddd8f0bbf67a73233bb6df733 + 1;
            I294ca2d54cee0e207eba2b6bc501af13d7576edac3409f1d345f26fe570947a2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icc1b7731fd55becb0c39c2ad581762a4053fa931b7944cfbf14ee41929363b6a);
            I94452304db6f03a077cc46cd087cc756c098f85885a9c8a60e1860ebb0b23a60    = I294ca2d54cee0e207eba2b6bc501af13d7576edac3409f1d345f26fe570947a2;

            Ib2ff21fa69dd26a3b35833b51981a6b4e03be26d774d933dd860357d347282e0 = I05970991b08e409add39bde806ea896adbd33912e59dfcc945540ff2b221e3a7 + ~I8e6a3df905c8c5778e1fd6e75b091c545389651762d9cb3e0d21b20d8dcee6ae + 1;
            Iee74dd10fa4b539456d95de7258116aa77db37667ec4ec2decfa968bf6f602aa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib2ff21fa69dd26a3b35833b51981a6b4e03be26d774d933dd860357d347282e0);
            I59d79bf88b865cc38882adc0e8d69f2a1556f9cef906cd558730ea7a902de6ce    = Iee74dd10fa4b539456d95de7258116aa77db37667ec4ec2decfa968bf6f602aa;

            Icf03aca159cc538c2d6f4b1b616e5c6c8dc4f66dfc24b50408e54d746671a222 = I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e + ~I554ab27e696a028f48da8ad39e2db6668b57ff692603a9562cd7e8780bfa491d + 1;
            I62b9c19449f50c6d47f459d20978c10e564edeec60593f2213ec4a45203a9b93 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icf03aca159cc538c2d6f4b1b616e5c6c8dc4f66dfc24b50408e54d746671a222);
            I022500b8d9cd3b589fb75b90c1b633a96fdc76c0e3e2ec514cf7b4ff3ccce1b6    = I62b9c19449f50c6d47f459d20978c10e564edeec60593f2213ec4a45203a9b93;

            Id934d373281e6054a71d367d79cddd1549b8048fc9fe481b15c8b8f6099e9468 = I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e + ~I1f070cf569961de917cbd287e7b14a2ad6e04a4474edfb92c095f6e9cea1efdc + 1;
            I85c9fd61717aec721a675c20933429f4e323f13065bcdbf79eee199d97d2e56b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id934d373281e6054a71d367d79cddd1549b8048fc9fe481b15c8b8f6099e9468);
            Id9936f1014242296259237c4aa19452ea56509e2d970ce60c72e7c4d18a66752    = I85c9fd61717aec721a675c20933429f4e323f13065bcdbf79eee199d97d2e56b;

            I381168c5956c61f426a711cb5861a659681cc9f9772accf6ecffd355ce8db307 = I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e + ~Ib423f5e14b109a601cf9e9d403a7b5c0ca0de8d665d065d8f317760c5705071d + 1;
            I23746c5cc5a886c61f469589a55b57fd6e8b77852b50e814c672a2c52802f253 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I381168c5956c61f426a711cb5861a659681cc9f9772accf6ecffd355ce8db307);
            Idad105c150f27de4777164385ed4e2123966f63d2b2ff32add6d18a95be2624d    = I23746c5cc5a886c61f469589a55b57fd6e8b77852b50e814c672a2c52802f253;

            Ic7195dd57a1287cdadc40d619ee55d7a59d4a02e624c74267ab5a631dc66a6c9 = I7c6003dc1100f7e40afedd83325b09245575489d7a9b1c7604eb81aeade0cf9e + ~Ic935d033e29fa4baba415347d379eeb1645c65388d3c7c9858ae48f5a098e2bd + 1;
            I806e92d3c392bf729c0f36bdc2b5d398ef947f073dcc733e4301aab45a73d08f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic7195dd57a1287cdadc40d619ee55d7a59d4a02e624c74267ab5a631dc66a6c9);
            Ice1023bfed1f964ccc66c7d914378cc899ac310a76f3d694302cc688bb560e45    = I806e92d3c392bf729c0f36bdc2b5d398ef947f073dcc733e4301aab45a73d08f;

            If27abe3474af746eb5d14fbe518daf8012c4ae8f65e9972aced680995387a413 = Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b + ~I6996b52f42eb9075a634fcdb07fafaf45c5aa99193446869751c4859e7c1f963 + 1;
            I9fd1bb95c6a2213084ff79a560a6264130dbc55ea0ee6b2702539e00fbfc67e3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If27abe3474af746eb5d14fbe518daf8012c4ae8f65e9972aced680995387a413);
            I372b0e45c0d1e8d30830bd3cac2c3082ec36f9af195380d0e1b7d62712123fa7    = I9fd1bb95c6a2213084ff79a560a6264130dbc55ea0ee6b2702539e00fbfc67e3;

            Ibc36ad96928d2d8544d21273b9764c7dc17dcf79447e8ad92b689f9c33debb62 = Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b + ~I332737561309225f302f64e49e8b3e4aa4dc35344858059b21e146e8cb84a466 + 1;
            I6644cc3a42774e6d8fa09e46158d631bf6b48b406b7981f8feed695d22959203 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibc36ad96928d2d8544d21273b9764c7dc17dcf79447e8ad92b689f9c33debb62);
            Ie98369c31ad7be164b6fc0f16fd6d1a5193f2b00a3eb10ee1cb478b4653b60fe    = I6644cc3a42774e6d8fa09e46158d631bf6b48b406b7981f8feed695d22959203;

            Ia3a1160cab48ed755a51597f93348a5ff2a29df29582523f0f1051175dcfd3a1 = Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b + ~I2d2817ad47b56d0a7ff72c326eabc6e2ffb1819a2748ffe3a4a42d3794cf2fc2 + 1;
            Iae221cbeaae99099c7066532f85d20ecf85ca760a449bb238696d7821a729c21 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia3a1160cab48ed755a51597f93348a5ff2a29df29582523f0f1051175dcfd3a1);
            I80f30106eccbcdd1f0aabed1521d2b09a4bb56a421079ec90f81527a903c6643    = Iae221cbeaae99099c7066532f85d20ecf85ca760a449bb238696d7821a729c21;

            I4b4f2557be01daf1e3a86e3900f7220915b80fb490425d6bfd0e6f2ac3d758d9 = Ia6e2ab2b5aec29f0e218ece9ed700f4cd4945e090ebcf67c3efb9c2c68f95b2b + ~I1f212ee134daea9d568f52fcdce6452048326c2dc243c60d25ee71b95ffea50d + 1;
            I304c658d3b58023c7c85b82e12d5e4eec7336cf6d04c3468e591bb77e4cce5ec = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4b4f2557be01daf1e3a86e3900f7220915b80fb490425d6bfd0e6f2ac3d758d9);
            I81349ebf72720f77a8902dc12d9cf986ddec6f8fe30f7f76f9f4dc54881708b5    = I304c658d3b58023c7c85b82e12d5e4eec7336cf6d04c3468e591bb77e4cce5ec;

            I59d501073967763b8f11f100cc0aa90180a85e7396d40479244bd2a74e1bbb81 = Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb + ~I8e8e17839b8f0cf30290c33a60662c784f062950716903854e36856a58f909b7 + 1;
            I57d74f096ffd259b46eb1b76f49ec20079d2b15d7453108f95f5f6aaf6a272f5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I59d501073967763b8f11f100cc0aa90180a85e7396d40479244bd2a74e1bbb81);
            Ic941f62ac4a004ce3dfdcdfc5312a3be16a5307024d1ad292754532cec3fc90b    = I57d74f096ffd259b46eb1b76f49ec20079d2b15d7453108f95f5f6aaf6a272f5;

            I51dd1d6d9f1dcdab1e85e392e5fffbbb22555f9bc89aaafd686ee55bd8dcd14d = Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb + ~Ic595c984782ebc89b61fa2a64e994aa66eb4979ab1e30e890886355dc247a67f + 1;
            I7e4b87e71ac1fd30a6139a3cf27f76002a1c67adf28eb8d4e382866afa224cb3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I51dd1d6d9f1dcdab1e85e392e5fffbbb22555f9bc89aaafd686ee55bd8dcd14d);
            I65c4ade7c4c23e62f5cd1846b0a739c70cd498087298f54c41f89bbd9677e705    = I7e4b87e71ac1fd30a6139a3cf27f76002a1c67adf28eb8d4e382866afa224cb3;

            If117910f998c5992518fd3258d34731a1dd45db76e7af467934d5c0b8b455c0c = Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb + ~Ibfb48072643b2cdc460b7a667940129aa243be78b6d57abbd483d5551fa36eba + 1;
            I3704a80d3cd58a300a6e4d721e00950f5166111d44d9827c6b492524d4c556c6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If117910f998c5992518fd3258d34731a1dd45db76e7af467934d5c0b8b455c0c);
            I4d548bf4a643564a906a42a32acc4fe6919c91f43890f1b921b9e42100b92e68    = I3704a80d3cd58a300a6e4d721e00950f5166111d44d9827c6b492524d4c556c6;

            I6414021c1267477ff6a5b8899ac081a7f3c840f899c3a08b1b42ca91d37f945d = Ife210366be61f39883479c5d877ceb632b1008531a90c85889267f92eb2ff4bb + ~I3a25f0d4a6f0fa33f493d9aec6fc7a318a826b3885a3cccf04e9b1a85bec345e + 1;
            I4e750ac2d9b11787d2cabe2f06aec65d630b6be5185d7ec5a3efa12565000e2d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6414021c1267477ff6a5b8899ac081a7f3c840f899c3a08b1b42ca91d37f945d);
            Id89fd01703e5a1c53c89a64885698fdf565b791620408fb963b53208a33e7f47    = I4e750ac2d9b11787d2cabe2f06aec65d630b6be5185d7ec5a3efa12565000e2d;

            I5375e515cadcd87ad137d29768eabc89cb773c65f1838f17762632fe6915b805 = Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952 + ~I31ea69d26acd05d303178076eb123a7b2bbfeca82c2690c54323889753261f1d + 1;
            Ia2b84466a2783970d94e38c4a99be0bd22b7e574580adb621eb579e8f9bf81b1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I5375e515cadcd87ad137d29768eabc89cb773c65f1838f17762632fe6915b805);
            I8467f29aa6da06588468e21697c56464c67e4809c135d2d41e38d9881715aee7    = Ia2b84466a2783970d94e38c4a99be0bd22b7e574580adb621eb579e8f9bf81b1;

            I1366c2561d741ee41e937b32668f5b2dae17f38f7ab9192ed8d4670e570096bf = Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952 + ~Iac3e25273f8b972112775f3aa57274eabadbc2da5eea147328f85a941b959bfd + 1;
            Ied4d22813a35e4cb32ffd1cdfddcdcc877dbfc83dd6d6780296ec5c5c9960925 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1366c2561d741ee41e937b32668f5b2dae17f38f7ab9192ed8d4670e570096bf);
            I55ee374c21e5aee6b0ada78409b18bdefed20abbf3dc5716c62daa87b418dcfa    = Ied4d22813a35e4cb32ffd1cdfddcdcc877dbfc83dd6d6780296ec5c5c9960925;

            I4ed1e2ce8c1861ad771d926c40a92a3335c27ed9c927da2c4b4c8d246f888cd8 = Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952 + ~I4b18b20124a63f85e812047188401b685693ae009c87ae337b840a7a3e03f140 + 1;
            I11bcf52f915e80d94647f8fa66ee0dbf0d31537d68a896fd62b4fdfd8e76aee6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4ed1e2ce8c1861ad771d926c40a92a3335c27ed9c927da2c4b4c8d246f888cd8);
            I4285be4ac50db4da7f720fe115c342ad8ecefdf6dbace4af4c9714009ae31e86    = I11bcf52f915e80d94647f8fa66ee0dbf0d31537d68a896fd62b4fdfd8e76aee6;

            I34dbafcdf27f8460fdfd7a329a955300c42889d6f99e9396df4fcf0a80d7e84a = Ia71089b0ed708e18d70ee2052b2dd9c29db42183caddd67a284132947d59d952 + ~Ifbee83b3613941d8ba27021c2fd37d0990a8af8fa3e0399f0f1f8a92ae18d273 + 1;
            Ibc1d752fb7dc31452424184c390d0348180fae8b0901eadef67aac5bfb0bc449 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I34dbafcdf27f8460fdfd7a329a955300c42889d6f99e9396df4fcf0a80d7e84a);
            If37e3544f587a047696dc53e30f6031f848e27a13e2328b2c38a4f51421954db    = Ibc1d752fb7dc31452424184c390d0348180fae8b0901eadef67aac5bfb0bc449;

            I9fbba72f6f8a1120c18220196387259e4e2ef9be67b89f4c4d941bd2716c16b1 = I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677 + ~I41b85a49eea9c0d773ecce66f0023338d3ee5a94e14a87c867a74960d30211cb + 1;
            I26105c08050f06741f732eb11726ecee4899cca05c21e1aa75eefb07c60b695f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9fbba72f6f8a1120c18220196387259e4e2ef9be67b89f4c4d941bd2716c16b1);
            Id9067d2f353cbef30dc828f16a97436418af2bf3e5fd19300471de394f710fff    = I26105c08050f06741f732eb11726ecee4899cca05c21e1aa75eefb07c60b695f;

            Iaf9bb39df39518f42c265087053d0e659319b41a5ce82aad117fb21646fc5811 = I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677 + ~I698accb14122caa36f489e7fc522e39188ee03651ef0c6670eecd60162cf2f0d + 1;
            Ib75010a3db964882380071e188e4d75235be279058fa470c1a758a97a7ab518b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iaf9bb39df39518f42c265087053d0e659319b41a5ce82aad117fb21646fc5811);
            I93150066a1cfdd9e59edd1d42cd2611eac0df4fdfbea33d913804f52dbd895a5    = Ib75010a3db964882380071e188e4d75235be279058fa470c1a758a97a7ab518b;

            I23a214695af25c30f017977039b6522a79e1ede0b71df88555b1a36a613ea32a = I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677 + ~I26c556de81da143a85c36f6ba98648e110114ab97302046b7aec581a62689a3d + 1;
            I32d23e06facbd4ea9378cd4d72ac744cfc0ddfc54bb1c22550b09176ea670372 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I23a214695af25c30f017977039b6522a79e1ede0b71df88555b1a36a613ea32a);
            Ie296c1317a499d9d35191ae9de6c681e2b521a2966b8837ffa470e3de6c8530d    = I32d23e06facbd4ea9378cd4d72ac744cfc0ddfc54bb1c22550b09176ea670372;

            I7d3dd2b2f1be7541867d824bf4cdda33f1e8e6acb187e6f78ee354a9030dcde4 = I4995d7eba85772ecb75824663a725b8c41dd18b265bef16a755c7c3c83bb3677 + ~Ia1c056993094512262fa3f3d38a2a46cd43eb08114e1af8c48ce2f6705d7297b + 1;
            I84baca35ef199aa658e78c93b7dd27049c57dc70d92194ae59ae657ac001470d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7d3dd2b2f1be7541867d824bf4cdda33f1e8e6acb187e6f78ee354a9030dcde4);
            I0aecd8795e3571b4b428903758f7dac78966a9a928f64c26a3e6f00fd61872ab    = I84baca35ef199aa658e78c93b7dd27049c57dc70d92194ae59ae657ac001470d;

            I242b12e2ea6f2cabed454cdd179b9a0b2ea51a43ac2c450f84ed2c650a2cf789 = Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab + ~Iccacefad631e33ec8e54f8261759ca110fefaa6fd9fad08940205708a7180eb1 + 1;
            I7cd8396ac94d8c37d3de99389d6b06115b7d36f1e31faf88cdf01c5662fcbbed = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I242b12e2ea6f2cabed454cdd179b9a0b2ea51a43ac2c450f84ed2c650a2cf789);
            I0bc6fa0d581c2d2fcce482d2821bf87f00bc84606afa8b56d7f4cd88bead4a3d    = I7cd8396ac94d8c37d3de99389d6b06115b7d36f1e31faf88cdf01c5662fcbbed;

            I66e51d57d162e80e54fc2e9bfa91dd74805a0cd6604ef63a5645f50242e2397d = Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab + ~Idb883f1d90a389f89c3e04f54dac20f205951bba3fd0a00e9432498c4def1131 + 1;
            I47f3b89a5acb9ee2c282930b7d311145f48b3aa49a1ebd406b76412db2042fa4 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I66e51d57d162e80e54fc2e9bfa91dd74805a0cd6604ef63a5645f50242e2397d);
            Idfee0ad9592b445c7afa92c1099d49c458d1eda5605ad06e6ec975e2d9103e11    = I47f3b89a5acb9ee2c282930b7d311145f48b3aa49a1ebd406b76412db2042fa4;

            I610a848a26543d03e396503018f1541e8a2647f8c97ebefcddab43e6cd91ad88 = Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab + ~I5059641c5d09a0369f6237643b75899865bff068e9aa8779d0befdbd53a6b754 + 1;
            I40748060a17eaeb7d8f1a828d0767e42c09c2c104161262b5adc72249d128df6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I610a848a26543d03e396503018f1541e8a2647f8c97ebefcddab43e6cd91ad88);
            Ic700c1c29d2fbb8e2e85fd9871082303e3dada09845afca88fd7c35f9d41affe    = I40748060a17eaeb7d8f1a828d0767e42c09c2c104161262b5adc72249d128df6;

            I16852d5801d3a353a9d084a0b9dd4fcc537eeb8277037f64f84d1fd1b1b42102 = Ib04cdb180dd05f2f8f4f9b10e30d1372641ccda9931757a47968f1c2a73cd9ab + ~I61e29bdef580f4f1057d7b4ffb5bbf37c67d3b8107d7979c2fce643282c7d861 + 1;
            I580aa2ffd81e1289f84a7d86e68cabc547ca6c8bb698bb648f6cf57491c18289 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I16852d5801d3a353a9d084a0b9dd4fcc537eeb8277037f64f84d1fd1b1b42102);
            Ie1342b74cd710b1a52ba3de5ca28ee42d03eaf53a42a6cedab9ecb6d987d7b55    = I580aa2ffd81e1289f84a7d86e68cabc547ca6c8bb698bb648f6cf57491c18289;

            Iefb3d17f1de1e179afcfcf9f8d209375b9cffd7efc7f3ae88ca55d6c58b0d7d6 = Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7 + ~I6f52a21dd933b23b7565abd508c69070b8cf652dc313689f62c7f04d7acb934b + 1;
            I89baba2fe1581baa53e6774b196896f7a0c32f88c5dcb0f6ccc7cd4911992b15 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iefb3d17f1de1e179afcfcf9f8d209375b9cffd7efc7f3ae88ca55d6c58b0d7d6);
            I69f8afa3d9aea957a3c1a9f3dbfd8ef8dc6370b228a7f67f0a27113c094992ed    = I89baba2fe1581baa53e6774b196896f7a0c32f88c5dcb0f6ccc7cd4911992b15;

            I1abfb953ea909659ae25d197a2ecbefc307fa6580318bf8dfd723883f2cb242d = Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7 + ~I80c7df909269b691013f9d178bc3e8c896d4d06ef4cc4b0ac42858888ae8b92a + 1;
            I2e381e0df584249b04ed891c499ded7e2d180a403ece202bb96f3cf8041dbbd8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1abfb953ea909659ae25d197a2ecbefc307fa6580318bf8dfd723883f2cb242d);
            I3b017b72afccffaac4ff923e52843d312e1cd5e1123575d6daf4692f81cfe748    = I2e381e0df584249b04ed891c499ded7e2d180a403ece202bb96f3cf8041dbbd8;

            I388e7ed193084e1a629828ccb5e027b54dff58603c1e644f81fa233d8c397511 = Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7 + ~I403d7b440509677065b38ca8634080a8edc4c8eae54a9923c50885861866a7d8 + 1;
            Id539ba7ee7b26dc8f610a6298e8fb42f50f810b490cd75ca72f0875a2271c8b3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I388e7ed193084e1a629828ccb5e027b54dff58603c1e644f81fa233d8c397511);
            I100b4afda393740a5fcf563e8e5fe34d5d7bfc439f2eedd77966bc9b37b3d602    = Id539ba7ee7b26dc8f610a6298e8fb42f50f810b490cd75ca72f0875a2271c8b3;

            Icd26d5b89d292b0466a08a131e8d00b1da2a54043a429e61b02f38a292c980fd = Ie6998e19aa82a9566f525ff1f8f99e09ce7d5def252d03a45ad929b79f0402b7 + ~Ib07a3587e3bfa70ff5dcb296b8595c5d15cb8a94efb13c3e5cc92cd3be3605ac + 1;
            I9826aba6d5de9618406c264016c229e048ccc60817b1edccef930d6e6bfc6a0d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icd26d5b89d292b0466a08a131e8d00b1da2a54043a429e61b02f38a292c980fd);
            Ieeaf4fb83c3c92f18b21f65ff2a951f74693fa6da2ec322ae6a4873d26729f51    = I9826aba6d5de9618406c264016c229e048ccc60817b1edccef930d6e6bfc6a0d;

            I1932bcf87fcb5256afa2f82da25621ca1cc06f6e256ab9b05d1b3589613bbe02 = I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5 + ~I78d7fbedde9ab5751194c52134dec1b83ea8d48c4ad77c0b3eb952143612ab71 + 1;
            Ic211c903aae638bfcdd91aa6d092f085204dad95f7e45bc78c9269816684ce42 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1932bcf87fcb5256afa2f82da25621ca1cc06f6e256ab9b05d1b3589613bbe02);
            I27ac039dc48350ce90d2a8a3953936d5f7c97ec1098fb20d853cd062f2d4a6f9    = Ic211c903aae638bfcdd91aa6d092f085204dad95f7e45bc78c9269816684ce42;

            I807bb4f93cb4990ea3d0b5f5bb5ee1c9e281eadf997a92a32fac10d917439ac6 = I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5 + ~I581a3a40f892233a7bd0dda3bb84e2e46095c27e45d53ed32ef5226f9d25ce43 + 1;
            I14d3a54a6919ec76c17e6d155fed5dd3848ea7e567f997f659d5a09a2100190b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I807bb4f93cb4990ea3d0b5f5bb5ee1c9e281eadf997a92a32fac10d917439ac6);
            I224433de24984b12aa905ae86eeaa53ec459acd68fefdba7aa1e8778abb89408    = I14d3a54a6919ec76c17e6d155fed5dd3848ea7e567f997f659d5a09a2100190b;

            I3ce261f7e73a1bc919627efb495dbeb739b6b9ef526e0d575ab46524d6f50092 = I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5 + ~If15171a1904299c55ffc5b4c9059900188c1c87caca3f4807c4498abe038becb + 1;
            Idfa486a97bc44780268cdfe3738e6c0a3fa58e51f0c4bad523ce7ab24b3fc471 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3ce261f7e73a1bc919627efb495dbeb739b6b9ef526e0d575ab46524d6f50092);
            Ice1b30668532ff63b6ead40f37366b805ea21a65f6fb7067bf9d3b5d08eced46    = Idfa486a97bc44780268cdfe3738e6c0a3fa58e51f0c4bad523ce7ab24b3fc471;

            Ic7138f5e1ef57f1e0d904946b13c6e16a293b6fba7db6266a9c40079e40c8e2c = I7aec2d2d99506db125ee20b66e67ad34234a375bc3ab5ae6220c942ad3f31ec5 + ~I8c443a2690956ee9d0171ca05534d698f75563cd74ec9f4de33c7e8dabe8105a + 1;
            Ib486f88deb674197e70cfa4b28061cca75c06176b05673ded7af5c62ffe15d5d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic7138f5e1ef57f1e0d904946b13c6e16a293b6fba7db6266a9c40079e40c8e2c);
            I2b6551d9c8b14c787afa552e23234fdbb63c8fdb8fb285416ff1b72a38e7d898    = Ib486f88deb674197e70cfa4b28061cca75c06176b05673ded7af5c62ffe15d5d;

            I7baf74b530afc8aa64e5a9f2b7879a0a6573eca1818262c1ac817c5940b0fd75 = I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093 + ~I3fe543ea18333fd169c6d6e692a5b42232e8abd2b14072a4daba9bacbe921d2f + 1;
            I958b582efc12bab546e1da193b5687e5c19e401a03bc7d6fa5c7bb1108ad911c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7baf74b530afc8aa64e5a9f2b7879a0a6573eca1818262c1ac817c5940b0fd75);
            I24ade58e2190b73f141a858e6812d93a49203181d6d427a29415d014a9cceec6    = I958b582efc12bab546e1da193b5687e5c19e401a03bc7d6fa5c7bb1108ad911c;

            Ide134ae79fa666de582a416826cc2d4a579d888b98b3b820f3c5e445767d002f = I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093 + ~I7a52610226b8a85bdc6a0b49cd74cc644d2fad0e8f98ee24c46ccd3664d0af24 + 1;
            I1fd2d5d75d3b779da0e3e1c3c66053704eac857ecae818b79be59c72e04e0b92 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ide134ae79fa666de582a416826cc2d4a579d888b98b3b820f3c5e445767d002f);
            I55affee832ae4e480ffb916ce8a5e3b12fb6429f1ccee3a8f9a668aeb8352f7e    = I1fd2d5d75d3b779da0e3e1c3c66053704eac857ecae818b79be59c72e04e0b92;

            I76566fde1f58392124d201e9b66f3a221ea658b9be074b36c54773b34997faa9 = I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093 + ~I9efd4f4bd4d8dfa270cb1c5a2e3f5c6cbfc3c5b672540ca268e0765170e6c748 + 1;
            If5f8b823e2d28fc1b521af24083f2fa271ac7a29129e8cc1cf8c5eba46fa4583 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I76566fde1f58392124d201e9b66f3a221ea658b9be074b36c54773b34997faa9);
            I3f2f052f1d132cf1a83172a044968741665a7b85e421658976109057a3d00ba1    = If5f8b823e2d28fc1b521af24083f2fa271ac7a29129e8cc1cf8c5eba46fa4583;

            Ie8db353155b2c11a919ec581a22860b11997a2ec74cc8be6c36b04716c9fa558 = I2974a4c4abea9efa23e0dde3ed6f33fd69512c386e814d1deb3775310c83b093 + ~I5dcbde9462714577263040534f0560b0c126ba001e959add92d0529cbc94bd9b + 1;
            Id068fbdc476f28f1695939e90fef8a08e2cd9434b1368ddefb14cdc950a76a2e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie8db353155b2c11a919ec581a22860b11997a2ec74cc8be6c36b04716c9fa558);
            Ibbe3cd91dfae5930a6ae5799a27b045ce6e0c59fe00a38b5fb4b1691949847f2    = Id068fbdc476f28f1695939e90fef8a08e2cd9434b1368ddefb14cdc950a76a2e;

            I54f9f4218a4fc5202873aa8c9e0fe7564af5e7c244d438f8c662117204056632 = I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a + ~I7dd3baf838ce22ecec10d3c1a3d0dd16582497f9e447038aa46bfd49571fcb4b + 1;
            Ia193fe333281870ef7d810f61721dd6c5557204828bec993bb47bf37c9ab46e8 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I54f9f4218a4fc5202873aa8c9e0fe7564af5e7c244d438f8c662117204056632);
            Icbbfd81a7f066da629076f9f7c26eb457be34298a6518cf45e67bb39e74f5f2a    = Ia193fe333281870ef7d810f61721dd6c5557204828bec993bb47bf37c9ab46e8;

            I7e64afd49b1b6224dd6a8f10660ef803524895019ee93a630209c21f66fdfb26 = I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a + ~I0dfd7663ac138a56ce3fe38c03c10675da9e417e38f56ea0fa4f9f1902d725b3 + 1;
            Ifedd253513982e9c918cb3e4a65f4a6034759bb977b8dc42b00ce4a97cbdd5ac = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7e64afd49b1b6224dd6a8f10660ef803524895019ee93a630209c21f66fdfb26);
            I762a7e10d310500a1080b7b46a9a30bb003c7a7d48011e96501a647e1de0cb66    = Ifedd253513982e9c918cb3e4a65f4a6034759bb977b8dc42b00ce4a97cbdd5ac;

            I813a94c07943df9b170773639811bb908b1dafdb2a89be0d53e81e2b98faecfb = I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a + ~I94ba926e07e8b3cbc5429ff6bf73020e95dda7b7c0059dc10ef646b2980bd80a + 1;
            I6ebc1aa84acf73083137d13ff8d907175d13ac8031ff97e186840f851182fa28 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I813a94c07943df9b170773639811bb908b1dafdb2a89be0d53e81e2b98faecfb);
            Idc9ce24f8fd9ca7372ef25d9e2b8414a4c8051c796f9ce64b91a6f3e70faeec6    = I6ebc1aa84acf73083137d13ff8d907175d13ac8031ff97e186840f851182fa28;

            I3a3f389915c4e6367d45081282db8a902b0acbee573fbb0da4c5d935043bc2ff = I3fc0df00109f90932c48899cf7c2cf31548373581e9bb59223b808f0be62c71a + ~I3872eb448ad521cf99b3a9d07ecde078320dcaaac45bd387137deaf5dec956b3 + 1;
            I7d39228cd05d50c7151740b19887493bd52a4504ce3b2090dc14baba0b03affc = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3a3f389915c4e6367d45081282db8a902b0acbee573fbb0da4c5d935043bc2ff);
            Iffe887b6857424a57f7b7bec156197556dd869c44a2eaa660fa66760cd88888a    = I7d39228cd05d50c7151740b19887493bd52a4504ce3b2090dc14baba0b03affc;

            I8a0fa39f59af823fa6b73d097b287483857fcaeb20ec459e4fb5812c8774a796 = Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223 + ~I4a4338f7d9bbbf60ef4dc6e821d22619911e41300b49e83d57a0a959218a05ae + 1;
            I3369e19a0c3d22229db15bfe65a56d3f45222928f405a8c28bb7dd5f5f6a96a1 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I8a0fa39f59af823fa6b73d097b287483857fcaeb20ec459e4fb5812c8774a796);
            Ie7328907da6b377ef494c54a5e6fc2f90992a99258967af4bc2205d0d42e9db1    = I3369e19a0c3d22229db15bfe65a56d3f45222928f405a8c28bb7dd5f5f6a96a1;

            Id0ab6ebd5d082a3d961cb6b58b59350db5bd2c3d85c08a14901f6573b80fa446 = Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223 + ~Id1fb56c160d418b26fe2b51dbe78addbbd2743e7a342e0b6bebd2e8d3cb1ce99 + 1;
            I6f621b228fdc4c92d7bd7bcdfe69acfae45c715d228e99fc566de1e72163faf2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id0ab6ebd5d082a3d961cb6b58b59350db5bd2c3d85c08a14901f6573b80fa446);
            I98616ac468624d04fcf2487684bc23bd20a87b719be4d4533f987ecb1bcc8d5c    = I6f621b228fdc4c92d7bd7bcdfe69acfae45c715d228e99fc566de1e72163faf2;

            Iccaddd2cbff52541bba9854cb236957b9ff6e50e07f2be5f60b08fb247e44962 = Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223 + ~I89b44baf278e7cf024304d7bc6cfa759a735e5da0cf25a96a83e29fa83d12bd8 + 1;
            I86236809a2da5af49885cd9a573af96295f9f16b79a784c7803681cf5494076f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iccaddd2cbff52541bba9854cb236957b9ff6e50e07f2be5f60b08fb247e44962);
            Ieb0d5850e57aa2cd83ee69ba71c85e9e047a9cc5b195da367a9f042a39559f47    = I86236809a2da5af49885cd9a573af96295f9f16b79a784c7803681cf5494076f;

            I9a6d992471765834fab17a42d3d419bedec8e1fa9eeb10617930e06d2aa2e5b8 = Ic31eee745f1d3ae70057b498f648074215f42fb1ee1d5acc271d846a64e87223 + ~I144443166f296f7fdfd616492bb4b1fe44e0353fa6b0fc822b3aec0c1ea0c894 + 1;
            I0bda102a3a10c710d14ca95940f86071834d6ed6cad335022b18ff8f2cee8602 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9a6d992471765834fab17a42d3d419bedec8e1fa9eeb10617930e06d2aa2e5b8);
            If6bf4d8f739928e726bca59f6307a2b78966853a5aeae6bb7dc4786660382ad9    = I0bda102a3a10c710d14ca95940f86071834d6ed6cad335022b18ff8f2cee8602;

            Ib78e3653ad432d8c12b68d0085fb8deeb5405ec0571e9153bf204f598fa23baf = If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911 + ~I9d7b0f41f5cd73f907351990b23117fcaae4302a36d194e6953b54d40361f8fe + 1;
            I00dc832ce34e281f748daed4bf56bc03e171d8124f2c72f7627ed6a5004de894 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib78e3653ad432d8c12b68d0085fb8deeb5405ec0571e9153bf204f598fa23baf);
            I3fc232b4e4ad45bd25aaed0b1306112944d63174fc4f473899349954e94895cd    = I00dc832ce34e281f748daed4bf56bc03e171d8124f2c72f7627ed6a5004de894;

            Idb9e9500623a940d82d7b77b7c613132875cd4287eec27e495a5d2a1fdb16f6d = If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911 + ~I8beede7aeefea570e5c65a76dbc5ce1f4eb114e444ea9b4636258bcefd9d5f34 + 1;
            Id5fb94774f7af4bb8c727a46f588f1266ec3fde633c58ef0844ea4f486782842 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idb9e9500623a940d82d7b77b7c613132875cd4287eec27e495a5d2a1fdb16f6d);
            I07c430087a2a880f756db41ba39cef794ad6d3b28723a7c22df5aa719bf585c2    = Id5fb94774f7af4bb8c727a46f588f1266ec3fde633c58ef0844ea4f486782842;

            Icc42075b4ed713ad08010e19baf3a6ca84a9dd07cdfa71d60c1b6d05634320db = If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911 + ~I102751a9d577151cf6f780ced3299363623ab308737d8483ccbe02118244d2bf + 1;
            I7fb0278bccf79ccd873d9a4bb72a48982ed0d6c1a8702c009bde652c84c90acb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icc42075b4ed713ad08010e19baf3a6ca84a9dd07cdfa71d60c1b6d05634320db);
            Iff963f656b33e8c5d0b4155f3d4ce0be5ec1c056727223d45af4ae070b006272    = I7fb0278bccf79ccd873d9a4bb72a48982ed0d6c1a8702c009bde652c84c90acb;

            I611cde8f0d43b4ca69572460c144fab6ea9088b62f7ee7ca6b2618893e002359 = If2dfa6763dabcb3d74d527102c1a0a0acd00644843f3908b293e60a3b65a3911 + ~I5445f1e35f9039ef623a77ce395c2a888153749fe8226e9b844b271c1c69d760 + 1;
            I345d4e8e18ce7ca6151e381d432ce605af1865671c5aa141b209d1818e2c06e0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I611cde8f0d43b4ca69572460c144fab6ea9088b62f7ee7ca6b2618893e002359);
            I44d78165b52487e966d2063495d2b76b8086031f3d3f0bac7713717f1e56b721    = I345d4e8e18ce7ca6151e381d432ce605af1865671c5aa141b209d1818e2c06e0;

            I41e79867cf93976d9e1db38f48b70e6fc09fe4ec448856483d064ed9ed2f5055 = Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8 + ~Ib0de9295b071389ca7b6bd34f7c9371614337b0be04ccd9ab9819a8e39ade463 + 1;
            I2b2c44feae2f93582dfa6ceaeff78800b79465d7cafdf52289855eba9ba3a236 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I41e79867cf93976d9e1db38f48b70e6fc09fe4ec448856483d064ed9ed2f5055);
            I6e5de0450866fddb6d15781d26a3df126ea57faea36d172ff9c08fbed711ea47    = I2b2c44feae2f93582dfa6ceaeff78800b79465d7cafdf52289855eba9ba3a236;

            Iad7a7d92a71ec5a2a4ecfae6f78716866da577038b41a649d32a5c4db56257ca = Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8 + ~Iae16b002804d17ac9e2c9655dda031f3f0ac10d703bc42079ee2a5fd3ede604f + 1;
            I1d109f4a8531b0b430e5010ec4e2619c94fa8502f3979e8450c9b1d09206660c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iad7a7d92a71ec5a2a4ecfae6f78716866da577038b41a649d32a5c4db56257ca);
            Ie4db811b4d839e478783694d956589c702666e122689ec06c5fcd299c782b1a7    = I1d109f4a8531b0b430e5010ec4e2619c94fa8502f3979e8450c9b1d09206660c;

            I73866569df6c4e95ef7273a1370e9da252db2d74b0df1884bbf87a80a05a8fc7 = Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8 + ~Id9db55519cb1208a2555678410c950b6fb31e5fb04a0ae12d6b0a9de4d750b43 + 1;
            I6a87ff2f8cc2aef5244068df9185b2f8a6b899cf3e6ad460439150b1f2dee99c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I73866569df6c4e95ef7273a1370e9da252db2d74b0df1884bbf87a80a05a8fc7);
            I23072d2753b8750a9cd8da42f6ec9fdce24f0ccf4c201e983c3aa96963421ed3    = I6a87ff2f8cc2aef5244068df9185b2f8a6b899cf3e6ad460439150b1f2dee99c;

            I90c36434a94834ebe700c144c2feb5f0b2a543bc43692f5a23b5b5495d417c64 = Ie7ab776436951de2bf23d5f129d8b172e1fab18d833a7a639cc4593e2630b4d8 + ~I5d9ebd6a6829c49b0e41f700d29bf8acf06a5dd87192846e5ca204ea8bf563eb + 1;
            I645eb770871cffae4c361144a6b3e428d61327c7379b25e3de9ec083b7d9e299 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I90c36434a94834ebe700c144c2feb5f0b2a543bc43692f5a23b5b5495d417c64);
            I96d2ff73be5717714513ef2406648446833f53abe34481e91be763d63d3f2d09    = I645eb770871cffae4c361144a6b3e428d61327c7379b25e3de9ec083b7d9e299;

            If3ae39f173044773979d138817d4e808bd30278aafc2968e47e95c79c1bdd88e = If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd + ~Ib398240cd12e68fb5b3ad4842123a4a16f27cfcae3db8bf1f38de24b82e272aa + 1;
            I1fc6e041dc759bd5cb34a694328c83cce92d4169f00f674238fcd140226fb7f5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If3ae39f173044773979d138817d4e808bd30278aafc2968e47e95c79c1bdd88e);
            If7d7e9843a2eed7a0478c5991a13e140b1ab83460cc8ea6a3bf24a85b8d8ae49    = I1fc6e041dc759bd5cb34a694328c83cce92d4169f00f674238fcd140226fb7f5;

            I417c9ec039c09269659f1426df4443750e00755cf0694b0fe5e508c563e114a5 = If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd + ~I7e3620302652666ddabcd16531a36e7af51722c39bffc4224f256a34ca33109c + 1;
            Ic803fc5440f03ab206425c2100f94823b03ff2a6d6c238ed7407fdf71237986d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I417c9ec039c09269659f1426df4443750e00755cf0694b0fe5e508c563e114a5);
            I61ea75f5f583a43e3691ab2462210c213f53492dd6a4a0a41abc406a7a828bd8    = Ic803fc5440f03ab206425c2100f94823b03ff2a6d6c238ed7407fdf71237986d;

            I3351df654db39d7ca929147d06b79348195c4dcac3d4f398ef2d7d4491a151bd = If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd + ~I29e9674dcb3b06489c5f9017b95878c6a75503e1dc4e2ba4c9c6a7a7cd74d885 + 1;
            Ice1dfd35c5faf0569fc1f6572561e2931d4616abed72917aa2f79010b9949786 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3351df654db39d7ca929147d06b79348195c4dcac3d4f398ef2d7d4491a151bd);
            I2668038e4b55b5d2fbdfcb8fdc56d43beaf4546ba92b39940b8f055a51d7013f    = Ice1dfd35c5faf0569fc1f6572561e2931d4616abed72917aa2f79010b9949786;

            I76e78b4f2c67b24b90b5ec2d4ad5f189296fdd4f21eb6eb8600fdfc9dead405d = If820e7019d1314708ad446f3b0dac6ae32b20beeed343bf05994e888c2ab60cd + ~I7e26d67803410d5079a43dbf6053aee09ff9b0242133282679c3beffd05aae02 + 1;
            Ida74a7b5fe7355a18199b5b942096f1655f787e2b340aa6954243923045f59a9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I76e78b4f2c67b24b90b5ec2d4ad5f189296fdd4f21eb6eb8600fdfc9dead405d);
            Ia29b333453d0a00fb718748060cc9eb198035cf24697fefdcc6b75b450e5fa6c    = Ida74a7b5fe7355a18199b5b942096f1655f787e2b340aa6954243923045f59a9;

            I9a7c4404df96e54123d0a04369056ed0844a3683e09535b029ff8896fd7bd60e = I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362 + ~I9b494d3414d329e4419da30566795e7b36627870c521c463cefbeb7b48196d3c + 1;
            Ibf7568c1b00603b724362101a10a23918bd964f364af6cc21399eca4c9a7f17b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9a7c4404df96e54123d0a04369056ed0844a3683e09535b029ff8896fd7bd60e);
            I9c17b85d3c4d97f0a7093e8007d812455859adb691cd79d2e41e78f95c44d2d4    = Ibf7568c1b00603b724362101a10a23918bd964f364af6cc21399eca4c9a7f17b;

            Iddb4bf2e6f1f1c5a0c910c4939447f53a9794ded6793cf9fd33eb927ff22833b = I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362 + ~I3390b463514e772ff0afe74698bc4850014fbe363d105ce3d0e8810706977682 + 1;
            I636a373b59d09734f347126322958163d4e21351a4fb1f1acccc9209429fd38d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iddb4bf2e6f1f1c5a0c910c4939447f53a9794ded6793cf9fd33eb927ff22833b);
            Idb9949cbe1d38f86e61e1cce9211aa264e0abfb2ea1afa05be251144a4a081b1    = I636a373b59d09734f347126322958163d4e21351a4fb1f1acccc9209429fd38d;

            If0c7c112ee1274d779fe816a1d31c0f6c98d88491fb96633839a9ee0277d1a88 = I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362 + ~I49a96e94f51c41ba36bb7a8d466771682602e2dbd6f65e13d7e858a60b554f3b + 1;
            Ifb235b2a210906a94a1dd95f01a9adcaf8fd76e786707e99bbfa8f0b4bf36e18 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If0c7c112ee1274d779fe816a1d31c0f6c98d88491fb96633839a9ee0277d1a88);
            I18216dc1eb7be60021a2be1d64303e6b9838aaaa2a9b1e6bdffd2a3789661432    = Ifb235b2a210906a94a1dd95f01a9adcaf8fd76e786707e99bbfa8f0b4bf36e18;

            I107b0aecdac212418e4f0054f31ea2a9e89dd7d4620ec8fff0725e7d29414853 = I66b5651f8fbe3ba1871094d322cc089670618e25393836718b1c459dac6df362 + ~I685960b47e49f3ff64eca0e1f26387605e48d325d533550beca6bd6d0f3abbd3 + 1;
            I9f513306dcc73f879dd824e41b5335820c03331e576edc90cf579cfeecfc74ff = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I107b0aecdac212418e4f0054f31ea2a9e89dd7d4620ec8fff0725e7d29414853);
            Id8f0e532c3fc4af615d6cf0967f8a54e6971c1f3572b4383c25360f5f8204ac3    = I9f513306dcc73f879dd824e41b5335820c03331e576edc90cf579cfeecfc74ff;

            Id2edbcc00e89016e0bd07ccb9dfab560cc91bf111ce3b460700435370e90e2fd = I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c + ~I29d04420073229582b38d6b3f7d9d638351e92073269d5528b09b080e5fd5670 + 1;
            I54e17ea4294cd67ff4fe7c421e38999b0b6c6eaac95124d86c6f19863061e935 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Id2edbcc00e89016e0bd07ccb9dfab560cc91bf111ce3b460700435370e90e2fd);
            Ia59883b6b96f3bbe38c2326bfca00e25d3b596e7ddf9287bbf70107666855849    = I54e17ea4294cd67ff4fe7c421e38999b0b6c6eaac95124d86c6f19863061e935;

            I35e88d9a4df07df57aa080c63822b5e79435d28c2f9655a449bd68dcc6aa7709 = I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c + ~If07308cb71758beb15e4a33e3770aba8021bd5572128b9bbc1c8db48e7f807b4 + 1;
            I122b25621999aa119574ea30fab73a0dfa43bb5da1e0e76082f0844cad371a4d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I35e88d9a4df07df57aa080c63822b5e79435d28c2f9655a449bd68dcc6aa7709);
            Ied4edbf18ed0371b7d1ffd53ca5d98f1344d1640b4ca9733d97af5ba5c1c2a5a    = I122b25621999aa119574ea30fab73a0dfa43bb5da1e0e76082f0844cad371a4d;

            I93523e2e245808a8657c66a68778e78a2b7d90f2d076f0be05a4ce53d5803d17 = I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c + ~I4e556f27c558f3d1f76d2ed4a3f0b1a68d74e5c0ce6370b9eec599e7f76f8bbf + 1;
            I32549ac0c631e47367790a831498738385979aada71ed9fa5d238c4128be632f = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I93523e2e245808a8657c66a68778e78a2b7d90f2d076f0be05a4ce53d5803d17);
            If9a4d7f44a518a3ab1ecc6bd5d4e05d8e8f78615ebada754f1ef1e7b13a0e956    = I32549ac0c631e47367790a831498738385979aada71ed9fa5d238c4128be632f;

            I0e18a6aa6a4f5814b2c895163df2b575a04229c654840b386f7654e0765ca631 = I0648a322ab540401b951800e8123a0a61c4a0fa58d22017fa3d2fc9d387e9c4c + ~Icf75218ad23cd1505d2d69d09c0305642a8be48b8a3b7aca4aa4d01a564ddebf + 1;
            I9ba7035cb5eb95ebff5d5d7e549a4ade921979bb4fa7e27f5810134ac2890d2c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0e18a6aa6a4f5814b2c895163df2b575a04229c654840b386f7654e0765ca631);
            I53fa59c42044794f03f617ff512486e58e173121f75b8dc3eb292e9246f7740f    = I9ba7035cb5eb95ebff5d5d7e549a4ade921979bb4fa7e27f5810134ac2890d2c;

            I0911515aa6dcfc8293b4c33ec6d3d7a6227c26e3de3ad8fb3aceca8473c37bc1 = Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7 + ~Ia55512c30a26e336794d389f3700b9153cea83619467b731571ba72a3a9374bf + 1;
            Ic14e91de88b33f4702b25a3e0b4485ba5165438366333847b3e2687934315ccd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0911515aa6dcfc8293b4c33ec6d3d7a6227c26e3de3ad8fb3aceca8473c37bc1);
            I9ae27a7b654a36e4265449d861213978965e4cc3bc7f36b77c6a77cde5e24f77    = Ic14e91de88b33f4702b25a3e0b4485ba5165438366333847b3e2687934315ccd;

            Iebc32b1def039cd8820e6149458d4008738f72a7ab9f73448bd352b362c0c852 = Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7 + ~Ic46278073f42d4eba79499cd6293cfcb33a74310e7b2ed4bff06f5cc63dc9ebd + 1;
            I119671afd256f916b0acec0f5212868cd2dab6bbbd5b158a5fd37320253cb913 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iebc32b1def039cd8820e6149458d4008738f72a7ab9f73448bd352b362c0c852);
            I9dd84c850b5e32710685c595cad935e3249afc0132b04ad8dec94cf13e16faf5    = I119671afd256f916b0acec0f5212868cd2dab6bbbd5b158a5fd37320253cb913;

            Iec3e7529badea1bdcf7d907613c7e25860e379167f064645f36c73bd50d9bb7a = Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7 + ~Ife11a6b34a661bffcf9f0147459d2f5a23d6c5460c59142668ee0f0506755225 + 1;
            I3350bfb01272aafbeca7b9bffcab3434116b885a4ecc32cd92680d122656906a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iec3e7529badea1bdcf7d907613c7e25860e379167f064645f36c73bd50d9bb7a);
            Id59c354fd382f5bb1b276d565cfc2a0d55444ebe928c144c3d0b5513d53e3787    = I3350bfb01272aafbeca7b9bffcab3434116b885a4ecc32cd92680d122656906a;

            Iff7936d861e3a88db1b8e9c2041b7f61a956e483c47f8f16d721acdb81f69c3e = Ic4ef1e901a5bebf22b640d40311ddd83379442eab80a261d827a174ccbc723d7 + ~Ic9adc8e66938cafc1f6974ab9e2fd71a29bcd6520e6fca93ce7bab4815494ed6 + 1;
            Ifce65e25bb01c5dd7349a1766ec452a1658f643d6bbe1f877493527cb46e568b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iff7936d861e3a88db1b8e9c2041b7f61a956e483c47f8f16d721acdb81f69c3e);
            Idab4a7def7105c2e615a9138bf503482df9a2c434aa1ee7c4937acf6d0e6bac1    = Ifce65e25bb01c5dd7349a1766ec452a1658f643d6bbe1f877493527cb46e568b;

            Idcb6f68f9742159aa2fe6947a2f9784ccd2b9d36bd3864ac8b6b38c842f5c5f4 = I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13 + ~I0421a9a7aa72d6f574071ffb4c65878f997e6dc2b605f0d8b351358b08c47ce3 + 1;
            I000e12e2ac3967d4da10fb33efdbb5d6e58d70ec6be81408ba9b7a0995925edf = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idcb6f68f9742159aa2fe6947a2f9784ccd2b9d36bd3864ac8b6b38c842f5c5f4);
            I0d0ba52491ed5f98c69d74967cefc454cb2be9dc40bbc5bfe16c8ace0231dd70    = I000e12e2ac3967d4da10fb33efdbb5d6e58d70ec6be81408ba9b7a0995925edf;

            I925b92518cdbfa9b8934753a60adb3c96413a57c111ab4beade1b677548443a9 = I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13 + ~Ia84ec437292f1ad3e702b4fa896a4f545cab7253574d294243af0c1e7de47155 + 1;
            Id202333f4219877a36045cd10102973d3a15c1dc91156e14961f1d09744c6a6d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I925b92518cdbfa9b8934753a60adb3c96413a57c111ab4beade1b677548443a9);
            I05291a3275d232592dd880dda626cf60a03a62c655a2cf4b811f5325a07eb5e1    = Id202333f4219877a36045cd10102973d3a15c1dc91156e14961f1d09744c6a6d;

            Ib7352b278443169fe5c6f9133c12c026cbc017f6a07531cd9c93b8d58344123c = I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13 + ~Ifc38f7d8250994e5e62716048122eabe81722a32478caab729cfb06aacfc09c2 + 1;
            I9a92d30f7a49d8556b1c480dfa0ab3a0dfee73aef8b8e5caa76e25a3df6742c3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib7352b278443169fe5c6f9133c12c026cbc017f6a07531cd9c93b8d58344123c);
            I141f0199ad8f1dcd707f6b0553ebd7fd04217fb960f13cf25e98511ed91bc7aa    = I9a92d30f7a49d8556b1c480dfa0ab3a0dfee73aef8b8e5caa76e25a3df6742c3;

            Ia8379750d4b5cb8da49adad32a77ec592f600fa74c5e099458eeeeb93ad133f0 = I37503844deac3cf45931e769cbdf17eb117b6dcd59576a1c1831f47fc3099e13 + ~I4f8e5bee14ab1e584593fc15140a36cf071f2949f1bc86fc3fb7dbfdeea7343c + 1;
            I45ee0619e5d6be949b89b7356b7d5a6c42d33e44c5a8885fe69eaacfc56ba8ad = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia8379750d4b5cb8da49adad32a77ec592f600fa74c5e099458eeeeb93ad133f0);
            I11a01802ccb6a01458a2cb2be3dea2f663acc531821edd809b95e10fb5a2def7    = I45ee0619e5d6be949b89b7356b7d5a6c42d33e44c5a8885fe69eaacfc56ba8ad;

            I2d2b275c4f7f134ee6a3999c3f0223d6b626df4441f891a9427d3d8f1f725fb7 = Id6e462224a7c7f18670d48e3a7c6d35465875f9638395e7dd87b3c494985d418 + ~I6efd033a5e005d772ae427cab43bfeacb72354d6905822aaf8d484125615d0f5 + 1;
            Id94d619696cf4cb1820576796ffef7f4fbe3a8a300c5fec44516ec9797164636 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2d2b275c4f7f134ee6a3999c3f0223d6b626df4441f891a9427d3d8f1f725fb7);
            Id76b3104f5a076b0f43f85da8b35a62b36a68d76bf8f26ff0667e085b37ce0e1    = Id94d619696cf4cb1820576796ffef7f4fbe3a8a300c5fec44516ec9797164636;

            I60ea282a4be819088dc3a40aad4a3031c831802d89e57d4c365a1a4d4ac86c3f = Id6e462224a7c7f18670d48e3a7c6d35465875f9638395e7dd87b3c494985d418 + ~Ia6058d7a3749f21a827ae6a0f4e792d6cd62ab37d668d607861bdf3985489d97 + 1;
            I82f65771b72b94319cef82f095d5719ff7dce631f5bc2769ca69634c978bb4ec = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I60ea282a4be819088dc3a40aad4a3031c831802d89e57d4c365a1a4d4ac86c3f);
            If5b73982b4248c4d2cc32bc28f0df8b37553ac0b034c0ebe3009bdfee069f642    = I82f65771b72b94319cef82f095d5719ff7dce631f5bc2769ca69634c978bb4ec;

            Ieadb5d27e6ce4c37e58646b5eacd57fb1a249461f9d16576dcc8bdf46bf4f3d8 = Id6e462224a7c7f18670d48e3a7c6d35465875f9638395e7dd87b3c494985d418 + ~Idbadcb95f603dca2fe62a931973c10429cefef4d6cad0b8e46cf34b2f7c7907b + 1;
            I6566d75140a54ab2f2f601ec74a46508751ac02ee7bf86bee304dfa07d54c8e2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ieadb5d27e6ce4c37e58646b5eacd57fb1a249461f9d16576dcc8bdf46bf4f3d8);
            I9e3cbc961652bd76ec24ad12037b6384d8690af30372a8e0e5a93c57e4fb7b70    = I6566d75140a54ab2f2f601ec74a46508751ac02ee7bf86bee304dfa07d54c8e2;

            I1eedc611ca90fc435e769af408fd45a0299a28c0ad26468af7e870bb5fa26608 = I2c0782e7324e49c90f18114dc327f50948f9bf80b906f202a50b101832a88baf + ~I73c8c2e52e23d992ea9758a361fb9550f0ac7f08bb93b6b26c6fab3b234720a6 + 1;
            I3a570d5967f92b4061a618a46c8d71292ae290fc212c5e3356651a7a69c22da7 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I1eedc611ca90fc435e769af408fd45a0299a28c0ad26468af7e870bb5fa26608);
            I7107302bbea73f0e5ff5ea2791a6d536cb04a165b68ef03ebeab0c0bfffe92cd    = I3a570d5967f92b4061a618a46c8d71292ae290fc212c5e3356651a7a69c22da7;

            I4872d474646c996a00b01718661c079771beab1291ba697119f4a0163b5b061d = I2c0782e7324e49c90f18114dc327f50948f9bf80b906f202a50b101832a88baf + ~I3a8f6218aa06df768133a9b95140db0cdd600a5d1a04a2004479693cecd87571 + 1;
            Id348d892485f4cc1abbc4a897aef1fb7fa4f27c61ff633c9582a1bf733f5d55c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4872d474646c996a00b01718661c079771beab1291ba697119f4a0163b5b061d);
            I561f05c657c3171c43fdfbb59215727da59d919f424597533b1890f7afe7cf07    = Id348d892485f4cc1abbc4a897aef1fb7fa4f27c61ff633c9582a1bf733f5d55c;

            I521983a9bbafb4754207a50436a99446235ae7c9cf0070958e99082cc336cc38 = I2c0782e7324e49c90f18114dc327f50948f9bf80b906f202a50b101832a88baf + ~I9f94e32610a6e83f5ca5d8eb0ad81277c7226ae8ffa7f1e734959a614bf1edd1 + 1;
            I0697f4ec5a674060a0fe012ca040842a7e13ab1391df2b3d09398a7ca857ba3b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I521983a9bbafb4754207a50436a99446235ae7c9cf0070958e99082cc336cc38);
            I81789766f2008122a36b608dce3f08425ac203a154b4e43f915e0e3ef19fa022    = I0697f4ec5a674060a0fe012ca040842a7e13ab1391df2b3d09398a7ca857ba3b;

            Ib0e28df62d3f3d60795ace1cb4975098004b434da3773f09b2f829c6ef7a8b21 = I3d8ccc88024eed4b5d118a6c3b8c06553fcfc8645a8569278e7e7e8d3b41597a + ~Iedb10f981e08498950a50589d8c2fd5dbff191f233da39d5819ddf2dc5172651 + 1;
            Ifad69639fb069c42f4ba17d17a3313ac3414b948dec1f6ad011824925fc5a7a9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib0e28df62d3f3d60795ace1cb4975098004b434da3773f09b2f829c6ef7a8b21);
            I678953f2ad317e167eea663eef2246d68cc67776d905877573ebcc39188a9a4d    = Ifad69639fb069c42f4ba17d17a3313ac3414b948dec1f6ad011824925fc5a7a9;

            I2a58a1a6247cd23a2e2d4ec408d68ca9f77d6331a8a67f975dfe0a1db72f2bcd = I3d8ccc88024eed4b5d118a6c3b8c06553fcfc8645a8569278e7e7e8d3b41597a + ~Icf3a16773d04781aa96eb511825cc59c609fc887b464a86c7839c57ddbba37db + 1;
            I604729a7799bbcf6bc10010a36ab4d0bd909a52c6ea58259e7c532c28c19b1d6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2a58a1a6247cd23a2e2d4ec408d68ca9f77d6331a8a67f975dfe0a1db72f2bcd);
            I048fdd325368b2b72c83a32e9ac2c0208f392416f178445db74ceeafe56c8408    = I604729a7799bbcf6bc10010a36ab4d0bd909a52c6ea58259e7c532c28c19b1d6;

            I2d712b4bb4e09ff4a0ff934bbaca37083bfe3fdd143d20c9f85ec220700af40b = I3d8ccc88024eed4b5d118a6c3b8c06553fcfc8645a8569278e7e7e8d3b41597a + ~Ie023df7145a8643ec413fd62bad9e4dafc719f7c882ae969eaccbce255ca7748 + 1;
            Ic42634514b28215593b2b52782e8b58dd3f1e9e4276619e8603c5de34b4acac5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2d712b4bb4e09ff4a0ff934bbaca37083bfe3fdd143d20c9f85ec220700af40b);
            I16b1a9836d7b38707938eb48bf60f17f049403d2fd29d5245798fd1ade1c2531    = Ic42634514b28215593b2b52782e8b58dd3f1e9e4276619e8603c5de34b4acac5;

            Ia36b5d24ca414ff96899820bbe3f5fc319b1e82dc558c2ec8af7559b6c45992e = Ice2f6ae40746fa0bd1c5b2db1aa0bac608899f3ec311d6e8459e126e446f7947 + ~Ic24e91afb654a0ee04d27daccc66b42d5e001a5962acd08aa73c3e962e1f2c88 + 1;
            I78f9a0c586ec95915e1628e57d58d38942d01562658ce91c4409571459bbda96 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia36b5d24ca414ff96899820bbe3f5fc319b1e82dc558c2ec8af7559b6c45992e);
            I48c21b6fc24c93dae3a01b55b280508297e0ff5101c7fbc7d17e823d9a31fb07    = I78f9a0c586ec95915e1628e57d58d38942d01562658ce91c4409571459bbda96;

            Ideabf29ace18ebaa3db078d782fa2d3b2db1422ddc35c86dbb12c94f172ac364 = Ice2f6ae40746fa0bd1c5b2db1aa0bac608899f3ec311d6e8459e126e446f7947 + ~I4408d142165f7f5bcee86e820e4ce79b4ecfe2134d8e50809080e0c27e4e2df9 + 1;
            I18c23544d10425853b73e8bd64411a829f4bd9fd145e5352cacd6ecf0c764945 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ideabf29ace18ebaa3db078d782fa2d3b2db1422ddc35c86dbb12c94f172ac364);
            I9d5c1ef1f35b4d40b4f20dcd2c33691152683bf308c95aa53adbf785defb75ef    = I18c23544d10425853b73e8bd64411a829f4bd9fd145e5352cacd6ecf0c764945;

            I82214920f75f46eb33a8b5e21ea60398b1c58a185ecc19b1ada4e7cb441e8773 = Ice2f6ae40746fa0bd1c5b2db1aa0bac608899f3ec311d6e8459e126e446f7947 + ~I3a210f2cb408bb61efba033b0ea8f1cda9a3341500248e1443840c24dfe04cea + 1;
            I5c79c03f571f276bfc03a16709012424498a1d7d53208213e600cd300cfddaf6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I82214920f75f46eb33a8b5e21ea60398b1c58a185ecc19b1ada4e7cb441e8773);
            Iec1baa5364573d0a9866494a039a3409a32b4665d4a79e2a729b54d370ecad97    = I5c79c03f571f276bfc03a16709012424498a1d7d53208213e600cd300cfddaf6;

            I193ddc6f5bac9d6f9e6599d78ec2c22aabe3032583f3dff87a62b3dca9074fa1 = I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec + ~Icf6cba7551eee2b4d2b53263af6fc190558f5b29af52c060adf5bc9116d56341 + 1;
            I2ce3e228247a767e41b5c376457e5be0d11aaef621b0d63d7683741f275b3f4e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I193ddc6f5bac9d6f9e6599d78ec2c22aabe3032583f3dff87a62b3dca9074fa1);
            I508c79d6f4d56ea0e8100825c438214e4b5087004f8a5041b4beb900509cfde8    = I2ce3e228247a767e41b5c376457e5be0d11aaef621b0d63d7683741f275b3f4e;

            I27be9ab07b6db7a211f0f2fc97fae8866b139ac8b76fb72d5b207866ef5dc538 = I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec + ~I5aff0a6c62deaff6e9d15280ae8c3cc326ae7f9ea6959dfa41a92c770b592cce + 1;
            Ie00142d305ce51cc78575481f10dda9c40010d6ae4a3fcb4435961983c8aa98c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I27be9ab07b6db7a211f0f2fc97fae8866b139ac8b76fb72d5b207866ef5dc538);
            Id55510ec558d15440325660ab2ac2cd9d4dd682c082479a742118c9ba1923cae    = Ie00142d305ce51cc78575481f10dda9c40010d6ae4a3fcb4435961983c8aa98c;

            I9c74de21b57f62df69930fb5dba0c0a81dcd57ea06cbcdd3e1dcbc9077a7396e = I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec + ~I6853348c8635a69100a45e6b2b255d6111daca84f2eb28629edd64f8c36f014c + 1;
            Ibd10325e424f3c8f0a460f2a4fe7bbffbfa3bc23e74abe4dfd6ec5b278e2c4be = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I9c74de21b57f62df69930fb5dba0c0a81dcd57ea06cbcdd3e1dcbc9077a7396e);
            I000c117a768755741005775b84eb6e4c406d2e29765ca9bbab991217963de8d2    = Ibd10325e424f3c8f0a460f2a4fe7bbffbfa3bc23e74abe4dfd6ec5b278e2c4be;

            I6a231da6c84868f89279c52b472159f3f28b097d98b55fa959cf8b65bd7357b7 = I4b20320f8be2127acc9ab378a4b87d242d1c8c041789919b7dbd706e7b4835ec + ~Ifd9d392bdf654a9146eebb9a670b75f4d74807786708350ceef7c79d54805ccc + 1;
            I47c4e3e3263c6533efa2dc2e7f1ec4150499e8360e38b1cfaa524071faadc4f5 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I6a231da6c84868f89279c52b472159f3f28b097d98b55fa959cf8b65bd7357b7);
            I95d510e99cd368229106d7ef60f9438bc186adb5359c9483b645b255a769df90    = I47c4e3e3263c6533efa2dc2e7f1ec4150499e8360e38b1cfaa524071faadc4f5;

            I2d28f08decf784d91ab2c0bb92cb9b95d798ec46ff319335f399bf55f24ca0c9 = I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8 + ~I9df56fb9c7b812f3ca5949962100efeb5889d69ff60754cb4eb3e0dd18376d45 + 1;
            Id2b48e805b3470041470bf0544dba31d75214a8834e8c456aebb8dc5a12e8656 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2d28f08decf784d91ab2c0bb92cb9b95d798ec46ff319335f399bf55f24ca0c9);
            I4cb9b54295972404ff2984e0b2a225773e067803925fc434674a5ef2439df4c3    = Id2b48e805b3470041470bf0544dba31d75214a8834e8c456aebb8dc5a12e8656;

            I2ce9a3e0eb6568348a715f3d26e23ff836ca88d2a48d62beb9b06f46ec986df3 = I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8 + ~I6c8cd97a5a950e00f0b9892a96d99ad1e5bae6c2db215bbb532060b753233aff + 1;
            I945dbc06fbc44959482d5670747fc5c6044a790ffc0a73ca0f41f150e8d59056 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2ce9a3e0eb6568348a715f3d26e23ff836ca88d2a48d62beb9b06f46ec986df3);
            Ied36baf05b90f7d785653eb1e7f699cfa84cd0a1eb3a985047f57e2885dad2ef    = I945dbc06fbc44959482d5670747fc5c6044a790ffc0a73ca0f41f150e8d59056;

            If13322a1bb24c2938298fda568b15f72bd6258fa12017507e5c8c34aa31969d9 = I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8 + ~Idd51d2eb571b7a35413e786a8a9437a5ef34a13b84d269e29c3319a4bb7531de + 1;
            I7d3a0a0dd3aea84fb203c8b51f1e4424f287b9ef01410f3cc5ac7e7579f2d4c0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If13322a1bb24c2938298fda568b15f72bd6258fa12017507e5c8c34aa31969d9);
            Id3947617c14deada0b43f71b47e700dbd8a1ac15820eed783d58774c249d5f24    = I7d3a0a0dd3aea84fb203c8b51f1e4424f287b9ef01410f3cc5ac7e7579f2d4c0;

            Ifb7752c1ee4d32c33015b0978e0bbc378b26a7467ea1c4983c2700f2372de3af = I8bda3b8333aea3c779a76564d604a3f7962fc7fb447ac140a1cab2a65e884fb8 + ~I3cf51d0ae95d4e3f7d0809785f84c5d25153742e5dd0d370235828d4f9c0d1cf + 1;
            I297e0d55dd6607cd32af52aac3e610ccf0fdb5e52f2ba250dd2c929616a33a8d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifb7752c1ee4d32c33015b0978e0bbc378b26a7467ea1c4983c2700f2372de3af);
            I846f9754b91cbdf37fc2662d5851bfffa4926c1ef01f4a23f20b02d9588ff3d4    = I297e0d55dd6607cd32af52aac3e610ccf0fdb5e52f2ba250dd2c929616a33a8d;

            I29cab53a69f72bbcf1812b364c9d4aca2dd9ca2159114ba63770ba7bf154c032 = Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421 + ~I5cbb1dce1049c737c8e052dd6b84121d353e3ee02202bcb8e5fa27261029c96d + 1;
            Id4d7fc501da443ac562b3578778aaea5dca1938dfb4563d14632481d1f453eb3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I29cab53a69f72bbcf1812b364c9d4aca2dd9ca2159114ba63770ba7bf154c032);
            I7485137b6eb30fbd6f06453139f9cd1ebeec411e566936bc598f0aefde881251    = Id4d7fc501da443ac562b3578778aaea5dca1938dfb4563d14632481d1f453eb3;

            I98b2432228e13880d555f5f32794fec8e0c4b85eb066e597f61dfae883cada43 = Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421 + ~I20a501f960ccd425135a3fcb8e667d68940a5950d939bca37d107d479984c038 + 1;
            I8aee3ea7ce652159455573562acaad5e41a877766e7fda11580be1d60194305d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I98b2432228e13880d555f5f32794fec8e0c4b85eb066e597f61dfae883cada43);
            I152ada5197e26088aadb2058a128099d201dc6e91d564b80b8e3930567a1a929    = I8aee3ea7ce652159455573562acaad5e41a877766e7fda11580be1d60194305d;

            I51bb519f0f46144969987729901cfa4e19f29f9703a5c2129ced5c6bf9c4531c = Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421 + ~I5c29250eb53f0eefc2332419b6c8e82f97741659657c08af97f8443954a5385f + 1;
            If787f037863d4eb15f1371255724977e8b67d17ffc783cb726ebec744a0ed62c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I51bb519f0f46144969987729901cfa4e19f29f9703a5c2129ced5c6bf9c4531c);
            Ic86eed327a12ce5bd475a6b82a5bdc31777526455fb541a8f4e842605bb34ddf    = If787f037863d4eb15f1371255724977e8b67d17ffc783cb726ebec744a0ed62c;

            I3865ea29a692b3a2567934ed101bc0dc34c941c7fa7c6fa6bd04a0670fea64c9 = Ie0b7e865d59f2c401a0c869f48b3fc7dcb7c938ef311f43b1006de1663017421 + ~I4fc7c4344699ed94536cb79d86f697e9da22498a2938b10360763aa9bad9da33 + 1;
            Iee4c52c7ebe29b796d3815def71a1869f8acb0bcdc109ad21b59ab2aa610c807 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3865ea29a692b3a2567934ed101bc0dc34c941c7fa7c6fa6bd04a0670fea64c9);
            Ic1a3e7a14eff1a6da9e96ddbd750086b011cdc44e8aa1189879b056fc48b3a27    = Iee4c52c7ebe29b796d3815def71a1869f8acb0bcdc109ad21b59ab2aa610c807;

            Ifc0ce7736e9c48c2d5e0e39ccf90c85218bd13a7e93695a158971e86e560a9b5 = I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e + ~I8d463b693ea969ef3023c411c0c9a1fbc49f81d348282c031b963bd8ce0527a3 + 1;
            I580713ee6afab29f13f6dbda18d77ae815138af729f981a455d34aca294bc4d3 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifc0ce7736e9c48c2d5e0e39ccf90c85218bd13a7e93695a158971e86e560a9b5);
            I215ee2b19d3ea96eedc62d8cb097051dad2d917dfb2eb2b0e1ed0ff697955765    = I580713ee6afab29f13f6dbda18d77ae815138af729f981a455d34aca294bc4d3;

            If5eeb2eea320a2012569a69de41e3e45dbf74bd9e8330a3c0a1b6fefc8994f01 = I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e + ~Iabd5561747d288862c0b289a28572fb5b0159a3fff7f79c59bf60f1612ec1e3f + 1;
            If18d826ce7582d4bf76e5968c9c86b08281682d30b790679e01e9aafa86f195c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If5eeb2eea320a2012569a69de41e3e45dbf74bd9e8330a3c0a1b6fefc8994f01);
            Ibbfd537ee459654bacd89b68f7d66565efcbdaa3838dc0847f83ba17c49b404b    = If18d826ce7582d4bf76e5968c9c86b08281682d30b790679e01e9aafa86f195c;

            Iacf07c5d8bc2563c377f66311c807d18c4cae1b4af253c3c55cb940c9d49257b = I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e + ~I4e6e6be5d9a7a85cc07a42c3a252e38fad4229a40bd68bec6728e7efa85984be + 1;
            Iff4ecb0f057c396e2e94c919920695cc67ad53f6b463c28baefee01ee00e4942 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iacf07c5d8bc2563c377f66311c807d18c4cae1b4af253c3c55cb940c9d49257b);
            Iccf845c102c65fc97a1244cb2c0182925c72e95fb4a9b0dc97379f5a32837612    = Iff4ecb0f057c396e2e94c919920695cc67ad53f6b463c28baefee01ee00e4942;

            I0c2168302de09a1bb09056d8e2f6cf9a4191a5151b99efe57fe8fec69e2c349c = I2d3ae3bd643723ef9b5bc0d3d4eee10916d64fdbf49fc42c50f3901e223f887e + ~If7b4cbde972a67fae839c5bc9ddfd64dc244041f6dd60f95c5329105ae08e460 + 1;
            Icb8d3dd7bb86ab8f1237c04d9d07d1d6046f07c618a3bd3308c59483260b7365 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0c2168302de09a1bb09056d8e2f6cf9a4191a5151b99efe57fe8fec69e2c349c);
            I32562e9f1cb6c7224d2efbd29f393e04c0d655e4bef402c2689cb946013f5d1f    = Icb8d3dd7bb86ab8f1237c04d9d07d1d6046f07c618a3bd3308c59483260b7365;

            I7aa29eeabf60e0de8e049cc83631713eecc92a33b00ab66889601b65a8584021 = Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf + ~I60b41ade4579462091cc59f1faf9f78f236a3bef12f893facebdf8e6b00096e7 + 1;
            I63450ac287a1e882703f7362bc499e7c779a7e68a1fbffd944aaf0e770fe18cb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7aa29eeabf60e0de8e049cc83631713eecc92a33b00ab66889601b65a8584021);
            I8ee1c7843334dc659003797fc7ec177037e184855e8e80063c6e490425de9446    = I63450ac287a1e882703f7362bc499e7c779a7e68a1fbffd944aaf0e770fe18cb;

            Ib7cd9e5a80b095f4c71eb6005d588f15ea498ecbf90748e128e42c0feee08dbe = Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf + ~Id73bbd3c91f1e5fe13f11e8849f77aad2ddaa35d1399140ceb5e133da8e11227 + 1;
            I1288c340fbff871d0fb4e5aab171e965bdf5b3b6cde30bb17f6a8d04ef546109 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib7cd9e5a80b095f4c71eb6005d588f15ea498ecbf90748e128e42c0feee08dbe);
            I5c6a9cfeb6a0354276fa86b65ea21b018e71d37b366f907012b41156aa22bfcb    = I1288c340fbff871d0fb4e5aab171e965bdf5b3b6cde30bb17f6a8d04ef546109;

            Ia9f187fb62e136eb42c8ab963813a504fbd8ed5f7390f608f923c3d5f8853a05 = Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf + ~I8a3b07f660ad94b304ffecabf47d3378d3ea73b1deccd771fd1982cec9f23e39 + 1;
            I559a54fedbda0d961279ffb3fc4d2eb644cf2b77f805acdfde54df03ba0c05f6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ia9f187fb62e136eb42c8ab963813a504fbd8ed5f7390f608f923c3d5f8853a05);
            I76041755b112a333460289875673d3f2b054918770d3a2cc46ab7a9f92b50eb5    = I559a54fedbda0d961279ffb3fc4d2eb644cf2b77f805acdfde54df03ba0c05f6;

            I482ab667b97b8e90796abc13f93d317377f279dcbd4c9699b5bf776cca58e12d = Ib6b661dd44e03bf1e3321c1c963e35e7f334f000eca05acfd994f33b86de8cbf + ~Icf608ba43019dffad0c708d49076088f2a4b5e126e76b3b2fefa5a0f1edeac7b + 1;
            I628a71f11553d99c7d0f19a7932ab7250a9448868d3e118479c70d70e1481ecb = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I482ab667b97b8e90796abc13f93d317377f279dcbd4c9699b5bf776cca58e12d);
            I30843beae9ebf34c0f73f773e1af0422e40b3ced201574b6f87f400cb37a7175    = I628a71f11553d99c7d0f19a7932ab7250a9448868d3e118479c70d70e1481ecb;

            Ic59104908c4c5eb1da72d1f877270cc3a75512d885653de8de2aaa5bc050ae87 = I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2 + ~I8060bc4cf825f705f2218152b6a7a8600692076ba01123cae35feec231f128dc + 1;
            If06e126d9560577dd7525491f2092e8e9c9ff9e64c0ef94b3d0ca2b61cb6392c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic59104908c4c5eb1da72d1f877270cc3a75512d885653de8de2aaa5bc050ae87);
            I7f99ba04346760d4ee2589662be79b19673e741f07d1b9c0c35b54d4bcd3cfc0    = If06e126d9560577dd7525491f2092e8e9c9ff9e64c0ef94b3d0ca2b61cb6392c;

            I2e28e3dc68c6c9d929ff4706e92b74d5b52de590d44dc846007d24a929cb60c9 = I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2 + ~I47b18bf83ed7f7e8a2c69814aafa41a66b6838a5a997d036c634f488f1c584f1 + 1;
            I42760d09b067c76aa603d685d09ef8a3fb0aeeeef30a19648ab2cc69233d8514 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I2e28e3dc68c6c9d929ff4706e92b74d5b52de590d44dc846007d24a929cb60c9);
            I311c88c2854536dbb8f578bdf98823eaf5888a7c772bc2c6f0cb49c9c9c79500    = I42760d09b067c76aa603d685d09ef8a3fb0aeeeef30a19648ab2cc69233d8514;

            I29c2a83008b667730e3fa038ef10d5c8c989348c36320071fe5a93d15a608d65 = I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2 + ~I55d6bfb606269d9d01dc348f732caf9cfdc7042c845744b7a25c0a74d0afefbe + 1;
            Iba06a153040bdb18311bb9c6826eddd28863470c44a75683bff1dbb5d03e1d39 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I29c2a83008b667730e3fa038ef10d5c8c989348c36320071fe5a93d15a608d65);
            I073f480ce57215d8a9930ab34bbed6bcf5e631613fced0e782749a390615672c    = Iba06a153040bdb18311bb9c6826eddd28863470c44a75683bff1dbb5d03e1d39;

            I7e9eb2043321328a9ced3e4d319e6963e60ba7928bec6115527f55f70cbb8db1 = I2c269a80fd6c291845bf9e97764622597ab62ea5c454022f07b532ff8a8d7dc2 + ~I0a5867bf6971ed11db3a6dc9af8cb356352990bbc3032878e82b6cb2ca8c402b + 1;
            Ifa64872cb59e066ea755fd8d50aa1fbdf10fbe3920e9ccbbad20c899f377207b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I7e9eb2043321328a9ced3e4d319e6963e60ba7928bec6115527f55f70cbb8db1);
            Iaef86ab80a38f09821c64eb7b93cf066c0ba40a4b315075fd4652eb82b687bff    = Ifa64872cb59e066ea755fd8d50aa1fbdf10fbe3920e9ccbbad20c899f377207b;

            If70d53608aa2878766b77726f3e0f650f572b7e89ea4df1a4504306868cc44be = I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987 + ~I8090d844610f0d62cc25a9c72c2d76d9d6783a067de9c9ea9d5a1f5c48744c70 + 1;
            Icc225eef673a329e451a89e36893eee8b9d8d9b8cfc911d6bf84a2ecafea5e4e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If70d53608aa2878766b77726f3e0f650f572b7e89ea4df1a4504306868cc44be);
            Id523ce79d9f7a6b24c5979c58855211eb2bde238c81e549064c23ec62a5c7a3d    = Icc225eef673a329e451a89e36893eee8b9d8d9b8cfc911d6bf84a2ecafea5e4e;

            Ifb7ec2a54d000887851d37b4b0f1be483d3caef91a4d07b19edbc19995fc77c4 = I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987 + ~I79d13cc47977ecb1fb0ca304be8c225a427063b4328cea4c4a227521a1f26018 + 1;
            I3bbfc044ed936cf51599cd8977c7bf894621c83e1e73c4cea372dc54a1d6c028 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifb7ec2a54d000887851d37b4b0f1be483d3caef91a4d07b19edbc19995fc77c4);
            Id27c2a1647e08c46fba102b41eceb3513a697df9876d76b23fc4118f16b479a0    = I3bbfc044ed936cf51599cd8977c7bf894621c83e1e73c4cea372dc54a1d6c028;

            Ib24004e855a53de1330e5ec4126e220205ba20169ae9ee4ec34135db389763bc = I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987 + ~Ic3f066b6b8dc09e89e9796c2b739b37e64af709758029ee21800f9fdf02c533d + 1;
            I809ac54f05fda9abf4917b1e555505f9eb41cf89a9a9fa098fd642e90bb635b0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib24004e855a53de1330e5ec4126e220205ba20169ae9ee4ec34135db389763bc);
            I54a09dd4115c1f70cff7fd7921120216494997fbc08a7e9eb8e59152ef12a9e6    = I809ac54f05fda9abf4917b1e555505f9eb41cf89a9a9fa098fd642e90bb635b0;

            If81c09fd3901cbccd2410864fc3e2d7087c400fab7cb319f6de0e030d706dc1b = I0faf7efe7eee34921c3aede5f7f6ae6f17639080bd6e9e4bc61595a59ad9f987 + ~I56253c88487a75fb5f830a66c0dd3172ff25795a2509eaf5367fe045f9e12b61 + 1;
            I3435109d555534fce5a4cccb9709c25bb5ea401158c144add8e4c09a6a68c8f6 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If81c09fd3901cbccd2410864fc3e2d7087c400fab7cb319f6de0e030d706dc1b);
            I5a2063e62c2c96b172ecad9fa950c0b42c413214e30d94796ca9c2b8c6bbe522    = I3435109d555534fce5a4cccb9709c25bb5ea401158c144add8e4c09a6a68c8f6;

            I3ec9f20d41034d8e73b2a9210188b70e7b2c68e62b25fcb5f140598043681a6a = Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3 + ~I799968e729d7842ce09a838203458d89b96fe9d2d7a5de0cbac32eefbf834898 + 1;
            I0fc48ba2f5bdf67aabf15071712eabd08121ca31614dbbfb3ce3eb7cf6287364 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3ec9f20d41034d8e73b2a9210188b70e7b2c68e62b25fcb5f140598043681a6a);
            If0c2c0785586996991da246fc01722deded4e3ca8550290626324c5908d770a5    = I0fc48ba2f5bdf67aabf15071712eabd08121ca31614dbbfb3ce3eb7cf6287364;

            I21d1d0816fb6a0c22f2e850ac9a2d9d1f582c218de0eae741d1c9916ad2bc5f9 = Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3 + ~I02962ee90b42f9b95262049bd2dcb7da2f43333787a578d5f5721681773db287 + 1;
            I36a6b8814b16f2a3e44bf1afffac6416088645e41a495b7dcf9053020718e983 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I21d1d0816fb6a0c22f2e850ac9a2d9d1f582c218de0eae741d1c9916ad2bc5f9);
            Icb2218fe2214af22ea6fff2b9ff3c8d1772fd9318efa83c7655b0dfee2f6ab4d    = I36a6b8814b16f2a3e44bf1afffac6416088645e41a495b7dcf9053020718e983;

            Iedde649e1098e7cafbda605e624786ca97ff3b6e68c7ee8be00b813d8ba5521a = Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3 + ~Ib36374f40465c181d1b8d65f23001a10ffaa250f0fd89077848e6a49a19c56dd + 1;
            Ibbfffde74fd960499ea7e7ce9dbd03e057746dd164bc9af0e585839225056f42 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iedde649e1098e7cafbda605e624786ca97ff3b6e68c7ee8be00b813d8ba5521a);
            I0c567cd54c6fded476f507a4a35d7d93fdbd2cd1c555e10edf313ddaf4b0d64f    = Ibbfffde74fd960499ea7e7ce9dbd03e057746dd164bc9af0e585839225056f42;

            Iee58ae84679865c9bfa421865961b359874636d1a9a6a85bda680627cf00cd2f = Idaf5e3fb95864b6c6a8fda88e35992ccda5287549564966df082eddd405a4cf3 + ~I199abcfe7a0dfbaa58ab1dbbb16223bd434b4ce5ed3a65633d506d668aa76f8c + 1;
            I0cfea5b22889a1b983f14e6d1c3bd847f20dd9cd96b0cafe80e1705be750eb96 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iee58ae84679865c9bfa421865961b359874636d1a9a6a85bda680627cf00cd2f);
            Ic49fb172f5523a522e94efd83b5827b8f63c2d8fd7c76263249d96a00a0e25ad    = I0cfea5b22889a1b983f14e6d1c3bd847f20dd9cd96b0cafe80e1705be750eb96;

            I00a07c03491a1f197d8ff004b3a7816850d0cd272e4ab9dd574ed104f730500a = I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96 + ~Ib1101385e86160606eeb12ff49ee86ca465f227b19c9bcad4811c6a0183c0ddc + 1;
            If34a395225bfb809ae5327b364a127aec5b1e5ef9e4fc9bad4baaa13cf13f661 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I00a07c03491a1f197d8ff004b3a7816850d0cd272e4ab9dd574ed104f730500a);
            Ibef81155a593cc991eb8f0da7ea8dbc27f3c935dc1fdf7b857110407ef449718    = If34a395225bfb809ae5327b364a127aec5b1e5ef9e4fc9bad4baaa13cf13f661;

            I0fa68b59aa1d936947137ecb31171e019a59aeadc82044e25faf04536b89d301 = I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96 + ~I44445d003eed631dd6933d4ade176469fe9a4ef0b21b0ee20067b5aae73704d8 + 1;
            I31edc2dea3cdd499a9a2035d2460448786e5a44b1d828d6486d7c3ccb959892b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0fa68b59aa1d936947137ecb31171e019a59aeadc82044e25faf04536b89d301);
            Id1c35604f896316440f1deadc55ea39d16307edf0e2ddea1d7d450c41dbbc705    = I31edc2dea3cdd499a9a2035d2460448786e5a44b1d828d6486d7c3ccb959892b;

            I4e3ea3d10bfb18320ffcdf21e5b7f279ab94cada35ceb624c8bbb1f5fed062ae = I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96 + ~I7c843a280d8a673e3c59a22f8bfbd5860c3284b189ffa281759aa44233eee225 + 1;
            I31d6cdf7439ddccefec7a19dfdc442d351d609dca8f14aa276c22741a45aecee = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4e3ea3d10bfb18320ffcdf21e5b7f279ab94cada35ceb624c8bbb1f5fed062ae);
            Ic00c95647ac3595e199e62c4d3e75956755ac952e4cea464b27066ad8f09415f    = I31d6cdf7439ddccefec7a19dfdc442d351d609dca8f14aa276c22741a45aecee;

            I37b48c08b0e188a8ae4c35cbe94bedbc2be0d8ccfe5dc8199fab4bf3a5c2b4c2 = I4c7ec78b196a19f74203005d69f4492537f9c9f6fa251d27b45ff0c0ba21de96 + ~I2ff52a8e46c22b626ca488ae87c88360d413ad08dfaa6701fe7b237d42c2cbe7 + 1;
            I2b2cba74c6c9eeade51d69171bf22d1de38947948b7af485a5e64aa9bd90d71a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I37b48c08b0e188a8ae4c35cbe94bedbc2be0d8ccfe5dc8199fab4bf3a5c2b4c2);
            I4d89a637472e8c4d071c44792883afdac1fe1c6ffa9d08f7259525884000b34e    = I2b2cba74c6c9eeade51d69171bf22d1de38947948b7af485a5e64aa9bd90d71a;

            I311137155e974b61171f0b9f85b3380cf230186a137daeece322108026a54fb4 = Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d + ~I52cf6523f0dd5f666334b2646768fe4499c699c8f6b27ec32ae325cc0981a515 + 1;
            I45a1490302e61b9172caa0feb0aea621e97a5a95b9e8c525d3ad875898955f02 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I311137155e974b61171f0b9f85b3380cf230186a137daeece322108026a54fb4);
            I081fd1385ec974da04b64bc5764efd6db252fefa40f518ed0ed4b01ce630064a    = I45a1490302e61b9172caa0feb0aea621e97a5a95b9e8c525d3ad875898955f02;

            I86d7cfde239760ee206e636d19402cb5decc9d170670b47874bb6e51950e797a = Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d + ~I289b4317d3472843dd49dc75a39395f8c39b9fc0c70000205510d08404d824a3 + 1;
            Ie22f10e98c9847ef82cfedf9cf3ca17fc0307139848522f58fe0ab8f92d253c2 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I86d7cfde239760ee206e636d19402cb5decc9d170670b47874bb6e51950e797a);
            I57c394b657ecd32691fcef200ba361abaffca7d8ddbc7bea22502a9f7bff9f5f    = Ie22f10e98c9847ef82cfedf9cf3ca17fc0307139848522f58fe0ab8f92d253c2;

            Icce39cddc9b07a5408d7b7cc73a0aee0ba96dd9b59ccb5f9da245a8115636e81 = Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d + ~I5eef24c8de2049e0e8bdd49346b6be22708a135d56c096907e50ecfbf3affdea + 1;
            Ia40a2c6be098446003dc0b6caccdf75cd1ecce9fac58135f83551b0029ef7032 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Icce39cddc9b07a5408d7b7cc73a0aee0ba96dd9b59ccb5f9da245a8115636e81);
            Ia14c31a81641330844c0c48e155c6f7630695ccf3e7238ad6eca01c8a45a104e    = Ia40a2c6be098446003dc0b6caccdf75cd1ecce9fac58135f83551b0029ef7032;

            If0c116c5bb5aa35db83ca1f71a49e32a260c13ce39a02cf3b683d3cebcdd412e = Ide8add98fb8e5ade41afcf207baba9c671e59b0a24f6e720bc116deaefa9217d + ~Ide088b881c7dabf6e2fab61eb4e5db3ea3750d7b72eb26cb79877bc23429efbe + 1;
            Ifcdbddb54d9293f008a7bf068e7733c4ce75f38ee2cbe8ab4247bc4200a604ac = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(If0c116c5bb5aa35db83ca1f71a49e32a260c13ce39a02cf3b683d3cebcdd412e);
            Iffdff1b757352d5f1174deb338f337fd8841ce8d132c2e0a16f18fc1a97313a2    = Ifcdbddb54d9293f008a7bf068e7733c4ce75f38ee2cbe8ab4247bc4200a604ac;

            Ibc1d7004fdb14267759bb0b179acbaf24853d6b0efe051dfd48de07495940dca = I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a + ~I3e5c11a25b8726c787dd0ffc08e93b671baf84832d9413eb7031a6fc17e8ad76 + 1;
            Icc54d76cca75160c97db719151bb55f2d112201e3812c72f002b3dba5e61575e = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibc1d7004fdb14267759bb0b179acbaf24853d6b0efe051dfd48de07495940dca);
            If8c3dafd18d6fabac3e4ec4dce257aba397ab0d341e25a1bb88f9e32909deb17    = Icc54d76cca75160c97db719151bb55f2d112201e3812c72f002b3dba5e61575e;

            Ib01b562cc42dd79d910091cbfd3ecb8cd0b386f396893baaee60076b8c04f906 = I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a + ~I2e063205340c315025edf32a4ba91e5f7cd39f37fc5800906a3862780cdf7d9a + 1;
            Id2df947b4126f71a866a204090780296b99e4ca990d0d27c7e3750ffb4d11451 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib01b562cc42dd79d910091cbfd3ecb8cd0b386f396893baaee60076b8c04f906);
            Ie4b741e2c3f5dbd43bba89fbaeb4cc6b309042b53629f8db67121eb22a656ee9    = Id2df947b4126f71a866a204090780296b99e4ca990d0d27c7e3750ffb4d11451;

            Ib1b3ee65ad4ddc6d66bedc912f129d315715913cb1517e24bfec0669f2b3ea04 = I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a + ~I29141cb56b9f52d74c42d689b180cfcfe7daf23ce573c1f4eaf21525370e5376 + 1;
            I8601156c6a18f07b4580760c232a62262c2eb8d656282d9710517b6bdb886459 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ib1b3ee65ad4ddc6d66bedc912f129d315715913cb1517e24bfec0669f2b3ea04);
            Ib1a3877a6c9f5b87fd3c2104782a0699748b68ef73a12291b34e914344db9d25    = I8601156c6a18f07b4580760c232a62262c2eb8d656282d9710517b6bdb886459;

            Ic2d2abe362d0a76e22e5bf3d902cf55d1091dce5ff18a17ec2b51dac09d2601d = I2634a7facad5d227f558bfebd58ecb90b4bf24d1adc41f06fdbab9364393aa8a + ~I5df56a6a00d4d8ca1c6b1a79e5f0e674482cb9541d86dd49c2ac361d86dcea1a + 1;
            I19e014466929e7ddd8d4a2a3f0fc6cb3d9eec8d39e8f7a81458043ccaaa90ee9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic2d2abe362d0a76e22e5bf3d902cf55d1091dce5ff18a17ec2b51dac09d2601d);
            Ieab221c067f0649e88f307dd8c46981653088853874e2a256b99f7b7a8bf93d5    = I19e014466929e7ddd8d4a2a3f0fc6cb3d9eec8d39e8f7a81458043ccaaa90ee9;

            Ic667337f6e8f713aef676104d2c4af6a634660e47835d615bb7b74af34c3e979 = I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df + ~Ic2bb8293812351030940ea0e0a882994714d60a4963e82e2291f6f2d386fce8e + 1;
            Ia24a2450394a5e7953feb8631095648c20bd71240699f481a0c3b748e665aa64 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic667337f6e8f713aef676104d2c4af6a634660e47835d615bb7b74af34c3e979);
            Ic80161feee5be9576086dd9d1ed8adca369a841f0052af01b2fe93d46af669b2    = Ia24a2450394a5e7953feb8631095648c20bd71240699f481a0c3b748e665aa64;

            Ic0a75ab618b9081cfdcd40620ad47ce4da348de800f33a88cae7bcee7ec46f3a = I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df + ~Ide8930fe855e6fb7dd5b689395a121a16f491421d448454c9c021f62753732c0 + 1;
            I5434f08cd24b915586080bec92103df0eb2a3d6d14ee496326046918db03b549 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic0a75ab618b9081cfdcd40620ad47ce4da348de800f33a88cae7bcee7ec46f3a);
            Iac4628a0a7bdc975990c2664a736112cdb2bf1b1b30f89ae1e6827a44bdb4474    = I5434f08cd24b915586080bec92103df0eb2a3d6d14ee496326046918db03b549;

            Ie6e50cae460faffae965f9ee7bcde9b12d5efb54a7d8f03d45a34cd1cf6e36d7 = I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df + ~I405b2f517ad52ec3c94eb9d1d695f6fb9700fbd32fb49fca23588911b5dd0ef5 + 1;
            I536c65ee87da658790b4273c04e7acefaa2baef5da84d48a9a53686c9ad20195 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie6e50cae460faffae965f9ee7bcde9b12d5efb54a7d8f03d45a34cd1cf6e36d7);
            I7da6920e7bb85e837e61b04ba09453237164470bf2eb7607af94194e05407bfe    = I536c65ee87da658790b4273c04e7acefaa2baef5da84d48a9a53686c9ad20195;

            Iac4ccc031aca350afe26f7ca6b09c8d4c124dbec5e0e705ba473f4c2834952f9 = I51fba9288b79659d99c3629d7356edc73dd5bc9c61c0ec58fbc9e4283717c2df + ~I16b3b3cdfef91e9cd5ab763bbcbe2188e61f45183118f5c735eff60965fe4138 + 1;
            I5ec53ebfd7533177d3d5a1d97e18c9e5f90e4caad316088f62d8bd0ec6bc983a = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iac4ccc031aca350afe26f7ca6b09c8d4c124dbec5e0e705ba473f4c2834952f9);
            Ie3ca82b8d601f023d408833c7b5445539ebf8f17bb678e486fb3f650b2e01d9d    = I5ec53ebfd7533177d3d5a1d97e18c9e5f90e4caad316088f62d8bd0ec6bc983a;

            Iedc1f868c50438002a4d97e96e0dac521014321ddc6d61e49b5eab223b997086 = Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481 + ~Ib4d2bee91a2ab56208d3d1f484e63f085a162ab9d482690dd3c5891a2a34d808 + 1;
            I1090417ca7c539e5bb1077d4b96824cac49fc6bd3253fb6d0348ec13edb97d2d = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Iedc1f868c50438002a4d97e96e0dac521014321ddc6d61e49b5eab223b997086);
            Ifc8ba6aad04e3418146443a14c520552e32ac2f43fabe430ef0d640b4262337e    = I1090417ca7c539e5bb1077d4b96824cac49fc6bd3253fb6d0348ec13edb97d2d;

            I18cd7259e4f753e93903dc1031fc51c25f000a37959e858574b79394f1dff508 = Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481 + ~Ia4205a1d01cb014ebf8e1d539dbe1c7270bf9bfa8eb7920b136417bdfb9f498e + 1;
            Ida31fcf4f48fdc3b391ca3e4d2c7b1c3ff6ce6ee53c2dfbbe1bc863514845a19 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I18cd7259e4f753e93903dc1031fc51c25f000a37959e858574b79394f1dff508);
            If1aa1bf1d7206ef9c00f8c1aafd738c03603858f9757a3f671242af1b139cc64    = Ida31fcf4f48fdc3b391ca3e4d2c7b1c3ff6ce6ee53c2dfbbe1bc863514845a19;

            Ie9395076cd1821b1a6cd391c4ce616cdbb0bc759a2a9f3a7ba32ec60b9c6015e = Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481 + ~I0bafe9c7cb10e6696f6b6dafb74a2113145f7ef1cb70496d068a61ba1de1bea1 + 1;
            I5b4f25d6b0cdd33c4b4f5f200eb9ca9d2ad68b01b48f7697100305c1456f35af = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ie9395076cd1821b1a6cd391c4ce616cdbb0bc759a2a9f3a7ba32ec60b9c6015e);
            I97205d95f7ff115112b2b1a7eb32bf70ff7c1e2fb431785547ed7f98d5fea0af    = I5b4f25d6b0cdd33c4b4f5f200eb9ca9d2ad68b01b48f7697100305c1456f35af;

            Ic30aa34e60dfa155b665def463cf115fe22112f358895a836b4179f33160134d = Iead0f188fe241b3a0ca8aed9e90c2e39bf6a7927468a47ea137d4a7d72c05481 + ~I78e49a2727c2f25a14e0f8937e6241f54246c8f42a643dc569f0249384909fb1 + 1;
            Ic98f738736b6b689361d5a77495e45e51874de01c86f1e7c10fe07e2c0f3ae82 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic30aa34e60dfa155b665def463cf115fe22112f358895a836b4179f33160134d);
            Ia6232cf34275276641c494e4f4cbd7a8796f1f946733ed0fe15d9e11cd8c740f    = Ic98f738736b6b689361d5a77495e45e51874de01c86f1e7c10fe07e2c0f3ae82;

            I577e72330edc830f5735c0ed269566f49c7fb3c4d196d3742fd1cf3c66cfcc95 = I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0 + ~I6822ca486e86051ea654b41b63bfefc12a2218ec87a88d8b5acc3e3c8a604c94 + 1;
            I347c2eca1405d163956cbc4ba007b08ae0a0a751bee7ecde367e2336fa308e26 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I577e72330edc830f5735c0ed269566f49c7fb3c4d196d3742fd1cf3c66cfcc95);
            I24883a74ba0e0eaf8efff93301dd4d714667c28020ff65d73e4056b2d014e287    = I347c2eca1405d163956cbc4ba007b08ae0a0a751bee7ecde367e2336fa308e26;

            I08b93985c2d4ce016468d10b7f0187ec3cd8a803308f2333bd361255e00977b6 = I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0 + ~If6fe8b42d897a8c92c628edac7869deee179622fa52fa779f2d9a0279791afc0 + 1;
            Ie0fdeb73844872fe9e7af165cda8d1c865df24e572180803760f4959f8e73ef0 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I08b93985c2d4ce016468d10b7f0187ec3cd8a803308f2333bd361255e00977b6);
            Ibdd97caada239a1152f2155c8cb9e25402600931810f6bafe34159894246d962    = Ie0fdeb73844872fe9e7af165cda8d1c865df24e572180803760f4959f8e73ef0;

            Idf041d85612e43dacf84491d005b30e93873e31c1b6e56df2e0ca7f0babdc5a6 = I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0 + ~I5b2b2323ba78f198e4c86b284772fed82ae708af1da14bfdf215a7b34f811204 + 1;
            I69baa1c18df6858ab86b75bb25b5f980db3508a861fc7da408a38ed95c910b16 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Idf041d85612e43dacf84491d005b30e93873e31c1b6e56df2e0ca7f0babdc5a6);
            I4ba3a78d1129b6b95ec4421b8dc75b90921b67ed09cc636c1fe08c778c9a4c87    = I69baa1c18df6858ab86b75bb25b5f980db3508a861fc7da408a38ed95c910b16;

            Ic9eb7815de9b84b1a3763dbf218de5d7d844ca252937b7685b20015bad378659 = I207a1ac11ab0cef656b0683d46a88f1b35052c55453db5a93d19f82aee01cba0 + ~I6563fc7a6bd595720441778baa975487126f50343c92ccba99218e274cf40336 + 1;
            I877a8619724696e16819de80d99f77e7ec18579f9e3cd99092f4ac0d358ab35c = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ic9eb7815de9b84b1a3763dbf218de5d7d844ca252937b7685b20015bad378659);
            Ia8fe4e59fc4b364c711cdef5a6718ae33543de2e35744d9cda4cf33f340d7add    = I877a8619724696e16819de80d99f77e7ec18579f9e3cd99092f4ac0d358ab35c;

            Ifa413778a53ec09ef3948f1ff255ab5b73d9243508614c057c59a153ad5289ea = I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219 + ~I01a734e70411ca4d260541915dfb0aa0eccbb88be6043a4a46e412d3b9f1e778 + 1;
            I97f8ce585d26cb40e221f7f8bff17e80cd5565540b9108ef64628053a3d547fa = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ifa413778a53ec09ef3948f1ff255ab5b73d9243508614c057c59a153ad5289ea);
            Ib0319b3fbdfab7c4df3ba7c1d710d7ca176cf8cd4223ea11fe12102cb5ac7f12    = I97f8ce585d26cb40e221f7f8bff17e80cd5565540b9108ef64628053a3d547fa;

            Ibc8a3b5a652d7343e1696747ac66770452a464ae8bbdd112799540acd80824d8 = I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219 + ~Ice95c4df972e8e6a31901269a2d291a70fe4e8dd1d86ea5ded5a16cb1c169890 + 1;
            Ibef17646fe9cd45fe72647539df79962a2f02d56819071f9e7740a099175decd = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibc8a3b5a652d7343e1696747ac66770452a464ae8bbdd112799540acd80824d8);
            Ice9d3685b31919d1cfe76a96ac6e1738ef6c66e069de55830f61665cb5bc0ca2    = Ibef17646fe9cd45fe72647539df79962a2f02d56819071f9e7740a099175decd;

            I3e50387897ad4d501a045ec8c1ed398fd84ff960cca94f41bd41fcd6462783bb = I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219 + ~I4a55baee8cbea583890824bd3ab4c4391b9d44203332575c030077c6e0e9f862 + 1;
            Ic2f933f79277b6967efca4d861031734f157410c96568f6370436fa3c94443d9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I3e50387897ad4d501a045ec8c1ed398fd84ff960cca94f41bd41fcd6462783bb);
            I36a3a77efd095e4c91274958f1ed4b9fc929f2b6794e4b879b8275f3a01ae48c    = Ic2f933f79277b6967efca4d861031734f157410c96568f6370436fa3c94443d9;

            I25ddd61dbf2b3f1b4024d769f62e690493ca0fdd01b3550226c9661ed9230fe1 = I39437fdaae54b8d3aec141f3a5d371da426bf8ec87ad02a2efe1f37bf11e3219 + ~Idc94a4d308c2e301c3d3524f1e20817f9b666827f340874b5adc763970f2efdc + 1;
            I34e2e324da2cf6bd7804e6c3d9a2e8af1ca0799f9a15e7c9597f812ee6679831 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I25ddd61dbf2b3f1b4024d769f62e690493ca0fdd01b3550226c9661ed9230fe1);
            I0643791cd1c7ee5c205da45ee4720229c6f7b61e98a7f642afc47506f6e10210    = I34e2e324da2cf6bd7804e6c3d9a2e8af1ca0799f9a15e7c9597f812ee6679831;

            I4dee2f1c5fecf86cc83b723fe96caccffdc564334698e43f9c04db5a25afc978 = Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884 + ~I93f4f945a6dfc45c0a002e0bd9251f56c68570c71e862e222a853f8855fb1165 + 1;
            I0784dbf1fd934c864e5c23e58e5636d5e4e72af359af2dc3cc1c11653a96d26b = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I4dee2f1c5fecf86cc83b723fe96caccffdc564334698e43f9c04db5a25afc978);
            I485c81ca3402c9b70ad8a10b749c0ee5e81569d1a64231a5fb25e3af8cc4abba    = I0784dbf1fd934c864e5c23e58e5636d5e4e72af359af2dc3cc1c11653a96d26b;

            Ibdf4b745b03013632bc0ac5142c9dfb98f197c78e95b71ce1074f84a5b5c96b4 = Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884 + ~Ie28b77da5cb0eae41811ec7dbc5f86111d64b794121eda9f2f0515324579f844 + 1;
            I1e024678e8d8668a4b3744b819e48699d59c21dd2856723a6af255d20bd83297 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(Ibdf4b745b03013632bc0ac5142c9dfb98f197c78e95b71ce1074f84a5b5c96b4);
            Ief695bef8a02a4f5e89c14ac6b89f84678cc7d7a9d71bf2a5e3c1abd44d1cbb2    = I1e024678e8d8668a4b3744b819e48699d59c21dd2856723a6af255d20bd83297;

            I0adfd7bea27acb0ef24fc07bb0649de5bc0ce7dca6226beef48e27cea9aa4df0 = Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884 + ~Iab63efeaac16bfc91c71a1a0819747c4576111221b2e355300a6e02adddb1aad + 1;
            Idadca14723005bf0db40379151927d667247f30071db43f735c3395db88dd110 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I0adfd7bea27acb0ef24fc07bb0649de5bc0ce7dca6226beef48e27cea9aa4df0);
            I0ce015383446aeba50b7677c9060a1e18dab91eb8040a718fcb7e104a700c29b    = Idadca14723005bf0db40379151927d667247f30071db43f735c3395db88dd110;

            I870372f2d3e9fcc2db983123cb83c7a6f1b5e9f022d915d5534425322e8957a8 = Ic0f894ce6262241ecffd6368658fc0ff6ffdc2566402a11ac08bd81afb590884 + ~I3167835472a3c4db7f1b7fbc1895c44e547122e9ad273066e6bdd43bccde11cb + 1;
            I0f94b265dac20d93ad623db13d43a951cd09643250c48e9d8f58e163ebb406c9 = Ie231944bb56504afd4cd4f051945212293ae680bfa7f185d00769b77d1dd196f(I870372f2d3e9fcc2db983123cb83c7a6f1b5e9f022d915d5534425322e8957a8);
            I9f790cf09f0d8b1c047cd0df401052898d374d930d5ccd784d142c544d8b54b6    = I0f94b265dac20d93ad623db13d43a951cd09643250c48e9d8f58e163ebb406c9;
end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
              Idd909220a9540c998e23f1b06cfca187d9d83bc0673aeafbd0ed6c20c9d39f4d <= {(SUM_LEN){1'b0}};
       end else begin
           if (I6d0b0c1a3968ec36626f19660bedfe0a538a7835edd2a21dd3f4ce0fe2c5c86b) begin
              if (Id76ecc370ac753fefd8cbdfb525a5868396234d646214915a49d70ad4cf925a7 <= HamDist_sum_mm) begin
                  Idd909220a9540c998e23f1b06cfca187d9d83bc0673aeafbd0ed6c20c9d39f4d <= Idd909220a9540c998e23f1b06cfca187d9d83bc0673aeafbd0ed6c20c9d39f4d + 1;
              end
           end
           else if (start_dec) begin
                  Idd909220a9540c998e23f1b06cfca187d9d83bc0673aeafbd0ed6c20c9d39f4d <= {(SUM_LEN){1'b0}};
           end
       end
   end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 I93c1856af28a13c1890271dc68b7b6cae884657bece4e0d452fce3ef922a9c12 <= 'h0;
       end else begin
          if (I47e3e3ab4fcba3cc4478ddd5e0ff92bb41fc8fb0403411b2b588ca51686b978d) begin
             if (HamDist_loop == 0)
                 I93c1856af28a13c1890271dc68b7b6cae884657bece4e0d452fce3ef922a9c12 <= HamDist_sum_mm;
             else
                 I93c1856af28a13c1890271dc68b7b6cae884657bece4e0d452fce3ef922a9c12 <= Iba7e42dfe0894a09d968f0190d344d90387e96a8048a01fbb5d05c15452f6ce3;
          end
       end
   end

   always_comb Iba7e42dfe0894a09d968f0190d344d90387e96a8048a01fbb5d05c15452f6ce3 = ((I93c1856af28a13c1890271dc68b7b6cae884657bece4e0d452fce3ef922a9c12 * HamDist_iir1 + HamDist_sum_mm *HamDist_iir2 + HamDist_iir3));



   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 Id76ecc370ac753fefd8cbdfb525a5868396234d646214915a49d70ad4cf925a7 <= {(SUM_LEN){1'b0}};
       end else begin
          if (I47e3e3ab4fcba3cc4478ddd5e0ff92bb41fc8fb0403411b2b588ca51686b978d) begin
             if (HamDist_loop == 0)
                 Id76ecc370ac753fefd8cbdfb525a5868396234d646214915a49d70ad4cf925a7 <= {(SUM_LEN){1'b0}};
             else
                 Id76ecc370ac753fefd8cbdfb525a5868396234d646214915a49d70ad4cf925a7 <= HamDist_sum_mm;
          end
       end
   end





   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          converged_loops_ended <= 1'b0;
          converged_pass_fail <= 1'b0;
       end else begin
          if (start_dec) begin
               converged_loops_ended <= 1'b0;
               converged_pass_fail <= 1'b0;
          end else begin
               if (Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e) begin
                       if (
                         (HamDist_sum_mm*100 > I93c1856af28a13c1890271dc68b7b6cae884657bece4e0d452fce3ef922a9c12 * HamDist_loop_percentage) ||
                         (Idd909220a9540c998e23f1b06cfca187d9d83bc0673aeafbd0ed6c20c9d39f4d > HamDist_loop_max)
                         ) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b0;
                       end else if (HamDist_sum_mm == 0) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b1;
                       end

               end  //Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e
               else begin // else I28391d3bc64ec15cbb090426b04aa6b7649c3cc85f11230bb0105e02d15e3624 Id34aef7affeaf78c7f4c29e3691a98e841168f86987161bc0d3906da392be76e
                    //wait for Ib9776d7ddf459c9ad5b0e1d6ac61e27befb5e99fd62446677600d7cacef544d0 start_dec to I913a4cb91be20332f3559f8070255d7ac3e6228bb423f4441551d3f783e7d4f4 I2ad8a7049d7c5511ac254f5f51fe70a046ebd884729056f0fe57f5160d467153 Ib4dc66dde806261bdda8607d8707aa727d308cd80272381a5583f63899918467
                    //converged_loops_ended <= 1'b0;
                    //converged_pass_fail <= 1'b0;
               end


          end  //start_dec
       end  //rstn
   end

//tmp_bit valid Ib8d31e852725afb1e26d53bab6095b2bff1749c9275be13ed1c05a56ed31ec09 I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0
// I9390298f3fb0c5b160498935d79cb139aef28e1c47358b4bbba61862b9c26e59 Ic501935a6b2b247d007e9860becbe4c13d6561af9fc8b73ba24c8b2a7a80cb22 I6e16db102267e6e7de7f08f9c28836861561b6ac5a9aec0d26e263c37267f54e I582967534d0f909d196b97f9e6921342777aea87b46fa52df165389db1fb8ccf I9ff94c3eb0c1d350b76101c553e6e70c1178b96fc7fd738182e39e2a3f1b9ebe or Ia70f53bb8550815bbefa894416109ff60708dbd3c7f57d1218df1f55d50fe467 Ib7bdf7a2d6e73e58d69a667ad9b63f706dd96bbbc4a8187914fc34646a1e003b
always_comb HamDist_cntr_inc_converged_valid = I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0;

//I1785cfc3bc6ac7738e8b38cdccd1af12563c2b9070e07af336a1bf8c0f772b6a Ia4c3ed04a95a3da14a9d235c83d868bed7c0f45cf7f3faa751ee8f50598d2211 Ib8d31e852725afb1e26d53bab6095b2bff1749c9275be13ed1c05a56ed31ec09 valid ??

always_comb I6d0b0c1a3968ec36626f19660bedfe0a538a7835edd2a21dd3f4ce0fe2c5c86b = I4b0c82ecfe5c4df9ab1b659484cba58f7d32110d375edf6450aa01ea77dde4c0;
always_comb hamming_code_calc_out             = I6d0b0c1a3968ec36626f19660bedfe0a538a7835edd2a21dd3f4ce0fe2c5c86b;


`ifdef ENCRYPT
`endif

endmodule

//C If029c1f097c0b6dc260a6c5304ad63ce886f7b6078deb247e269b295dd8c9555: I5f75057e98eefa9da67b1a59d3d184f5c0315a905ebe0f6ddfe89aef6413c683 I148de9c5a7a44d19e56cd9ae1a554bf67847afb0c58f6e12fa29ac7ddfca9940:0.100000 I3955f8fd92cda2c17a22e4cccf13c595bc7975089af39fd576cb1be59c0b8269:2.197225 percent_probability_int:'d4500

 //I6ede6cac45f64ed08afc0391ecf38a70942e66382fdad32454a8e52bbe5673d2 I59e61154e1a87dffab5b71a93bf419a969a0a85ae8e300adf0c479acfdc2a59c valid I5694d08a2e53ffcae0c3103e5ad6f6076abd960eb1f8a56577040bc1028f702b I98c1eb4ee93476743763878fcb96a25fbc9a175074d64004779ecb5242f645e6
//y_int:
 //44010bdd34c9a17a9dc5c9798ef00a0604fe89b67904e634be0b
//If3db4f2de25b43f2d2b33fab02836601f68e9641146eacef45de90905b65ab10:
 //0200400200100008100880c0000680200320002200
//C If029c1f097c0b6dc260a6c5304ad63ce886f7b6078deb247e269b295dd8c9555: I5f75057e98eefa9da67b1a59d3d184f5c0315a905ebe0f6ddfe89aef6413c683 I148de9c5a7a44d19e56cd9ae1a554bf67847afb0c58f6e12fa29ac7ddfca9940:0.038462 I3955f8fd92cda2c17a22e4cccf13c595bc7975089af39fd576cb1be59c0b8269:3.218876 percent_probability_int:'d6592
