//`include "GF2_LDPC_flogtanh_0x0000f_assign_inc.sv"
//always_comb begin
              I00c7f323bbe2c226738efd26b205128d['h00000] = 
          (!flogtanh_sel['h0000f]) ? 
                       Iaf491f5f8d1574e1cb610cbd3edeca68['h00000] : //%
                       Iaf491f5f8d1574e1cb610cbd3edeca68['h00001] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00001] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h00002] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00002] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h00004] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00003] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h00006] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00004] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h00008] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00005] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h0000a] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00006] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h0000c] ;
//end
//always_comb begin // 
               I00c7f323bbe2c226738efd26b205128d['h00007] =  Iaf491f5f8d1574e1cb610cbd3edeca68['h0000e] ;
//end
