//`include "GF2_LDPC_flogtanh_0x00004_assign_inc.sv"
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00000] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00000] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00001] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00001] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00002] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00003] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00002] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00004] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00005] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00003] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00006] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00007] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00004] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00008] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00009] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00005] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0000a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0000b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00006] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0000c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0000d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00007] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0000e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0000f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00008] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00010] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00011] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00009] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00012] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00013] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00014] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00015] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00016] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00017] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00018] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00019] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0001a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0001b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0001c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0001d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0001e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0001f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00010] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00020] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00021] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00011] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00022] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00023] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00012] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00024] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00025] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00013] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00026] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00027] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00014] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00028] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00029] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00015] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0002a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0002b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00016] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0002c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0002d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00017] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0002e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0002f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00018] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00030] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00031] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00019] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00032] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00033] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00034] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00035] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00036] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00037] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00038] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00039] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0003a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0003b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0003c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0003d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0003e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0003f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00020] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00040] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00041] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00021] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00042] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00043] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00022] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00044] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00045] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00023] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00046] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00047] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00024] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00048] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00049] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00025] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0004a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0004b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00026] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0004c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0004d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00027] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0004e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0004f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00028] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00050] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00051] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00029] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00052] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00053] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00054] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00055] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00056] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00057] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00058] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00059] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0005a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0005b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0005c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0005d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0005e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0005f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00030] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00060] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00061] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00031] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00062] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00063] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00032] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00064] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00065] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00033] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00066] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00067] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00034] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00068] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00069] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00035] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0006a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0006b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00036] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0006c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0006d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00037] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0006e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0006f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00038] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00070] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00071] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00039] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00072] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00073] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00074] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00075] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00076] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00077] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00078] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00079] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0007a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0007b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0007c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0007d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0007e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0007f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00040] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00080] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00081] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00041] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00082] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00083] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00042] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00084] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00085] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00043] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00086] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00087] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00044] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00088] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00089] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00045] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0008a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0008b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00046] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0008c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0008d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00047] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0008e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0008f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00048] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00090] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00091] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00049] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00092] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00093] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00094] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00095] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00096] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00097] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00098] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00099] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0009a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0009b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0009c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0009d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0009e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0009f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00050] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00051] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00052] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00053] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00054] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000a9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00055] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000aa] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ab] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00056] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ac] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ad] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00057] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ae] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000af] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00058] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00059] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000b9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ba] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000bb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000bc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000bd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000be] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000bf] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00060] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00061] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00062] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00063] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00064] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000c9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00065] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ca] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000cb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00066] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000cc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000cd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00067] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ce] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000cf] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00068] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00069] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000d9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000da] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000db] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000dc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000dd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000de] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000df] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00070] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00071] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00072] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00073] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00074] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000e9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00075] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ea] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000eb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00076] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ec] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ed] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00077] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ee] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ef] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00078] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00079] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000f9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000fa] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000fb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000fc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000fd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000fe] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h000ff] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00080] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00100] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00101] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00081] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00102] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00103] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00082] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00104] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00105] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00083] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00106] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00107] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00084] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00108] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00109] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00085] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0010a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0010b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00086] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0010c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0010d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00087] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0010e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0010f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00088] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00110] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00111] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00089] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00112] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00113] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00114] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00115] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00116] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00117] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00118] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00119] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0011a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0011b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0011c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0011d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0011e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0011f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00090] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00120] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00121] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00091] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00122] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00123] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00092] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00124] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00125] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00093] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00126] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00127] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00094] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00128] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00129] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00095] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0012a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0012b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00096] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0012c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0012d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00097] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0012e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0012f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00098] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00130] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00131] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00099] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00132] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00133] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00134] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00135] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00136] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00137] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00138] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00139] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0013a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0013b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0013c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0013d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0013e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0013f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a0] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00140] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00141] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a1] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00142] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00143] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a2] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00144] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00145] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a3] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00146] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00147] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00148] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00149] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a5] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0014a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0014b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a6] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0014c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0014d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0014e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0014f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a8] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00150] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00151] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00152] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00153] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000aa] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00154] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00155] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ab] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00156] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00157] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ac] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00158] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00159] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ad] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0015a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0015b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ae] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0015c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0015d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000af] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0015e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0015f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b0] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00160] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00161] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b1] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00162] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00163] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b2] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00164] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00165] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b3] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00166] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00167] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00168] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00169] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b5] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0016a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0016b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b6] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0016c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0016d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0016e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0016f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b8] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00170] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00171] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00172] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00173] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ba] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00174] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00175] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bb] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00176] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00177] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bc] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00178] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00179] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bd] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0017a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0017b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000be] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0017c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0017d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bf] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0017e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0017f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c0] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00180] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00181] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c1] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00182] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00183] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c2] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00184] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00185] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c3] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00186] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00187] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00188] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00189] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c5] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0018a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0018b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c6] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0018c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0018d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0018e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0018f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c8] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00190] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00191] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00192] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00193] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ca] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00194] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00195] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cb] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00196] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00197] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cc] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00198] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00199] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cd] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0019a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0019b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ce] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0019c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0019d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cf] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0019e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0019f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d0] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d1] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d2] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d3] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001a9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d5] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001aa] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ab] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d6] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ac] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ad] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ae] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001af] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d8] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000da] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000db] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000dc] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001b9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000dd] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ba] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001bb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000de] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001bc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001bd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000df] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001be] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001bf] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e0] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e1] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e2] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e3] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001c9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e5] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ca] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001cb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e6] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001cc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001cd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ce] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001cf] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e8] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ea] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000eb] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ec] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001d9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ed] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001da] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001db] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ee] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001dc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001dd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ef] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001de] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001df] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f0] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f1] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f2] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f3] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001e9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f5] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ea] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001eb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f6] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ec] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ed] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ee] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ef] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f8] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f1] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f3] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fa] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f5] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fb] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f7] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fc] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001f9] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fd] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001fa] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001fb] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fe] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001fc] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001fd] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ff] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001fe] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h001ff] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00100] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00200] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00201] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00101] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00202] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00203] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00102] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00204] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00205] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00103] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00206] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00207] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00104] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00208] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00209] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00105] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0020a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0020b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00106] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0020c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0020d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00107] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0020e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0020f] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00108] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00210] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00211] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00109] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00212] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00213] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00214] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00215] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00216] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00217] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00218] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00219] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0021a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0021b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0021c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0021d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0021e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0021f] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00110] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00220] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00111] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00222] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00223] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00112] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00224] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00225] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00113] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00226] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00227] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00114] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00228] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00229] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00115] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0022a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0022b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00116] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0022c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0022d] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00117] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0022e] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00118] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00230] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00231] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00119] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00232] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00233] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00234] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00235] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00236] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00237] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00238] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0023a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0023b] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0023c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0023d] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0023e] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00120] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00240] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00241] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00121] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00242] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00243] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00122] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00244] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00245] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00123] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00246] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00124] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00248] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00249] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00125] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0024a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0024b] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00126] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0024c] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00127] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0024e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0024f] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00128] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00250] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00129] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00252] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00253] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00254] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00255] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00256] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00258] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00259] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0025a] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012e] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0025c] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0025d] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012f] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0025e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0025f] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00130] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00260] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00131] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00262] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00263] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00132] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00264] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00133] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00266] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00267] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00134] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00268] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00135] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0026a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0026b] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00136] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0026c] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00137] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0026e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0026f] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00138] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00270] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00139] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00272] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00273] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00274] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00276] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00277] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00278] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0027a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0027b] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0027c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0027e] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00140] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00280] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00281] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00141] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00282] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00142] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00284] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00285] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00143] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00144] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00288] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00145] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0028a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0028b] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00146] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0028c] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00147] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0028e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0028f] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00148] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00149] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00292] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014a] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00294] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00295] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00298] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0029a] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0029b] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0029c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0029e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00150] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00151] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00152] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002a4] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00153] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002a6] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002a7] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00154] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00155] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002aa] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00156] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ac] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ad] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00157] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00158] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002b0] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00159] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002b2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002b3] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002b8] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ba] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002bb] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002be] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00160] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c1] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00161] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00162] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00163] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c6] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00164] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c8] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002c9] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00165] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00166] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00167] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00168] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002d0] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00169] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002d2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002d3] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002d8] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002da] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002db] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00170] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00171] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002e2] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00172] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002e4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002e5] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00173] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00174] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00175] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00176] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00177] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002ee] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00178] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002f0] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002f1] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00179] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002f8] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017d] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002fa] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002fb] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h002fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00180] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00181] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00182] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00183] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00306] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00184] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00308] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00309] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00185] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0030a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00186] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0030c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00187] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0030e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00188] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00189] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00314] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018b] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00316] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00317] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0031a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0031c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0031e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00190] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00191] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00192] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00324] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00193] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00326] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00327] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00194] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00195] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0032a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00196] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0032c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00197] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0032e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00198] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00199] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00336] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019c] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00338] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00339] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0033a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0033c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0033e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0034a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0034c] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a7] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0034e] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0034f] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0035a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0035c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0035e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00366] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00368] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00369] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0036a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0036c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0036e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0037a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0037c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0037e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00386] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c4] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00388] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00389] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0038a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0038c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0038e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0039a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0039c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0039e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003b0] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d9] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003b2] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003b3] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003f2] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fa] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003f4] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003f5] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h003fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00200] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00201] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00202] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00203] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00204] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00205] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0040a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00206] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0040c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00207] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0040e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00208] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00209] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0041a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0041c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0041e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00210] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00211] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00212] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00213] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00214] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00215] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0042a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00216] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0042c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00217] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0042e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00218] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00219] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0043a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0043c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0043e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00220] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00221] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00222] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00223] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00224] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00225] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0044a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00226] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0044c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00227] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0044e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00228] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00229] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0045a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0045c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0045e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00230] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00231] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00232] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00233] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00234] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00235] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0046a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00236] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0046c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00237] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0046e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00238] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00239] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0047a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0047c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0047e] ;
//end
//always_comb begin
              Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00240] = 
          (!flogtanh_sel['h00004]) ? 
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00480] : //%
                       I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00481] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00241] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00242] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00243] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00244] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00245] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0048a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00246] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0048c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00247] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0048e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00248] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00249] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0049a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0049c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0049e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00250] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00251] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00252] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00253] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00254] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00255] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00256] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00257] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00258] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00259] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00260] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00261] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00262] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00263] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00264] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00265] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00266] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00267] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00268] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00269] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00270] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00271] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00272] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00273] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00274] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00275] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00276] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00277] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00278] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00279] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h004fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00280] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00281] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00282] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00283] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00284] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00285] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0050a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00286] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0050c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00287] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0050e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00288] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00289] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0051a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0051c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0051e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00290] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00291] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00292] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00293] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00294] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00295] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0052a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00296] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0052c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00297] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0052e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00298] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00299] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0053a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0053c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0053e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0054a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0054c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0054e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0055a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0055c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0055e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0056a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0056c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0056e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0057a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0057c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0057e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0058a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0058c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0058e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0059a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0059c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0059e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h005fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00300] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00301] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00302] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00303] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00304] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00305] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0060a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00306] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0060c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00307] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0060e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00308] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00309] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0061a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0061c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0061e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00310] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00311] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00312] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00313] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00314] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00315] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0062a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00316] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0062c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00317] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0062e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00318] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00319] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0063a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0063c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0063e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00320] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00321] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00322] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00323] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00324] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00325] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0064a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00326] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0064c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00327] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0064e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00328] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00329] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0065a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0065c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0065e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00330] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00331] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00332] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00333] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00334] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00335] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0066a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00336] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0066c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00337] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0066e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00338] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00339] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0067a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0067c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0067e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00340] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00341] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00342] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00343] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00344] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00345] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0068a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00346] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0068c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00347] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0068e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00348] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00349] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0069a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0069c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0069e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00350] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00351] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00352] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00353] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00354] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00355] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00356] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00357] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00358] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00359] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00360] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00361] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00362] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00363] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00364] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00365] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00366] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00367] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00368] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00369] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00370] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00371] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00372] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00373] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00374] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00375] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00376] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00377] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00378] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00379] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h006fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00380] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00381] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00382] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00383] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00384] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00385] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0070a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00386] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0070c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00387] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0070e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00388] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00389] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0071a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0071c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0071e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00390] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00391] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00392] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00393] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00394] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00395] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0072a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00396] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0072c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00397] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0072e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00398] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00399] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0073a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0073c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0073e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0074a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0074c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0074e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0075a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0075c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0075e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0076a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0076c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0076e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0077a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0077c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0077e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0078a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0078c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0078e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0079a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0079c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0079e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h007fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00400] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00401] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00402] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00403] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00404] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00405] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0080a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00406] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0080c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00407] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0080e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00408] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00409] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0081a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0081c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0081e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00410] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00411] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00412] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00413] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00414] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00415] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0082a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00416] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0082c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00417] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0082e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00418] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00419] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0083a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0083c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0083e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00420] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00421] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00422] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00423] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00424] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00425] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0084a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00426] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0084c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00427] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0084e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00428] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00429] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0085a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0085c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0085e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00430] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00431] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00432] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00433] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00434] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00435] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0086a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00436] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0086c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00437] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0086e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00438] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00439] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0087a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0087c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0087e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00440] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00441] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00442] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00443] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00444] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00445] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0088a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00446] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0088c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00447] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0088e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00448] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00449] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0089a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0089c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0089e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00450] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00451] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00452] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00453] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00454] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00455] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00456] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00457] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00458] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00459] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00460] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00461] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00462] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00463] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00464] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00465] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00466] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00467] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00468] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00469] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00470] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00471] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00472] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00473] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00474] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00475] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00476] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00477] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00478] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00479] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h008fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00480] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00481] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00482] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00483] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00484] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00485] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0090a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00486] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0090c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00487] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0090e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00488] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00489] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0091a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0091c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0091e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00490] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00491] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00492] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00493] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00494] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00495] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0092a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00496] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0092c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00497] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0092e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00498] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00499] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0093a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0093c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0093e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0094a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0094c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0094e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0095a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0095c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0095e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0096a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0096c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0096e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0097a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0097c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0097e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0098a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0098c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0098e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0099a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0099c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0099e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h009fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00500] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00501] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00502] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00503] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00504] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00505] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00506] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00507] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00508] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00509] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00510] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00511] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00512] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00513] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00514] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00515] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00516] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00517] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00518] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00519] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00520] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00521] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00522] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00523] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00524] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00525] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00526] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00527] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00528] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00529] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00530] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00531] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00532] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00533] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00534] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00535] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00536] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00537] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00538] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00539] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00540] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00541] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00542] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00543] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00544] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00545] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00546] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00547] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00548] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00549] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00550] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00551] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00552] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00553] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00554] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00555] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00556] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00557] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00558] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00559] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00560] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00561] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00562] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00563] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00564] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00565] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00566] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00567] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00568] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00569] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00570] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00571] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00572] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00573] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00574] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00575] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00576] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00577] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00578] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00579] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00580] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00581] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00582] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00583] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00584] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00585] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00586] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00587] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00588] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00589] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00590] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00591] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00592] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00593] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00594] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00595] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00596] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00597] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00598] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00599] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00600] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00601] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00602] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00603] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00604] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00605] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00606] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00607] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00608] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00609] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00610] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00611] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00612] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00613] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00614] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00615] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00616] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00617] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00618] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00619] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00620] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00621] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00622] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00623] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00624] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00625] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00626] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00627] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00628] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00629] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00630] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00631] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00632] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00633] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00634] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00635] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00636] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00637] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00638] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00639] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00640] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00641] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00642] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00643] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00644] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00645] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00646] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00647] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00648] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00649] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00650] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00651] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00652] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00653] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00654] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00655] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00656] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00657] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00658] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00659] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00660] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00661] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00662] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00663] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00664] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00665] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00666] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00667] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00668] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00669] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00670] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00671] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00672] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00673] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00674] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00675] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00676] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00677] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00678] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00679] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00680] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00681] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00682] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00683] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00684] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00685] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00686] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00687] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00688] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00689] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00690] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00691] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00692] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00693] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00694] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00695] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00696] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00697] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00698] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00699] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00700] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00701] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00702] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00703] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00704] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00705] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00706] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00707] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00708] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00709] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00710] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00711] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00712] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00713] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00714] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00715] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00716] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00717] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00718] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00719] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00720] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00721] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00722] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00723] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00724] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00725] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00726] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00727] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00728] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00729] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00730] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00731] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00732] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00733] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00734] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00735] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00736] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00737] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00738] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00739] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00740] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00741] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00742] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00743] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00744] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00745] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00746] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00747] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00748] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00749] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00750] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00751] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00752] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00753] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00754] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00755] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00756] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00757] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00758] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00759] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00760] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00761] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00762] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00763] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00764] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00765] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00766] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00767] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00768] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00769] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00770] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00771] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00772] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00773] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00774] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00775] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00776] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00777] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00778] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00779] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00780] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00781] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00782] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00783] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00784] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00785] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00786] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00787] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00788] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00789] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00790] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00791] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00792] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00793] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00794] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00795] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00796] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00797] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00798] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00799] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h00ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00800] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00801] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00802] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00803] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00804] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00805] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0100a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00806] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0100c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00807] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0100e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00808] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00809] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0101a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0101c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0101e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00810] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00811] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00812] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00813] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00814] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00815] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0102a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00816] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0102c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00817] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0102e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00818] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00819] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0103a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0103c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0103e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00820] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00821] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00822] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00823] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00824] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00825] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0104a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00826] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0104c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00827] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0104e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00828] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00829] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0105a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0105c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0105e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00830] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00831] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00832] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00833] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00834] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00835] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0106a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00836] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0106c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00837] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0106e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00838] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00839] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0107a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0107c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0107e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00840] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00841] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00842] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00843] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00844] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00845] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0108a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00846] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0108c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00847] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0108e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00848] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00849] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0109a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0109c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0109e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00850] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00851] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00852] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00853] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00854] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00855] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00856] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00857] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00858] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00859] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00860] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00861] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00862] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00863] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00864] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00865] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00866] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00867] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00868] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00869] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00870] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00871] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00872] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00873] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00874] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00875] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00876] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00877] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00878] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00879] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h010fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00880] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00881] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00882] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00883] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00884] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00885] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0110a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00886] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0110c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00887] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0110e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00888] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00889] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0111a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0111c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0111e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00890] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00891] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00892] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00893] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00894] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00895] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0112a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00896] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0112c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00897] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0112e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00898] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00899] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0113a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0113c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0113e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0114a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0114c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0114e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0115a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0115c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0115e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0116a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0116c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0116e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0117a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0117c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0117e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0118a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0118c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0118e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0119a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0119c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0119e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h011fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00900] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00901] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00902] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00903] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00904] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00905] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0120a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00906] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0120c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00907] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0120e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00908] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00909] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0121a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0121c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0121e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00910] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00911] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00912] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00913] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00914] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00915] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0122a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00916] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0122c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00917] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0122e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00918] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00919] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0123a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0123c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0123e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00920] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00921] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00922] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00923] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00924] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00925] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0124a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00926] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0124c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00927] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0124e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00928] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00929] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0125a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0125c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0125e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00930] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00931] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00932] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00933] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00934] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00935] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0126a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00936] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0126c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00937] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0126e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00938] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00939] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0127a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0127c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0127e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00940] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00941] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00942] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00943] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00944] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00945] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0128a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00946] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0128c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00947] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0128e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00948] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00949] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0129a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0129c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0129e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00950] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00951] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00952] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00953] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00954] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00955] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00956] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00957] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00958] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00959] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00960] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00961] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00962] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00963] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00964] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00965] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00966] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00967] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00968] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00969] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00970] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00971] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00972] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00973] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00974] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00975] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00976] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00977] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00978] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00979] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h012fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00980] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00981] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00982] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00983] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00984] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00985] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0130a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00986] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0130c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00987] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0130e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00988] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00989] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0131a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0131c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0131e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00990] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00991] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00992] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00993] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00994] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00995] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0132a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00996] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0132c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00997] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0132e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00998] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00999] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0133a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0133c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0133e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0134a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0134c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0134e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0135a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0135c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0135e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0136a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0136c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0136e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0137a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0137c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0137e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0138a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0138c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0138e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0139a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0139c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0139e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h013fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0140a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0140c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0140e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0141a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0141c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0141e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0142a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0142c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0142e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0143a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0143c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0143e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0144a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0144c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0144e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0145a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0145c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0145e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0146a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0146c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0146e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0147a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0147c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0147e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0148a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0148c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0148e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0149a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0149c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0149e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h014fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0150a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0150c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0150e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0151a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0151c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0151e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0152a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0152c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0152e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0153a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0153c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0153e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0154a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0154c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0154e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0155a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0155c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0155e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0156a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0156c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0156e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0157a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0157c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0157e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0158a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0158c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0158e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00acb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00acc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00acd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0159a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ace] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0159c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00acf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0159e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ada] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00adb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00adc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00add] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ade] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00adf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h015fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0160a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0160c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0160e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0161a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0161c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0161e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0162a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0162c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0162e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0163a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0163c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0163e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0164a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0164c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0164e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0165a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0165c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0165e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0166a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0166c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0166e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0167a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0167c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0167e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0168a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0168c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0168e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0169a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0169c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0169e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h016fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0170a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0170c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0170e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0171a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0171c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0171e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0172a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0172c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0172e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0173a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0173c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0173e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0174a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0174c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0174e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00baa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0175a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0175c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00baf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0175e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0176a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0176c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0176e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0177a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0177c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0177e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0178a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0178c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0178e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0179a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0179c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0179e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00beb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h017fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0180a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0180c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0180e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0181a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0181c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0181e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0182a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0182c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0182e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0183a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0183c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0183e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0184a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0184c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0184e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0185a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0185c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0185e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0186a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0186c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0186e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0187a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0187c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0187e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0188a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0188c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0188e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0189a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0189c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0189e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h018fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0190a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0190c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0190e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0191a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0191c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0191e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0192a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0192c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0192e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0193a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0193c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0193e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0194a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0194c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0194e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00caa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0195a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0195c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00caf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0195e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0196a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0196c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0196e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0197a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0197c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0197e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0198a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0198c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0198e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ccb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ccc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ccd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0199a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0199c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ccf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0199e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ceb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ced] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h019fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00daa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00daf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ddb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ddc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ddd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ddf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00deb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ded] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00def] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ead] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ecb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ecc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ecd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ece] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ecf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00edb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00edc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00edd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ede] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00edf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00faa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00faf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00feb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h01ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01000] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01001] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01002] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01003] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01004] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01005] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0200a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01006] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0200c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01007] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0200e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01008] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01009] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0201a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0201c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0201e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01010] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01011] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01012] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01013] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01014] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01015] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0202a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01016] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0202c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01017] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0202e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01018] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01019] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0203a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0203c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0203e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01020] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01021] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01022] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01023] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01024] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01025] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0204a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01026] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0204c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01027] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0204e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01028] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01029] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0205a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0205c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0205e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01030] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01031] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01032] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01033] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01034] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01035] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0206a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01036] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0206c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01037] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0206e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01038] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01039] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0207a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0207c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0207e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01040] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01041] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01042] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01043] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01044] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01045] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0208a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01046] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0208c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01047] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0208e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01048] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01049] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0209a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0209c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0209e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01050] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01051] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01052] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01053] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01054] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01055] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01056] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01057] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01058] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01059] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01060] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01061] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01062] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01063] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01064] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01065] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01066] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01067] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01068] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01069] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01070] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01071] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01072] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01073] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01074] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01075] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01076] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01077] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01078] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01079] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h020fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01080] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01081] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01082] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01083] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01084] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01085] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0210a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01086] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0210c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01087] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0210e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01088] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01089] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0211a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0211c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0211e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01090] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01091] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01092] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01093] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01094] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01095] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0212a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01096] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0212c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01097] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0212e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01098] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01099] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0213a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0213c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0213e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0214a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0214c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0214e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0215a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0215c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0215e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0216a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0216c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0216e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0217a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0217c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0217e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0218a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0218c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0218e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0219a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0219c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0219e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h021fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01100] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01101] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01102] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01103] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01104] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01105] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0220a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01106] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0220c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01107] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0220e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01108] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01109] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0221a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0221c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0221e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01110] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01111] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01112] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01113] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01114] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01115] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0222a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01116] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0222c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01117] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0222e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01118] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01119] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0223a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0223c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0223e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01120] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01121] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01122] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01123] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01124] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01125] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0224a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01126] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0224c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01127] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0224e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01128] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01129] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0225a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0225c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0225e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01130] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01131] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01132] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01133] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01134] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01135] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0226a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01136] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0226c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01137] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0226e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01138] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01139] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0227a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0227c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0227e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01140] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01141] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01142] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01143] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01144] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01145] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0228a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01146] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0228c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01147] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0228e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01148] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01149] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0229a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0229c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0229e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01150] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01151] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01152] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01153] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01154] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01155] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01156] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01157] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01158] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01159] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01160] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01161] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01162] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01163] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01164] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01165] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01166] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01167] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01168] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01169] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01170] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01171] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01172] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01173] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01174] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01175] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01176] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01177] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01178] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01179] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h022fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01180] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01181] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01182] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01183] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01184] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01185] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0230a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01186] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0230c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01187] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0230e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01188] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01189] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0231a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0231c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0231e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01190] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01191] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01192] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01193] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01194] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01195] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0232a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01196] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0232c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01197] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0232e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01198] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01199] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0233a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0233c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0233e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0234a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0234c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0234e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0235a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0235c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0235e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0236a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0236c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0236e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0237a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0237c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0237e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0238a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0238c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0238e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0239a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0239c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0239e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h023fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01200] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01201] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01202] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01203] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01204] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01205] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0240a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01206] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0240c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01207] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0240e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01208] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01209] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0241a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0241c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0241e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01210] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01211] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01212] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01213] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01214] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01215] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0242a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01216] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0242c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01217] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0242e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01218] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01219] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0243a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0243c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0243e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01220] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01221] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01222] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01223] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01224] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01225] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0244a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01226] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0244c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01227] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0244e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01228] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01229] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0245a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0245c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0245e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01230] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01231] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01232] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01233] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01234] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01235] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0246a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01236] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0246c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01237] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0246e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01238] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01239] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0247a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0247c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0247e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01240] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01241] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01242] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01243] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01244] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01245] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0248a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01246] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0248c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01247] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0248e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01248] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01249] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0249a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0249c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0249e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01250] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01251] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01252] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01253] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01254] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01255] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01256] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01257] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01258] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01259] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01260] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01261] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01262] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01263] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01264] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01265] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01266] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01267] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01268] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01269] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01270] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01271] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01272] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01273] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01274] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01275] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01276] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01277] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01278] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01279] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h024fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01280] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01281] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01282] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01283] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01284] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01285] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0250a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01286] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0250c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01287] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0250e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01288] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01289] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0251a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0251c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0251e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01290] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01291] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01292] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01293] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01294] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01295] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0252a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01296] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0252c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01297] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0252e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01298] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01299] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0253a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0253c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0253e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0254a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0254c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0254e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0255a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0255c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0255e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0256a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0256c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0256e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0257a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0257c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0257e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0258a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0258c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0258e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0259a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0259c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0259e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h025fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01300] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01301] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01302] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01303] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01304] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01305] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0260a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01306] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0260c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01307] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0260e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01308] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01309] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0261a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0261c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0261e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01310] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01311] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01312] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01313] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01314] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01315] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0262a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01316] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0262c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01317] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0262e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01318] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01319] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0263a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0263c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0263e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01320] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01321] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01322] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01323] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01324] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01325] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0264a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01326] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0264c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01327] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0264e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01328] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01329] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0265a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0265c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0265e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01330] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01331] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01332] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01333] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01334] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01335] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0266a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01336] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0266c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01337] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0266e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01338] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01339] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0267a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0267c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0267e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01340] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01341] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01342] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01343] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01344] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01345] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0268a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01346] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0268c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01347] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0268e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01348] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01349] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0269a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0269c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0269e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01350] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01351] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01352] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01353] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01354] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01355] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01356] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01357] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01358] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01359] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01360] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01361] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01362] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01363] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01364] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01365] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01366] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01367] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01368] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01369] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01370] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01371] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01372] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01373] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01374] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01375] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01376] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01377] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01378] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01379] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h026fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01380] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01381] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01382] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01383] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01384] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01385] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0270a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01386] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0270c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01387] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0270e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01388] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01389] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0271a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0271c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0271e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01390] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01391] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01392] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01393] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01394] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01395] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0272a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01396] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0272c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01397] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0272e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01398] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01399] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0273a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0273c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0273e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0274a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0274c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0274e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0275a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0275c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0275e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0276a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0276c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0276e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0277a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0277c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0277e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0278a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0278c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0278e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0279a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0279c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0279e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h027fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01400] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01401] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01402] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01403] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01404] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01405] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0280a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01406] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0280c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01407] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0280e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01408] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01409] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0281a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0281c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0281e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01410] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01411] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01412] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01413] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01414] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01415] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0282a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01416] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0282c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01417] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0282e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01418] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01419] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0283a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0283c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0283e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01420] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01421] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01422] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01423] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01424] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01425] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0284a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01426] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0284c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01427] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0284e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01428] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01429] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0285a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0285c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0285e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01430] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01431] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01432] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01433] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01434] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01435] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0286a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01436] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0286c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01437] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0286e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01438] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01439] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0287a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0287c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0287e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01440] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01441] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01442] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01443] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01444] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01445] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0288a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01446] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0288c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01447] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0288e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01448] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01449] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0289a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0289c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0289e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01450] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01451] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01452] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01453] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01454] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01455] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01456] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01457] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01458] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01459] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01460] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01461] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01462] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01463] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01464] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01465] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01466] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01467] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01468] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01469] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01470] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01471] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01472] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01473] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01474] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01475] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01476] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01477] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01478] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01479] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h028fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01480] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01481] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01482] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01483] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01484] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01485] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0290a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01486] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0290c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01487] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0290e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01488] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01489] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0291a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0291c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0291e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01490] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01491] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01492] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01493] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01494] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01495] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0292a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01496] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0292c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01497] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0292e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01498] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01499] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0293a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0293c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0293e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0294a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0294c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0294e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0295a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0295c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0295e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0296a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0296c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0296e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0297a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0297c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0297e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0298a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0298c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0298e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0299a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0299c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0299e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h029fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01500] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01501] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01502] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01503] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01504] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01505] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01506] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01507] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01508] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01509] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01510] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01511] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01512] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01513] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01514] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01515] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01516] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01517] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01518] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01519] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01520] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01521] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01522] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01523] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01524] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01525] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01526] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01527] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01528] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01529] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01530] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01531] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01532] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01533] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01534] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01535] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01536] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01537] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01538] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01539] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01540] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01541] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01542] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01543] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01544] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01545] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01546] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01547] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01548] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01549] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01550] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01551] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01552] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01553] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01554] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01555] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01556] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01557] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01558] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01559] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01560] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01561] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01562] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01563] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01564] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01565] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01566] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01567] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01568] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01569] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01570] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01571] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01572] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01573] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01574] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01575] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01576] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01577] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01578] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01579] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01580] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01581] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01582] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01583] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01584] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01585] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01586] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01587] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01588] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01589] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01590] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01591] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01592] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01593] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01594] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01595] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01596] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01597] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01598] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01599] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01600] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01601] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01602] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01603] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01604] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01605] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01606] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01607] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01608] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01609] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01610] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01611] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01612] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01613] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01614] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01615] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01616] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01617] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01618] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01619] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01620] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01621] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01622] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01623] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01624] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01625] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01626] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01627] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01628] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01629] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01630] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01631] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01632] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01633] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01634] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01635] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01636] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01637] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01638] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01639] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01640] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01641] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01642] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01643] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01644] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01645] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01646] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01647] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01648] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01649] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01650] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01651] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01652] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01653] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01654] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01655] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01656] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01657] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01658] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01659] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01660] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01661] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01662] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01663] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01664] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01665] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01666] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01667] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01668] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01669] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01670] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01671] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01672] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01673] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01674] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01675] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01676] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01677] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01678] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01679] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01680] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01681] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01682] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01683] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01684] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01685] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01686] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01687] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01688] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01689] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01690] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01691] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01692] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01693] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01694] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01695] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01696] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01697] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01698] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01699] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01700] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01701] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01702] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01703] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01704] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01705] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01706] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01707] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01708] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01709] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01710] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01711] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01712] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01713] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01714] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01715] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01716] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01717] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01718] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01719] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01720] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01721] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01722] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01723] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01724] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01725] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01726] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01727] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01728] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01729] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01730] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01731] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01732] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01733] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01734] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01735] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01736] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01737] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01738] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01739] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01740] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01741] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01742] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01743] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01744] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01745] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01746] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01747] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01748] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01749] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01750] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01751] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01752] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01753] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01754] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01755] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01756] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01757] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01758] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01759] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01760] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01761] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01762] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01763] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01764] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01765] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01766] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01767] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01768] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01769] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01770] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01771] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01772] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01773] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01774] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01775] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01776] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01777] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01778] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01779] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01780] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01781] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01782] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01783] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01784] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01785] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01786] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01787] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01788] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01789] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01790] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01791] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01792] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01793] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01794] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01795] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01796] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01797] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01798] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01799] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h02ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01800] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01801] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01802] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01803] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01804] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01805] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0300a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01806] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0300c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01807] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0300e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01808] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01809] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0301a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0301c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0301e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01810] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01811] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01812] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01813] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01814] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01815] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0302a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01816] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0302c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01817] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0302e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01818] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01819] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0303a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0303c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0303e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01820] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01821] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01822] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01823] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01824] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01825] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0304a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01826] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0304c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01827] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0304e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01828] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01829] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0305a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0305c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0305e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01830] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01831] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01832] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01833] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01834] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01835] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0306a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01836] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0306c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01837] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0306e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01838] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01839] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0307a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0307c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0307e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01840] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01841] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01842] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01843] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01844] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01845] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0308a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01846] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0308c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01847] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0308e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01848] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01849] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0309a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0309c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0309e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01850] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01851] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01852] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01853] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01854] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01855] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01856] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01857] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01858] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01859] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01860] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01861] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01862] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01863] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01864] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01865] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01866] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01867] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01868] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01869] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01870] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01871] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01872] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01873] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01874] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01875] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01876] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01877] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01878] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01879] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h030fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01880] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01881] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01882] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01883] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01884] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01885] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0310a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01886] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0310c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01887] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0310e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01888] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01889] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0311a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0311c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0311e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01890] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01891] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01892] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01893] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01894] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01895] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0312a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01896] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0312c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01897] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0312e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01898] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01899] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0313a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0313c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0313e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0314a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0314c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0314e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0315a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0315c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0315e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0316a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0316c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0316e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0317a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0317c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0317e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0318a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0318c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0318e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0319a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0319c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0319e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h031fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01900] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01901] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01902] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01903] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01904] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01905] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0320a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01906] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0320c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01907] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0320e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01908] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01909] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0321a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0321c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0321e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01910] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01911] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01912] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01913] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01914] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01915] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0322a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01916] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0322c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01917] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0322e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01918] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01919] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0323a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0323c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0323e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01920] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01921] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01922] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01923] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01924] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01925] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0324a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01926] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0324c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01927] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0324e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01928] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01929] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0325a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0325c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0325e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01930] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01931] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01932] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01933] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01934] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01935] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0326a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01936] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0326c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01937] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0326e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01938] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01939] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0327a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0327c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0327e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01940] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01941] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01942] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01943] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01944] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01945] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0328a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01946] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0328c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01947] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0328e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01948] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01949] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0329a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0329c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0329e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01950] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01951] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01952] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01953] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01954] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01955] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01956] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01957] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01958] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01959] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01960] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01961] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01962] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01963] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01964] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01965] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01966] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01967] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01968] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01969] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01970] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01971] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01972] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01973] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01974] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01975] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01976] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01977] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01978] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01979] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h032fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01980] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01981] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01982] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01983] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01984] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01985] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0330a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01986] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0330c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01987] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0330e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01988] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01989] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0331a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0331c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0331e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01990] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01991] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01992] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01993] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01994] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01995] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0332a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01996] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0332c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01997] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0332e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01998] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01999] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0333a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0333c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0333e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0334a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0334c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0334e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0335a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0335c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0335e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0336a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0336c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0336e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0337a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0337c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0337e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0338a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0338c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0338e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0339a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0339c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0339e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h033fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0340a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0340c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0340e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0341a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0341c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0341e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0342a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0342c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0342e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0343a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0343c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0343e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0344a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0344c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0344e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0345a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0345c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0345e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0346a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0346c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0346e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0347a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0347c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0347e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0348a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0348c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0348e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0349a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0349c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0349e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h034fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0350a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0350c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0350e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0351a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0351c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0351e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0352a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0352c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0352e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0353a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0353c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0353e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0354a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0354c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0354e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0355a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0355c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0355e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0356a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0356c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0356e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0357a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0357c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0357e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0358a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0358c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0358e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01acb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01acc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01acd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0359a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ace] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0359c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01acf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0359e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ada] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01adb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01adc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01add] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ade] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01adf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h035fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0360a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0360c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0360e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0361a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0361c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0361e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0362a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0362c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0362e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0363a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0363c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0363e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0364a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0364c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0364e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0365a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0365c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0365e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0366a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0366c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0366e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0367a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0367c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0367e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0368a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0368c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0368e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0369a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0369c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0369e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h036fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0370a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0370c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0370e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0371a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0371c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0371e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0372a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0372c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0372e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0373a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0373c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0373e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0374a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0374c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0374e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01baa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0375a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0375c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01baf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0375e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0376a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0376c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0376e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0377a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0377c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0377e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0378a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0378c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0378e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0379a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0379c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0379e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01beb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h037fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0380a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0380c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0380e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0381a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0381c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0381e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0382a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0382c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0382e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0383a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0383c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0383e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0384a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0384c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0384e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0385a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0385c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0385e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0386a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0386c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0386e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0387a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0387c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0387e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0388a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0388c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0388e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0389a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0389c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0389e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h038fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0390a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0390c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0390e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0391a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0391c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0391e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0392a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0392c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0392e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0393a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0393c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0393e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0394a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0394c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0394e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01caa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0395a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0395c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01caf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0395e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0396a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0396c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0396e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0397a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0397c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0397e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0398a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0398c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0398e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ccb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ccc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ccd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0399a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0399c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ccf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0399e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ceb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ced] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h039fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01daa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01daf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ddb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ddc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ddd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ddf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01deb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ded] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01def] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ead] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ecb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ecc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ecd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ece] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ecf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01edb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01edc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01edd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ede] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01edf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01faa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01faf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01feb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h03ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02000] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02001] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02002] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02003] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02004] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02005] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0400a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02006] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0400c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02007] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0400e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02008] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02009] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0401a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0401c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0401e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02010] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02011] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02012] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02013] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02014] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02015] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0402a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02016] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0402c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02017] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0402e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02018] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02019] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0403a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0403c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0403e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02020] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02021] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02022] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02023] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02024] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02025] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0404a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02026] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0404c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02027] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0404e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02028] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02029] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0405a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0405c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0405e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02030] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02031] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02032] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02033] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02034] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02035] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0406a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02036] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0406c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02037] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0406e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02038] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02039] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0407a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0407c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0407e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02040] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02041] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02042] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02043] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02044] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02045] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0408a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02046] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0408c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02047] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0408e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02048] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02049] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0409a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0409c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0409e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02050] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02051] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02052] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02053] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02054] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02055] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02056] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02057] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02058] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02059] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02060] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02061] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02062] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02063] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02064] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02065] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02066] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02067] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02068] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02069] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02070] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02071] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02072] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02073] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02074] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02075] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02076] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02077] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02078] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02079] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h040fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02080] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02081] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02082] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02083] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02084] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02085] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0410a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02086] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0410c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02087] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0410e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02088] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02089] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0411a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0411c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0411e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02090] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02091] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02092] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02093] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02094] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02095] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0412a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02096] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0412c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02097] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0412e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02098] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02099] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0413a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0413c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0413e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0414a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0414c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0414e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0415a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0415c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0415e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0416a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0416c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0416e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0417a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0417c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0417e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0418a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0418c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0418e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0419a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0419c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0419e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h041fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02100] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02101] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02102] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02103] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02104] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02105] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0420a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02106] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0420c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02107] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0420e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02108] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02109] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0421a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0421c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0421e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02110] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02111] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02112] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02113] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02114] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02115] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0422a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02116] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0422c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02117] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0422e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02118] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02119] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0423a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0423c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0423e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02120] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02121] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02122] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02123] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02124] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02125] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0424a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02126] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0424c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02127] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0424e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02128] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02129] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0425a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0425c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0425e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02130] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02131] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02132] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02133] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02134] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02135] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0426a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02136] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0426c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02137] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0426e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02138] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02139] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0427a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0427c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0427e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02140] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02141] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02142] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02143] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02144] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02145] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0428a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02146] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0428c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02147] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0428e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02148] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02149] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0429a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0429c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0429e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02150] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02151] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02152] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02153] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02154] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02155] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02156] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02157] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02158] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02159] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02160] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02161] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02162] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02163] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02164] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02165] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02166] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02167] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02168] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02169] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02170] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02171] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02172] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02173] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02174] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02175] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02176] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02177] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02178] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02179] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h042fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02180] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02181] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02182] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02183] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02184] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02185] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0430a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02186] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0430c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02187] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0430e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02188] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02189] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0431a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0431c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0431e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02190] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02191] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02192] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02193] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02194] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02195] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0432a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02196] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0432c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02197] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0432e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02198] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02199] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0433a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0433c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0433e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0434a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0434c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0434e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0435a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0435c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0435e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0436a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0436c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0436e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0437a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0437c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0437e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0438a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0438c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0438e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0439a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0439c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0439e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h043fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02200] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02201] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02202] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02203] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02204] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02205] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0440a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02206] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0440c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02207] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0440e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02208] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02209] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0441a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0441c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0441e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02210] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02211] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02212] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02213] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02214] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02215] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0442a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02216] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0442c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02217] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0442e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02218] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02219] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0443a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0443c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0443e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02220] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02221] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02222] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02223] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02224] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02225] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0444a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02226] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0444c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02227] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0444e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02228] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02229] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0445a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0445c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0445e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02230] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02231] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02232] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02233] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02234] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02235] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0446a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02236] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0446c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02237] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0446e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02238] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02239] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0447a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0447c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0447e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02240] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02241] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02242] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02243] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02244] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02245] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0448a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02246] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0448c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02247] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0448e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02248] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02249] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0449a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0449c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0449e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02250] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02251] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02252] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02253] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02254] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02255] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02256] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02257] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02258] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02259] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02260] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02261] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02262] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02263] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02264] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02265] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02266] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02267] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02268] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02269] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02270] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02271] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02272] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02273] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02274] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02275] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02276] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02277] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02278] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02279] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h044fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02280] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02281] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02282] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02283] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02284] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02285] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0450a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02286] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0450c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02287] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0450e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02288] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02289] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0451a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0451c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0451e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02290] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02291] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02292] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02293] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02294] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02295] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0452a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02296] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0452c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02297] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0452e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02298] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02299] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0453a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0453c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0453e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0454a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0454c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0454e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0455a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0455c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0455e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0456a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0456c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0456e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0457a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0457c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0457e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0458a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0458c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0458e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0459a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0459c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0459e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h045fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02300] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02301] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02302] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02303] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02304] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02305] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0460a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02306] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0460c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02307] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0460e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02308] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02309] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0461a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0461c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0461e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02310] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02311] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02312] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02313] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02314] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02315] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0462a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02316] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0462c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02317] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0462e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02318] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02319] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0463a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0463c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0463e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02320] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02321] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02322] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02323] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02324] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02325] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0464a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02326] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0464c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02327] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0464e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02328] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02329] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0465a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0465c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0465e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02330] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02331] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02332] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02333] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02334] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02335] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0466a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02336] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0466c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02337] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0466e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02338] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02339] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0467a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0467c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0467e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02340] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02341] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02342] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02343] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02344] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02345] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0468a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02346] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0468c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02347] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0468e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02348] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02349] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0469a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0469c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0469e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02350] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02351] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02352] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02353] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02354] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02355] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02356] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02357] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02358] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02359] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02360] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02361] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02362] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02363] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02364] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02365] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02366] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02367] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02368] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02369] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02370] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02371] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02372] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02373] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02374] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02375] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02376] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02377] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02378] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02379] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h046fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02380] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02381] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02382] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02383] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02384] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02385] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0470a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02386] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0470c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02387] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0470e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02388] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02389] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0471a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0471c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0471e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02390] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02391] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02392] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02393] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02394] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02395] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0472a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02396] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0472c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02397] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0472e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02398] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02399] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0473a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0473c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0473e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0474a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0474c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0474e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0475a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0475c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0475e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0476a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0476c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0476e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0477a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0477c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0477e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0478a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0478c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0478e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0479a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0479c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0479e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h047fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02400] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02401] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02402] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02403] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02404] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02405] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0480a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02406] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0480c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02407] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0480e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02408] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02409] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0481a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0481c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0481e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02410] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02411] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02412] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02413] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02414] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02415] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0482a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02416] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0482c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02417] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0482e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02418] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02419] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0483a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0483c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0483e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02420] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02421] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02422] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02423] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02424] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02425] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0484a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02426] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0484c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02427] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0484e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02428] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02429] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0485a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0485c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0485e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02430] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02431] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02432] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02433] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02434] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02435] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0486a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02436] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0486c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02437] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0486e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02438] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02439] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0487a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0487c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0487e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02440] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02441] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02442] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02443] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02444] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02445] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0488a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02446] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0488c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02447] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0488e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02448] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02449] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0489a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0489c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0489e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02450] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02451] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02452] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02453] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02454] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02455] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02456] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02457] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02458] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02459] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02460] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02461] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02462] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02463] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02464] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02465] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02466] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02467] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02468] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02469] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02470] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02471] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02472] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02473] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02474] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02475] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02476] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02477] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02478] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02479] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h048fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02480] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02481] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02482] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02483] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02484] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02485] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0490a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02486] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0490c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02487] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0490e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02488] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02489] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0491a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0491c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0491e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02490] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02491] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02492] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02493] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02494] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02495] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0492a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02496] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0492c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02497] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0492e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02498] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02499] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0493a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0493c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0493e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0494a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0494c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0494e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0495a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0495c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0495e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0496a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0496c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0496e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0497a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0497c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0497e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0498a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0498c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0498e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0499a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0499c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0499e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h049fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02500] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02501] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02502] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02503] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02504] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02505] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02506] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02507] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02508] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02509] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02510] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02511] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02512] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02513] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02514] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02515] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02516] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02517] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02518] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02519] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02520] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02521] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02522] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02523] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02524] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02525] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02526] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02527] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02528] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02529] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02530] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02531] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02532] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02533] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02534] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02535] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02536] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02537] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02538] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02539] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02540] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02541] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02542] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02543] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02544] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02545] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02546] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02547] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02548] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02549] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02550] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02551] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02552] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02553] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02554] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02555] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02556] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02557] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02558] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02559] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02560] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02561] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02562] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02563] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02564] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02565] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02566] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02567] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02568] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02569] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02570] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02571] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02572] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02573] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02574] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02575] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02576] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02577] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02578] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02579] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02580] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02581] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02582] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02583] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02584] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02585] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02586] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02587] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02588] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02589] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02590] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02591] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02592] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02593] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02594] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02595] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02596] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02597] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02598] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02599] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02600] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02601] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02602] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02603] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02604] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02605] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02606] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02607] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02608] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02609] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02610] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02611] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02612] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02613] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02614] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02615] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02616] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02617] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02618] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02619] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02620] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02621] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02622] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02623] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02624] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02625] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02626] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02627] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02628] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02629] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02630] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02631] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02632] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02633] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02634] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02635] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02636] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02637] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02638] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02639] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02640] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02641] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02642] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02643] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02644] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02645] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02646] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02647] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02648] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02649] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02650] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02651] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02652] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02653] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02654] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02655] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02656] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02657] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02658] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02659] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02660] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02661] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02662] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02663] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02664] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02665] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02666] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02667] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02668] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02669] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02670] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02671] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02672] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02673] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02674] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02675] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02676] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02677] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02678] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02679] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02680] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02681] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02682] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02683] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02684] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02685] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02686] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02687] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02688] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02689] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02690] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02691] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02692] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02693] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02694] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02695] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02696] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02697] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02698] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02699] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02700] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02701] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02702] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02703] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02704] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02705] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02706] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02707] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02708] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02709] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02710] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02711] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02712] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02713] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02714] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02715] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02716] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02717] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02718] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02719] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02720] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02721] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02722] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02723] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02724] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02725] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02726] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02727] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02728] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02729] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02730] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02731] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02732] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02733] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02734] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02735] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02736] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02737] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02738] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02739] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02740] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02741] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02742] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02743] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02744] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02745] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02746] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02747] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02748] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02749] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02750] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02751] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02752] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02753] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02754] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02755] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02756] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02757] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02758] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02759] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02760] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02761] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02762] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02763] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02764] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02765] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02766] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02767] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02768] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02769] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02770] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02771] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02772] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02773] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02774] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02775] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02776] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02777] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02778] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02779] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02780] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02781] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02782] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02783] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02784] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02785] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02786] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02787] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02788] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02789] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02790] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02791] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02792] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02793] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02794] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02795] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02796] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02797] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02798] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02799] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h04ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02800] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02801] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02802] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02803] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02804] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02805] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0500a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02806] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0500c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02807] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0500e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02808] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02809] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0501a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0501c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0501e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02810] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02811] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02812] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02813] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02814] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02815] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0502a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02816] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0502c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02817] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0502e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02818] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02819] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0503a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0503c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0503e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02820] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02821] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02822] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02823] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02824] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02825] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0504a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02826] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0504c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02827] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0504e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02828] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02829] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0505a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0505c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0505e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02830] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02831] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02832] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02833] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02834] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02835] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0506a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02836] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0506c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02837] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0506e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02838] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02839] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0507a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0507c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0507e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02840] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02841] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02842] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02843] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02844] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02845] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0508a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02846] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0508c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02847] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0508e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02848] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02849] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0509a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0509c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0509e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02850] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02851] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02852] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02853] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02854] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02855] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02856] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02857] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02858] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02859] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02860] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02861] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02862] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02863] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02864] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02865] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02866] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02867] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02868] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02869] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02870] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02871] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02872] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02873] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02874] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02875] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02876] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02877] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02878] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02879] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h050fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02880] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02881] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02882] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02883] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02884] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02885] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0510a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02886] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0510c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02887] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0510e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02888] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02889] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0511a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0511c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0511e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02890] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02891] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02892] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02893] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02894] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02895] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0512a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02896] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0512c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02897] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0512e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02898] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02899] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0513a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0513c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0513e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0514a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0514c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0514e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0515a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0515c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0515e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0516a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0516c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0516e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0517a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0517c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0517e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0518a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0518c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0518e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0519a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0519c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0519e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h051fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02900] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02901] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02902] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02903] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02904] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02905] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0520a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02906] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0520c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02907] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0520e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02908] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02909] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0521a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0521c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0521e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02910] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02911] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02912] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02913] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02914] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02915] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0522a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02916] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0522c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02917] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0522e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02918] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02919] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0523a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0523c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0523e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02920] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02921] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02922] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02923] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02924] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02925] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0524a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02926] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0524c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02927] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0524e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02928] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02929] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0525a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0525c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0525e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02930] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02931] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02932] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02933] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02934] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02935] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0526a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02936] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0526c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02937] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0526e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02938] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02939] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0527a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0527c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0527e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02940] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02941] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02942] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02943] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02944] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02945] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0528a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02946] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0528c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02947] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0528e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02948] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02949] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0529a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0529c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0529e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02950] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02951] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02952] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02953] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02954] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02955] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02956] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02957] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02958] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02959] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02960] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02961] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02962] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02963] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02964] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02965] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02966] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02967] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02968] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02969] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02970] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02971] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02972] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02973] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02974] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02975] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02976] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02977] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02978] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02979] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h052fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02980] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02981] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02982] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02983] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02984] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02985] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0530a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02986] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0530c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02987] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0530e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02988] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02989] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0531a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0531c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0531e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02990] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02991] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02992] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02993] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02994] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02995] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0532a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02996] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0532c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02997] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0532e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02998] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02999] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0533a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0533c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0533e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0534a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0534c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0534e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0535a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0535c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0535e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0536a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0536c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0536e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0537a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0537c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0537e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0538a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0538c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0538e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0539a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0539c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0539e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h053fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0540a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0540c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0540e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0541a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0541c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0541e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0542a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0542c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0542e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0543a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0543c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0543e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0544a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0544c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0544e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0545a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0545c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0545e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0546a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0546c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0546e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0547a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0547c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0547e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0548a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0548c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0548e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0549a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0549c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0549e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h054fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0550a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0550c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0550e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0551a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0551c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0551e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0552a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0552c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0552e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0553a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0553c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0553e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0554a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0554c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0554e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0555a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0555c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0555e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0556a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0556c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0556e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0557a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0557c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0557e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0558a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0558c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0558e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02acb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02acc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02acd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0559a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ace] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0559c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02acf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0559e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ada] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02adb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02adc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02add] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ade] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02adf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h055fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0560a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0560c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0560e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0561a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0561c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0561e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0562a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0562c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0562e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0563a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0563c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0563e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0564a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0564c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0564e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0565a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0565c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0565e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0566a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0566c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0566e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0567a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0567c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0567e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0568a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0568c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0568e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0569a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0569c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0569e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h056fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0570a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0570c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0570e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0571a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0571c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0571e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0572a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0572c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0572e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0573a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0573c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0573e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0574a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0574c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0574e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02baa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0575a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0575c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02baf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0575e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0576a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0576c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0576e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0577a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0577c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0577e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0578a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0578c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0578e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0579a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0579c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0579e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02beb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h057fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0580a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0580c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0580e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0581a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0581c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0581e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0582a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0582c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0582e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0583a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0583c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0583e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0584a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0584c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0584e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0585a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0585c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0585e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0586a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0586c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0586e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0587a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0587c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0587e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0588a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0588c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0588e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0589a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0589c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0589e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h058fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0590a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0590c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0590e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0591a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0591c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0591e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0592a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0592c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0592e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0593a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0593c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0593e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0594a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0594c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0594e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02caa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0595a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0595c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02caf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0595e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0596a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0596c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0596e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0597a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0597c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0597e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0598a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0598c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0598e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ccb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ccc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ccd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0599a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0599c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ccf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0599e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ceb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ced] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h059fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02daa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02daf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ddb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ddc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ddd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ddf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02deb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ded] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02def] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ead] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ecb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ecc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ecd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ece] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ecf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02edb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02edc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02edd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ede] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02edf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02faa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02faf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02feb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h05ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03000] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03001] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03002] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03003] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03004] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03005] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0600a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03006] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0600c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03007] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0600e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03008] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03009] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0601a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0601c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0601e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03010] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03011] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03012] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03013] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03014] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03015] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0602a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03016] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0602c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03017] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0602e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03018] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03019] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0603a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0603c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0603e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03020] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03021] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03022] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03023] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03024] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03025] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0604a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03026] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0604c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03027] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0604e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03028] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03029] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0605a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0605c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0605e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03030] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03031] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03032] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03033] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03034] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03035] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0606a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03036] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0606c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03037] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0606e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03038] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03039] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0607a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0607c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0607e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03040] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03041] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03042] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03043] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03044] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03045] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0608a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03046] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0608c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03047] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0608e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03048] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03049] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0609a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0609c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0609e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03050] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03051] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03052] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03053] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03054] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03055] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03056] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03057] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03058] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03059] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03060] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03061] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03062] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03063] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03064] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03065] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03066] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03067] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03068] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03069] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03070] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03071] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03072] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03073] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03074] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03075] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03076] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03077] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03078] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03079] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h060fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03080] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03081] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03082] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03083] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03084] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03085] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0610a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03086] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0610c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03087] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0610e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03088] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03089] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0611a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0611c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0611e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03090] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03091] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03092] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03093] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03094] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03095] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0612a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03096] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0612c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03097] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0612e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03098] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03099] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0613a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0613c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0613e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0614a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0614c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0614e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0615a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0615c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0615e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0616a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0616c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0616e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0617a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0617c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0617e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0618a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0618c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0618e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0619a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0619c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0619e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h061fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03100] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03101] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03102] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03103] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03104] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03105] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0620a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03106] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0620c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03107] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0620e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03108] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03109] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0621a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0621c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0621e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03110] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03111] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03112] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03113] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03114] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03115] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0622a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03116] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0622c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03117] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0622e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03118] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03119] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0623a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0623c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0623e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03120] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03121] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03122] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03123] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03124] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03125] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0624a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03126] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0624c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03127] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0624e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03128] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03129] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0625a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0625c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0625e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03130] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03131] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03132] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03133] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03134] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03135] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0626a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03136] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0626c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03137] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0626e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03138] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03139] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0627a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0627c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0627e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03140] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03141] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03142] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03143] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03144] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03145] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0628a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03146] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0628c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03147] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0628e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03148] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03149] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0629a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0629c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0629e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03150] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03151] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03152] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03153] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03154] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03155] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03156] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03157] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03158] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03159] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03160] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03161] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03162] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03163] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03164] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03165] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03166] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03167] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03168] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03169] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03170] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03171] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03172] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03173] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03174] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03175] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03176] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03177] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03178] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03179] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h062fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03180] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03181] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03182] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03183] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03184] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03185] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0630a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03186] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0630c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03187] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0630e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03188] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03189] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0631a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0631c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0631e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03190] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03191] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03192] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03193] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03194] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03195] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0632a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03196] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0632c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03197] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0632e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03198] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03199] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0633a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0633c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0633e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0634a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0634c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0634e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0635a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0635c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0635e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0636a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0636c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0636e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0637a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0637c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0637e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0638a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0638c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0638e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0639a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0639c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0639e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h063fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03200] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03201] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03202] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03203] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03204] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03205] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0640a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03206] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0640c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03207] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0640e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03208] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03209] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0641a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0641c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0641e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03210] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03211] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03212] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03213] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03214] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03215] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0642a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03216] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0642c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03217] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0642e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03218] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03219] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0643a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0643c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0643e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03220] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03221] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03222] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03223] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03224] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03225] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0644a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03226] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0644c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03227] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0644e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03228] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03229] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0645a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0645c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0645e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03230] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03231] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03232] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03233] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03234] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03235] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0646a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03236] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0646c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03237] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0646e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03238] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03239] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0647a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0647c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0647e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03240] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03241] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03242] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03243] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03244] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03245] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0648a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03246] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0648c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03247] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0648e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03248] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03249] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0649a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0649c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0649e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03250] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03251] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03252] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03253] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03254] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03255] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03256] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03257] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03258] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03259] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03260] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03261] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03262] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03263] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03264] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03265] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03266] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03267] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03268] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03269] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03270] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03271] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03272] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03273] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03274] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03275] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03276] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03277] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03278] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03279] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h064fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03280] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03281] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03282] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03283] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03284] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03285] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0650a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03286] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0650c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03287] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0650e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03288] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03289] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0651a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0651c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0651e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03290] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03291] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03292] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03293] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03294] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03295] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0652a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03296] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0652c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03297] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0652e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03298] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03299] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0653a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0653c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0653e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0654a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0654c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0654e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0655a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0655c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0655e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0656a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0656c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0656e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0657a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0657c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0657e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0658a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0658c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0658e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0659a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0659c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0659e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h065fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03300] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03301] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03302] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03303] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03304] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03305] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0660a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03306] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0660c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03307] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0660e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03308] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03309] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0661a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0661c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0661e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03310] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03311] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03312] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03313] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03314] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03315] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0662a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03316] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0662c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03317] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0662e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03318] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03319] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0663a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0663c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0663e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03320] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03321] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03322] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03323] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03324] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03325] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0664a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03326] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0664c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03327] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0664e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03328] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03329] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0665a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0665c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0665e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03330] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03331] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03332] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03333] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03334] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03335] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0666a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03336] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0666c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03337] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0666e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03338] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03339] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0667a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0667c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0667e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03340] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03341] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03342] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03343] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03344] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03345] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0668a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03346] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0668c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03347] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0668e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03348] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03349] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0669a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0669c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0669e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03350] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03351] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03352] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03353] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03354] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03355] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03356] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03357] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03358] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03359] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03360] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03361] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03362] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03363] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03364] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03365] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03366] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03367] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03368] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03369] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03370] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03371] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03372] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03373] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03374] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03375] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03376] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03377] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03378] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03379] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h066fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03380] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03381] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03382] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03383] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03384] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03385] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0670a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03386] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0670c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03387] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0670e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03388] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03389] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0671a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0671c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0671e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03390] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03391] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03392] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03393] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03394] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03395] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0672a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03396] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0672c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03397] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0672e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03398] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03399] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0673a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0673c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0673e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0674a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0674c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0674e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0675a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0675c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0675e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0676a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0676c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0676e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0677a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0677c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0677e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0678a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0678c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0678e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0679a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0679c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0679e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h067fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03400] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03401] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03402] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03403] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03404] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03405] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0680a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03406] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0680c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03407] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0680e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03408] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03409] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0681a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0681c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0681e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03410] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03411] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03412] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03413] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03414] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03415] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0682a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03416] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0682c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03417] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0682e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03418] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03419] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0683a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0683c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0683e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03420] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03421] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03422] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03423] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03424] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03425] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0684a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03426] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0684c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03427] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0684e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03428] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03429] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0685a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0685c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0685e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03430] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03431] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03432] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03433] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03434] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03435] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0686a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03436] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0686c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03437] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0686e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03438] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03439] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0687a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0687c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0687e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03440] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03441] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03442] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03443] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03444] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03445] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0688a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03446] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0688c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03447] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0688e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03448] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03449] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0689a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0689c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0689e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03450] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03451] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03452] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03453] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03454] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03455] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03456] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03457] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03458] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03459] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03460] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03461] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03462] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03463] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03464] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03465] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03466] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03467] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03468] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03469] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03470] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03471] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03472] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03473] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03474] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03475] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03476] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03477] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03478] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03479] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h068fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03480] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03481] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03482] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03483] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03484] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03485] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0690a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03486] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0690c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03487] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0690e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03488] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03489] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0691a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0691c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0691e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03490] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03491] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03492] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03493] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03494] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03495] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0692a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03496] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0692c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03497] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0692e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03498] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03499] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0693a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0693c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0693e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0694a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0694c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0694e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0695a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0695c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0695e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0696a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0696c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0696e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0697a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0697c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0697e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0698a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0698c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0698e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0699a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0699c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0699e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h069fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03500] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03501] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03502] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03503] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03504] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03505] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03506] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03507] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03508] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03509] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03510] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03511] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03512] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03513] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03514] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03515] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03516] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03517] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03518] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03519] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03520] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03521] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03522] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03523] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03524] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03525] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03526] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03527] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03528] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03529] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03530] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03531] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03532] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03533] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03534] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03535] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03536] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03537] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03538] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03539] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03540] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03541] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03542] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03543] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03544] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03545] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03546] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03547] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03548] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03549] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03550] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03551] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03552] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03553] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03554] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03555] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03556] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03557] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03558] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03559] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03560] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03561] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03562] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03563] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03564] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03565] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03566] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03567] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03568] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03569] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03570] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03571] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03572] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03573] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03574] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03575] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03576] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03577] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03578] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03579] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03580] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03581] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03582] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03583] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03584] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03585] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03586] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03587] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03588] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03589] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03590] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03591] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03592] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03593] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03594] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03595] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03596] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03597] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03598] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03599] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03600] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03601] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03602] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03603] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03604] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03605] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03606] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03607] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03608] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03609] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03610] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03611] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03612] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03613] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03614] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03615] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03616] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03617] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03618] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03619] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03620] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03621] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03622] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03623] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03624] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03625] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03626] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03627] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03628] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03629] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03630] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03631] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03632] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03633] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03634] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03635] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03636] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03637] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03638] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03639] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03640] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03641] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03642] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03643] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03644] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03645] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03646] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03647] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03648] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03649] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03650] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03651] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03652] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03653] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03654] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03655] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03656] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03657] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03658] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03659] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03660] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03661] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03662] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03663] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03664] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03665] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03666] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03667] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03668] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03669] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03670] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03671] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03672] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03673] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03674] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03675] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03676] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03677] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03678] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03679] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03680] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03681] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03682] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03683] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03684] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03685] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03686] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03687] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03688] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03689] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03690] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03691] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03692] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03693] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03694] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03695] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03696] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03697] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03698] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03699] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03700] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03701] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03702] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03703] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03704] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03705] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03706] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03707] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03708] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03709] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03710] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03711] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03712] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03713] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03714] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03715] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03716] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03717] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03718] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03719] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03720] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03721] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03722] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03723] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03724] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03725] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03726] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03727] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03728] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03729] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03730] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03731] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03732] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03733] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03734] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03735] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03736] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03737] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03738] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03739] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03740] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03741] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03742] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03743] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03744] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03745] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03746] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03747] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03748] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03749] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03750] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03751] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03752] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03753] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03754] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03755] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03756] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03757] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03758] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03759] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03760] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03761] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03762] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03763] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03764] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03765] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03766] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03767] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03768] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03769] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03770] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03771] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03772] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03773] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03774] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03775] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03776] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03777] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03778] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03779] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03780] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03781] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03782] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03783] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03784] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03785] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03786] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03787] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03788] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03789] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03790] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03791] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03792] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03793] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03794] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03795] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03796] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03797] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03798] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03799] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h06ffe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03800] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07000] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03801] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07002] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03802] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07004] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03803] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07006] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03804] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07008] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03805] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0700a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03806] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0700c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03807] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0700e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03808] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07010] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03809] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07012] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07014] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07016] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07018] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0701a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0701c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0701e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03810] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07020] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03811] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07022] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03812] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07024] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03813] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07026] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03814] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07028] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03815] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0702a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03816] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0702c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03817] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0702e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03818] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07030] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03819] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07032] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07034] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07036] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07038] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0703a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0703c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0703e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03820] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07040] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03821] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07042] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03822] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07044] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03823] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07046] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03824] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07048] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03825] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0704a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03826] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0704c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03827] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0704e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03828] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07050] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03829] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07052] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07054] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07056] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07058] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0705a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0705c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0705e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03830] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07060] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03831] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07062] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03832] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07064] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03833] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07066] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03834] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07068] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03835] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0706a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03836] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0706c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03837] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0706e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03838] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07070] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03839] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07072] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07074] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07076] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07078] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0707a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0707c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0707e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03840] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07080] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03841] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07082] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03842] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07084] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03843] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07086] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03844] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07088] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03845] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0708a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03846] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0708c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03847] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0708e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03848] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07090] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03849] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07092] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07094] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07096] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07098] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0709a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0709c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0709e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03850] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03851] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03852] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03853] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03854] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03855] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03856] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03857] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03858] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03859] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03860] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03861] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03862] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03863] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03864] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03865] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03866] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03867] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03868] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03869] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03870] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03871] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03872] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03873] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03874] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03875] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03876] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03877] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03878] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03879] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h070fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03880] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07100] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03881] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07102] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03882] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07104] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03883] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07106] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03884] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07108] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03885] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0710a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03886] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0710c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03887] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0710e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03888] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07110] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03889] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07112] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07114] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07116] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07118] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0711a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0711c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0711e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03890] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07120] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03891] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07122] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03892] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07124] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03893] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07126] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03894] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07128] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03895] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0712a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03896] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0712c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03897] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0712e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03898] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07130] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03899] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07132] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07134] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07136] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07138] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0713a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0713c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0713e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07140] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07142] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07144] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07146] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07148] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0714a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0714c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0714e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07150] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07152] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07154] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07156] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07158] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0715a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0715c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0715e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07160] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07162] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07164] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07166] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07168] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0716a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0716c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0716e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07170] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07172] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07174] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07176] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07178] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0717a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0717c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0717e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07180] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07182] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07184] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07186] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07188] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0718a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0718c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0718e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07190] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07192] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07194] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07196] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07198] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0719a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0719c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0719e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h071fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03900] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07200] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03901] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07202] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03902] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07204] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03903] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07206] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03904] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07208] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03905] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0720a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03906] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0720c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03907] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0720e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03908] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07210] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03909] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07212] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07214] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07216] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07218] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0721a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0721c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0721e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03910] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07220] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03911] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07222] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03912] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07224] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03913] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07226] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03914] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07228] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03915] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0722a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03916] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0722c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03917] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0722e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03918] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07230] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03919] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07232] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07234] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07236] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07238] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0723a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0723c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0723e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03920] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07240] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03921] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07242] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03922] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07244] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03923] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07246] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03924] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07248] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03925] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0724a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03926] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0724c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03927] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0724e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03928] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07250] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03929] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07252] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07254] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07256] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07258] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0725a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0725c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0725e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03930] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07260] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03931] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07262] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03932] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07264] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03933] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07266] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03934] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07268] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03935] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0726a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03936] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0726c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03937] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0726e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03938] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07270] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03939] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07272] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07274] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07276] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07278] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0727a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0727c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0727e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03940] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07280] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03941] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07282] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03942] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07284] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03943] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07286] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03944] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07288] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03945] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0728a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03946] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0728c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03947] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0728e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03948] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07290] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03949] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07292] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07294] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07296] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07298] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0729a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0729c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0729e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03950] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03951] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03952] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03953] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03954] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03955] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03956] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03957] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03958] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03959] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03960] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03961] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03962] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03963] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03964] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03965] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03966] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03967] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03968] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03969] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03970] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03971] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03972] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03973] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03974] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03975] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03976] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03977] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03978] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03979] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h072fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03980] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07300] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03981] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07302] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03982] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07304] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03983] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07306] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03984] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07308] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03985] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0730a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03986] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0730c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03987] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0730e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03988] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07310] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03989] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07312] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07314] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07316] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07318] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0731a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0731c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0731e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03990] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07320] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03991] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07322] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03992] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07324] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03993] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07326] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03994] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07328] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03995] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0732a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03996] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0732c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03997] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0732e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03998] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07330] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03999] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07332] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07334] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07336] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07338] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0733a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0733c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0733e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07340] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07342] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07344] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07346] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07348] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0734a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0734c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0734e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07350] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07352] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039aa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07354] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07356] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07358] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0735a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0735c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039af] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0735e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07360] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07362] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07364] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07366] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07368] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0736a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0736c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0736e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07370] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07372] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07374] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039bb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07376] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039bc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07378] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039bd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0737a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039be] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0737c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039bf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0737e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07380] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07382] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07384] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07386] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07388] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0738a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0738c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0738e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07390] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07392] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07394] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039cb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07396] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039cc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07398] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039cd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0739a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0739c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039cf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0739e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039da] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039db] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039dc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039dd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039de] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039df] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039eb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h073fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07400] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07402] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07404] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07406] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07408] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0740a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0740c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0740e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07410] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07412] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07414] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07416] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07418] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0741a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0741c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0741e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07420] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07422] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07424] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07426] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07428] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0742a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0742c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0742e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07430] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07432] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07434] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07436] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07438] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0743a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0743c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0743e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07440] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07442] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07444] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07446] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07448] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0744a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0744c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0744e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07450] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07452] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07454] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07456] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07458] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0745a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0745c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0745e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07460] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07462] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07464] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07466] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07468] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0746a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0746c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0746e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07470] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07472] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07474] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07476] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07478] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0747a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0747c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0747e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07480] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07482] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07484] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07486] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07488] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0748a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0748c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0748e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07490] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07492] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07494] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07496] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07498] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0749a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0749c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0749e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h074fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07500] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07502] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07504] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07506] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07508] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0750a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0750c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0750e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07510] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07512] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07514] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07516] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07518] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0751a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0751c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0751e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07520] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07522] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07524] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07526] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07528] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0752a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0752c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0752e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07530] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07532] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07534] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07536] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07538] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0753a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0753c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0753e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07540] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07542] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07544] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07546] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07548] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0754a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0754c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0754e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07550] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07552] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07554] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07556] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07558] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0755a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0755c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0755e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07560] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07562] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07564] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07566] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07568] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0756a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0756c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0756e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07570] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07572] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07574] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07576] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07578] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0757a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0757c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0757e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07580] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07582] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07584] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07586] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07588] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0758a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0758c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0758e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07590] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07592] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07594] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03acb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07596] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03acc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07598] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03acd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0759a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ace] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0759c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03acf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0759e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ada] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03adb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03adc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03add] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ade] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03adf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h075fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07600] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07602] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07604] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07606] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07608] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0760a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0760c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0760e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07610] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07612] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07614] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07616] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07618] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0761a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0761c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0761e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07620] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07622] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07624] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07626] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07628] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0762a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0762c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0762e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07630] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07632] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07634] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07636] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07638] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0763a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0763c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0763e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07640] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07642] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07644] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07646] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07648] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0764a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0764c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0764e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07650] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07652] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07654] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07656] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07658] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0765a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0765c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0765e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07660] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07662] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07664] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07666] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07668] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0766a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0766c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0766e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07670] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07672] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07674] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07676] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07678] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0767a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0767c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0767e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07680] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07682] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07684] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07686] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07688] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0768a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0768c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0768e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07690] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07692] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07694] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07696] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07698] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0769a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0769c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0769e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h076fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07700] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07702] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07704] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07706] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07708] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0770a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0770c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0770e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07710] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07712] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07714] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07716] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07718] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0771a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0771c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0771e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07720] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07722] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07724] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07726] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07728] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0772a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0772c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0772e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07730] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07732] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07734] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07736] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07738] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0773a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0773c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0773e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07740] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07742] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07744] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07746] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07748] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0774a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0774c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0774e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07750] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07752] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03baa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07754] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07756] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07758] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0775a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0775c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03baf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0775e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07760] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07762] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07764] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07766] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07768] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0776a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0776c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0776e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07770] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07772] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07774] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07776] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07778] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0777a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0777c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0777e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07780] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07782] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07784] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07786] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07788] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0778a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0778c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0778e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07790] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07792] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07794] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07796] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07798] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0779a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0779c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0779e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03beb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h077fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07800] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07802] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07804] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07806] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07808] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0780a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0780c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0780e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07810] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07812] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07814] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07816] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07818] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0781a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0781c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0781e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07820] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07822] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07824] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07826] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07828] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0782a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0782c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0782e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07830] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07832] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07834] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07836] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07838] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0783a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0783c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0783e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07840] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07842] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07844] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07846] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07848] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0784a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0784c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0784e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07850] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07852] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07854] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07856] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07858] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0785a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0785c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0785e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07860] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07862] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07864] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07866] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07868] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0786a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0786c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0786e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07870] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07872] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07874] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07876] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07878] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0787a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0787c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0787e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07880] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07882] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07884] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07886] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07888] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0788a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0788c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0788e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07890] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07892] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07894] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07896] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07898] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0789a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0789c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0789e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h078fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07900] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07902] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07904] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07906] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07908] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0790a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0790c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0790e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07910] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07912] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07914] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07916] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07918] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0791a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0791c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0791e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07920] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07922] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07924] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07926] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07928] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0792a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0792c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0792e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07930] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07932] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07934] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07936] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07938] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0793a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0793c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0793e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07940] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07942] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07944] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07946] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07948] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0794a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0794c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0794e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07950] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07952] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03caa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07954] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07956] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07958] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0795a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0795c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03caf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0795e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07960] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07962] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07964] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07966] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07968] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0796a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0796c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0796e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07970] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07972] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07974] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07976] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07978] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0797a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0797c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0797e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07980] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07982] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07984] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07986] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07988] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0798a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0798c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0798e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07990] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07992] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07994] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ccb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07996] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ccc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07998] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ccd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0799a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0799c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ccf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h0799e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079a0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079a2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079a4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079a6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079a8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079aa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079b0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079b2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079b4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079b6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079b8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079bc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079be] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079c0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079c2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079c4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079c6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079c8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079cc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079d0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079d2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079d4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ceb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079d6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079d8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ced] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079da] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079dc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079de] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079e0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079e2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079e4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079e6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079e8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079ee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079f0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079f2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079f4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079f6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079f8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079fa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079fc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h079fe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07a9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ab0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ab2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ab4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ab6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ab8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07abc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07abe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ac0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ac2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ac4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ac6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ac8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07acc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ace] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ad0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ad2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ad4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ad6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ad8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ada] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07adc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ade] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ae0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ae2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ae4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ae6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ae8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07aee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07af0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07af2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07af4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07af6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07af8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07afa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07afc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07afe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03daa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03daf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07b9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ba0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ba2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ba4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ba6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ba8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07baa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ddb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ddc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ddd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ddf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03deb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ded] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03def] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07be0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07be2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07be4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07be6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07be8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07bfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07c9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ca0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ca2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ca4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ca6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ca8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07caa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ccc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ce0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ce2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ce4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ce6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ce8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cf0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cf2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cf4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cf6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cf8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07cfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eaa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ead] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eaf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ecb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ecc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ecd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ece] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ecf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07d9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07da0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07da2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07da4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07da6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07da8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07daa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07db0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07db2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07db4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03edb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07db6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03edc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07db8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03edd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ede] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03edf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eeb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ddc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07de0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07de2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07de4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07de6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07de8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07df0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07df2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07df4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07df6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07df8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dfa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dfc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07dfe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f00] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f01] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f02] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f03] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f04] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f05] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f06] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f07] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f08] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f09] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f10] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f11] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f12] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f13] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f14] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f15] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f16] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f17] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f18] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f19] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f20] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f21] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f22] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f23] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f24] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f25] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f26] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f27] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f28] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f29] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f30] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f31] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f32] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f33] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f34] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f35] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f36] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f37] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f38] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f39] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f40] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f41] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f42] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f43] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f44] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f45] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f46] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f47] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f48] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f49] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07e9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f50] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ea0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f51] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ea2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f52] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ea4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f53] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ea6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f54] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ea8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f55] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eaa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f56] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f57] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f58] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f59] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ebc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ebe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f60] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ec0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f61] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ec2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f62] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ec4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f63] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ec6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f64] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ec8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f65] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f66] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ecc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f67] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ece] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f68] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ed0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f69] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ed2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ed4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ed6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ed8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07edc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ede] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f70] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ee0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f71] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ee2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f72] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ee4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f73] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ee6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f74] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ee8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f75] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f76] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f77] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07eee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f78] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ef0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f79] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ef2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ef4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ef6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ef8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07efa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07efc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07efe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f80] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f00] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f81] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f02] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f82] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f04] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f83] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f06] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f84] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f08] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f85] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f0a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f86] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f0c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f87] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f0e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f88] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f10] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f89] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f12] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f14] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f16] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f18] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f1a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f1c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f1e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f90] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f20] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f91] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f22] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f92] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f24] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f93] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f26] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f94] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f28] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f95] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f2a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f96] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f2c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f97] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f2e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f98] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f30] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f99] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f32] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9a] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f34] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9b] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f36] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9c] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f38] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9d] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f3a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9e] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f3c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9f] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f3e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f40] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f42] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f44] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f46] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f48] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f4a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f4c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f4e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f50] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f52] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03faa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f54] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fab] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f56] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fac] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f58] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fad] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f5a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fae] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f5c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03faf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f5e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f60] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f62] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f64] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f66] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f68] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f6a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f6c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f6e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f70] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f72] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fba] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f74] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f76] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f78] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f7a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f7c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f7e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f80] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f82] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f84] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f86] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f88] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f8a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f8c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f8e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f90] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f92] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fca] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f94] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fcb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f96] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fcc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f98] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fcd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f9a] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fce] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f9c] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fcf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07f9e] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fa0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fa2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fa4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fa6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fa8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07faa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fac] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fae] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fb0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fb2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fda] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fb4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fdb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fb6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fdc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fb8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fdd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fba] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fde] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fbc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fdf] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fbe] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fc0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fc2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fc4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fc6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fc8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fca] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fcc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fce] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fd0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fd2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fea] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fd4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03feb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fd6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fec] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fd8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fed] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fda] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fee] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fdc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fef] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fde] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff0] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fe0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff1] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fe2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff2] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fe4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff3] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fe6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff4] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fe8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff5] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fea] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff6] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fec] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff7] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07fee] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff8] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ff0] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff9] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ff2] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffa] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ff4] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffb] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ff6] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffc] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ff8] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffd] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ffa] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffe] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ffc] ;
//end
//always_comb begin // 
               Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fff] =  I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1['h07ffe] ;
//end
