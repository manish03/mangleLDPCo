 reg  ['h1f:0] [$clog2('h7000+1)-1:0] If72de6675c42172560d5d150642f3da8 ;
