              Id8535704c02d21b31bba0f979b865ce2 = 
          (!flogtanh_sel[7]) ? 
                       Ida9cf0ff6fe9afcde8fb6e10f4a2a9a3: 
                       I9ff622ac8ef93a7d8d1bf5f91cd0f972;
              I4b9150498657596ba1fcdcf43bc2644b = 
          (!flogtanh_sel[7]) ? 
                       I35a5875790032fa907cbfff6be72a604: 
                       Ica42b16ad8703e0088757d8a95c17578;
