 reg  ['hfff:0] [$clog2('h7000+1)-1:0] I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e ;
