//`include "GF2_LDPC_flogtanh_0x00005_assign_inc.sv"
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00000] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00000] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00001] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00001] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00002] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00003] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00002] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00004] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00005] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00003] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00006] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00007] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00004] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00008] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00009] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00005] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0000a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0000b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00006] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0000c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0000d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00007] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0000e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0000f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00008] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00010] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00011] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00009] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00012] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00013] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0000a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00014] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00015] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0000b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00016] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00017] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0000c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00018] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00019] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0000d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0001a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0001b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0000e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0001c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0001d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0000f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0001e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0001f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00010] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00020] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00021] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00011] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00022] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00023] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00012] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00024] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00025] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00013] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00026] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00027] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00014] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00028] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00029] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00015] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0002a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0002b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00016] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0002c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0002d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00017] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0002e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0002f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00018] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00030] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00031] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00019] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00032] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00033] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0001a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00034] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00035] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0001b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00036] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00037] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0001c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00038] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00039] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0001d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0003a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0003b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0001e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0003c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0003d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0001f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0003e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0003f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00020] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00040] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00041] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00021] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00042] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00043] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00022] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00044] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00045] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00023] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00046] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00047] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00024] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00048] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00049] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00025] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0004a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0004b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00026] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0004c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0004d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00027] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0004e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0004f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00028] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00050] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00051] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00029] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00052] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00053] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0002a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00054] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00055] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0002b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00056] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00057] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0002c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00058] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00059] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0002d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0005a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0005b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0002e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0005c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0005d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0002f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0005e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0005f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00030] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00060] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00061] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00031] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00062] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00063] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00032] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00064] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00065] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00033] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00066] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00067] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00034] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00068] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00069] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00035] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0006a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0006b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00036] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0006c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0006d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00037] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0006e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0006f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00038] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00070] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00071] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00039] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00072] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00073] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0003a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00074] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00075] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0003b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00076] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00077] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0003c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00078] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00079] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0003d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0007a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0007b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0003e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0007c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0007d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0003f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0007e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0007f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00040] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00080] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00081] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00041] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00082] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00083] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00042] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00084] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00085] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00043] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00086] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00087] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00044] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00088] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00089] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00045] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0008a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0008b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00046] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0008c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0008d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00047] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0008e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0008f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00048] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00090] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00091] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00049] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00092] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00093] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0004a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00094] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00095] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0004b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00096] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00097] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0004c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00098] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00099] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0004d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0009a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0009b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0004e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0009c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0009d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0004f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0009e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0009f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00050] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000a0] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000a1] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00051] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000a2] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000a3] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00052] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000a4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000a5] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00053] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000a6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000a7] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00054] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000a8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000a9] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00055] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000aa] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000ab] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00056] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ac] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000ad] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00057] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ae] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000af] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00058] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000b0] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000b1] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00059] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000b2] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000b3] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0005a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000b4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000b5] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0005b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000b6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000b7] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0005c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000b8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000b9] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0005d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ba] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000bb] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0005e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000bc] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000bd] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0005f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000be] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000bf] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00060] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000c0] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000c1] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00061] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000c2] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000c3] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00062] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000c4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000c5] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00063] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000c6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000c7] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00064] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000c8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000c9] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00065] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ca] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000cb] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00066] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000cc] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000cd] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00067] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ce] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000cf] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00068] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000d0] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000d1] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00069] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000d2] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000d3] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0006a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000d4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000d5] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0006b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000d6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000d7] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0006c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000d8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000d9] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0006d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000da] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000db] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0006e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000dc] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000dd] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0006f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000de] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000df] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00070] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000e0] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000e1] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00071] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000e2] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000e3] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00072] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000e4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000e5] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00073] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000e6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000e7] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00074] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000e8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000e9] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00075] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ea] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000eb] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00076] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ec] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000ed] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00077] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000ee] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000ef] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00078] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000f0] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000f1] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00079] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000f2] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000f3] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0007a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000f4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000f5] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0007b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000f6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000f7] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0007c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000f8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000f9] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0007d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000fa] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000fb] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0007e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000fc] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000fd] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0007f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h000fe] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h000ff] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00080] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00100] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00101] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00081] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00102] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00103] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00082] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00104] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00105] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00083] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00106] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00107] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00084] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00108] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00109] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00085] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0010a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0010b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00086] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0010c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0010d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00087] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0010e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0010f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00088] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00110] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00111] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00089] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00112] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00113] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0008a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00114] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00115] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0008b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00116] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00117] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0008c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00118] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00119] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0008d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0011a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0011b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0008e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0011c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0011d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0008f] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0011e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0011f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00090] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00120] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00121] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00091] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00122] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00123] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00092] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00124] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00125] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00093] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00126] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00127] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00094] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00128] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00129] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00095] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0012a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0012b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00096] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0012c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0012d] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00097] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0012e] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0012f] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00098] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00130] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00131] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00099] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00132] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00133] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0009a] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00134] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00135] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0009b] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00136] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00137] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0009c] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00138] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00139] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0009d] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0013a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0013b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h0009e] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0013c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0013d] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0009f] =  I0310077d53ae4ed9904df42e3f81c634['h0013e] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a0] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00140] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00141] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a1] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00142] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00143] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a2] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00144] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00145] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a3] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00146] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00147] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000a4] =  I0310077d53ae4ed9904df42e3f81c634['h00148] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a5] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0014a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0014b] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a6] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0014c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0014d] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000a7] =  I0310077d53ae4ed9904df42e3f81c634['h0014e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000a8] =  I0310077d53ae4ed9904df42e3f81c634['h00150] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000a9] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00152] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00153] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000aa] =  I0310077d53ae4ed9904df42e3f81c634['h00154] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000ab] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00156] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00157] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000ac] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00158] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00159] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ad] =  I0310077d53ae4ed9904df42e3f81c634['h0015a] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000ae] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0015c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0015d] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000af] =  I0310077d53ae4ed9904df42e3f81c634['h0015e] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000b0] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00160] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00161] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000b1] =  I0310077d53ae4ed9904df42e3f81c634['h00162] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000b2] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00164] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00165] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000b3] =  I0310077d53ae4ed9904df42e3f81c634['h00166] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000b4] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00168] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00169] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000b5] =  I0310077d53ae4ed9904df42e3f81c634['h0016a] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000b6] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0016c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0016d] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000b7] =  I0310077d53ae4ed9904df42e3f81c634['h0016e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000b8] =  I0310077d53ae4ed9904df42e3f81c634['h00170] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000b9] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00172] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00173] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ba] =  I0310077d53ae4ed9904df42e3f81c634['h00174] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000bb] =  I0310077d53ae4ed9904df42e3f81c634['h00176] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000bc] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00178] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00179] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000bd] =  I0310077d53ae4ed9904df42e3f81c634['h0017a] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000be] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0017c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0017d] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000bf] =  I0310077d53ae4ed9904df42e3f81c634['h0017e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c0] =  I0310077d53ae4ed9904df42e3f81c634['h00180] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c1] =  I0310077d53ae4ed9904df42e3f81c634['h00182] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000c2] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00184] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00185] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c3] =  I0310077d53ae4ed9904df42e3f81c634['h00186] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c4] =  I0310077d53ae4ed9904df42e3f81c634['h00188] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000c5] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0018a] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0018b] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c6] =  I0310077d53ae4ed9904df42e3f81c634['h0018c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c7] =  I0310077d53ae4ed9904df42e3f81c634['h0018e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000c8] =  I0310077d53ae4ed9904df42e3f81c634['h00190] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000c9] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00192] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00193] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ca] =  I0310077d53ae4ed9904df42e3f81c634['h00194] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000cb] =  I0310077d53ae4ed9904df42e3f81c634['h00196] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000cc] =  I0310077d53ae4ed9904df42e3f81c634['h00198] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000cd] =  I0310077d53ae4ed9904df42e3f81c634['h0019a] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000ce] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h0019c] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h0019d] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000cf] =  I0310077d53ae4ed9904df42e3f81c634['h0019e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d0] =  I0310077d53ae4ed9904df42e3f81c634['h001a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d1] =  I0310077d53ae4ed9904df42e3f81c634['h001a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d2] =  I0310077d53ae4ed9904df42e3f81c634['h001a4] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000d3] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h001a6] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h001a7] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d4] =  I0310077d53ae4ed9904df42e3f81c634['h001a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d5] =  I0310077d53ae4ed9904df42e3f81c634['h001aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d6] =  I0310077d53ae4ed9904df42e3f81c634['h001ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d7] =  I0310077d53ae4ed9904df42e3f81c634['h001ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d8] =  I0310077d53ae4ed9904df42e3f81c634['h001b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000d9] =  I0310077d53ae4ed9904df42e3f81c634['h001b2] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000da] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h001b4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h001b5] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000db] =  I0310077d53ae4ed9904df42e3f81c634['h001b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000dc] =  I0310077d53ae4ed9904df42e3f81c634['h001b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000dd] =  I0310077d53ae4ed9904df42e3f81c634['h001ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000de] =  I0310077d53ae4ed9904df42e3f81c634['h001bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000df] =  I0310077d53ae4ed9904df42e3f81c634['h001be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e0] =  I0310077d53ae4ed9904df42e3f81c634['h001c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e1] =  I0310077d53ae4ed9904df42e3f81c634['h001c2] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000e2] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h001c4] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h001c5] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e3] =  I0310077d53ae4ed9904df42e3f81c634['h001c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e4] =  I0310077d53ae4ed9904df42e3f81c634['h001c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e5] =  I0310077d53ae4ed9904df42e3f81c634['h001ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e6] =  I0310077d53ae4ed9904df42e3f81c634['h001cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e7] =  I0310077d53ae4ed9904df42e3f81c634['h001ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e8] =  I0310077d53ae4ed9904df42e3f81c634['h001d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000e9] =  I0310077d53ae4ed9904df42e3f81c634['h001d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ea] =  I0310077d53ae4ed9904df42e3f81c634['h001d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000eb] =  I0310077d53ae4ed9904df42e3f81c634['h001d6] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000ec] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h001d8] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h001d9] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ed] =  I0310077d53ae4ed9904df42e3f81c634['h001da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ee] =  I0310077d53ae4ed9904df42e3f81c634['h001dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ef] =  I0310077d53ae4ed9904df42e3f81c634['h001de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f0] =  I0310077d53ae4ed9904df42e3f81c634['h001e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f1] =  I0310077d53ae4ed9904df42e3f81c634['h001e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f2] =  I0310077d53ae4ed9904df42e3f81c634['h001e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f3] =  I0310077d53ae4ed9904df42e3f81c634['h001e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f4] =  I0310077d53ae4ed9904df42e3f81c634['h001e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f5] =  I0310077d53ae4ed9904df42e3f81c634['h001ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f6] =  I0310077d53ae4ed9904df42e3f81c634['h001ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f7] =  I0310077d53ae4ed9904df42e3f81c634['h001ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f8] =  I0310077d53ae4ed9904df42e3f81c634['h001f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000f9] =  I0310077d53ae4ed9904df42e3f81c634['h001f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000fa] =  I0310077d53ae4ed9904df42e3f81c634['h001f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000fb] =  I0310077d53ae4ed9904df42e3f81c634['h001f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000fc] =  I0310077d53ae4ed9904df42e3f81c634['h001f8] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h000fd] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h001fa] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h001fb] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000fe] =  I0310077d53ae4ed9904df42e3f81c634['h001fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h000ff] =  I0310077d53ae4ed9904df42e3f81c634['h001fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00100] =  I0310077d53ae4ed9904df42e3f81c634['h00200] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00101] =  I0310077d53ae4ed9904df42e3f81c634['h00202] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00102] =  I0310077d53ae4ed9904df42e3f81c634['h00204] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00103] =  I0310077d53ae4ed9904df42e3f81c634['h00206] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00104] =  I0310077d53ae4ed9904df42e3f81c634['h00208] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00105] =  I0310077d53ae4ed9904df42e3f81c634['h0020a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00106] =  I0310077d53ae4ed9904df42e3f81c634['h0020c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00107] =  I0310077d53ae4ed9904df42e3f81c634['h0020e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00108] =  I0310077d53ae4ed9904df42e3f81c634['h00210] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00109] =  I0310077d53ae4ed9904df42e3f81c634['h00212] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0010a] =  I0310077d53ae4ed9904df42e3f81c634['h00214] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0010b] =  I0310077d53ae4ed9904df42e3f81c634['h00216] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0010c] =  I0310077d53ae4ed9904df42e3f81c634['h00218] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0010d] =  I0310077d53ae4ed9904df42e3f81c634['h0021a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0010e] =  I0310077d53ae4ed9904df42e3f81c634['h0021c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0010f] =  I0310077d53ae4ed9904df42e3f81c634['h0021e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00110] =  I0310077d53ae4ed9904df42e3f81c634['h00220] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00111] =  I0310077d53ae4ed9904df42e3f81c634['h00222] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00112] =  I0310077d53ae4ed9904df42e3f81c634['h00224] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00113] =  I0310077d53ae4ed9904df42e3f81c634['h00226] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00114] =  I0310077d53ae4ed9904df42e3f81c634['h00228] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00115] =  I0310077d53ae4ed9904df42e3f81c634['h0022a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00116] =  I0310077d53ae4ed9904df42e3f81c634['h0022c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00117] =  I0310077d53ae4ed9904df42e3f81c634['h0022e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00118] =  I0310077d53ae4ed9904df42e3f81c634['h00230] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00119] =  I0310077d53ae4ed9904df42e3f81c634['h00232] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0011a] =  I0310077d53ae4ed9904df42e3f81c634['h00234] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0011b] =  I0310077d53ae4ed9904df42e3f81c634['h00236] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0011c] =  I0310077d53ae4ed9904df42e3f81c634['h00238] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0011d] =  I0310077d53ae4ed9904df42e3f81c634['h0023a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0011e] =  I0310077d53ae4ed9904df42e3f81c634['h0023c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0011f] =  I0310077d53ae4ed9904df42e3f81c634['h0023e] ;
//end
//always_comb begin
              Ifcca41d795dde8a35d1654b9520c92e7['h00120] = 
          (!flogtanh_sel['h00005]) ? 
                       I0310077d53ae4ed9904df42e3f81c634['h00240] : //%
                       I0310077d53ae4ed9904df42e3f81c634['h00241] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00121] =  I0310077d53ae4ed9904df42e3f81c634['h00242] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00122] =  I0310077d53ae4ed9904df42e3f81c634['h00244] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00123] =  I0310077d53ae4ed9904df42e3f81c634['h00246] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00124] =  I0310077d53ae4ed9904df42e3f81c634['h00248] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00125] =  I0310077d53ae4ed9904df42e3f81c634['h0024a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00126] =  I0310077d53ae4ed9904df42e3f81c634['h0024c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00127] =  I0310077d53ae4ed9904df42e3f81c634['h0024e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00128] =  I0310077d53ae4ed9904df42e3f81c634['h00250] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00129] =  I0310077d53ae4ed9904df42e3f81c634['h00252] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0012a] =  I0310077d53ae4ed9904df42e3f81c634['h00254] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0012b] =  I0310077d53ae4ed9904df42e3f81c634['h00256] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0012c] =  I0310077d53ae4ed9904df42e3f81c634['h00258] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0012d] =  I0310077d53ae4ed9904df42e3f81c634['h0025a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0012e] =  I0310077d53ae4ed9904df42e3f81c634['h0025c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0012f] =  I0310077d53ae4ed9904df42e3f81c634['h0025e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00130] =  I0310077d53ae4ed9904df42e3f81c634['h00260] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00131] =  I0310077d53ae4ed9904df42e3f81c634['h00262] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00132] =  I0310077d53ae4ed9904df42e3f81c634['h00264] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00133] =  I0310077d53ae4ed9904df42e3f81c634['h00266] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00134] =  I0310077d53ae4ed9904df42e3f81c634['h00268] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00135] =  I0310077d53ae4ed9904df42e3f81c634['h0026a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00136] =  I0310077d53ae4ed9904df42e3f81c634['h0026c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00137] =  I0310077d53ae4ed9904df42e3f81c634['h0026e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00138] =  I0310077d53ae4ed9904df42e3f81c634['h00270] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00139] =  I0310077d53ae4ed9904df42e3f81c634['h00272] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0013a] =  I0310077d53ae4ed9904df42e3f81c634['h00274] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0013b] =  I0310077d53ae4ed9904df42e3f81c634['h00276] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0013c] =  I0310077d53ae4ed9904df42e3f81c634['h00278] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0013d] =  I0310077d53ae4ed9904df42e3f81c634['h0027a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0013e] =  I0310077d53ae4ed9904df42e3f81c634['h0027c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0013f] =  I0310077d53ae4ed9904df42e3f81c634['h0027e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00140] =  I0310077d53ae4ed9904df42e3f81c634['h00280] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00141] =  I0310077d53ae4ed9904df42e3f81c634['h00282] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00142] =  I0310077d53ae4ed9904df42e3f81c634['h00284] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00143] =  I0310077d53ae4ed9904df42e3f81c634['h00286] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00144] =  I0310077d53ae4ed9904df42e3f81c634['h00288] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00145] =  I0310077d53ae4ed9904df42e3f81c634['h0028a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00146] =  I0310077d53ae4ed9904df42e3f81c634['h0028c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00147] =  I0310077d53ae4ed9904df42e3f81c634['h0028e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00148] =  I0310077d53ae4ed9904df42e3f81c634['h00290] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00149] =  I0310077d53ae4ed9904df42e3f81c634['h00292] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0014a] =  I0310077d53ae4ed9904df42e3f81c634['h00294] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0014b] =  I0310077d53ae4ed9904df42e3f81c634['h00296] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0014c] =  I0310077d53ae4ed9904df42e3f81c634['h00298] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0014d] =  I0310077d53ae4ed9904df42e3f81c634['h0029a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0014e] =  I0310077d53ae4ed9904df42e3f81c634['h0029c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0014f] =  I0310077d53ae4ed9904df42e3f81c634['h0029e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00150] =  I0310077d53ae4ed9904df42e3f81c634['h002a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00151] =  I0310077d53ae4ed9904df42e3f81c634['h002a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00152] =  I0310077d53ae4ed9904df42e3f81c634['h002a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00153] =  I0310077d53ae4ed9904df42e3f81c634['h002a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00154] =  I0310077d53ae4ed9904df42e3f81c634['h002a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00155] =  I0310077d53ae4ed9904df42e3f81c634['h002aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00156] =  I0310077d53ae4ed9904df42e3f81c634['h002ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00157] =  I0310077d53ae4ed9904df42e3f81c634['h002ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00158] =  I0310077d53ae4ed9904df42e3f81c634['h002b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00159] =  I0310077d53ae4ed9904df42e3f81c634['h002b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0015a] =  I0310077d53ae4ed9904df42e3f81c634['h002b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0015b] =  I0310077d53ae4ed9904df42e3f81c634['h002b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0015c] =  I0310077d53ae4ed9904df42e3f81c634['h002b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0015d] =  I0310077d53ae4ed9904df42e3f81c634['h002ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0015e] =  I0310077d53ae4ed9904df42e3f81c634['h002bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0015f] =  I0310077d53ae4ed9904df42e3f81c634['h002be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00160] =  I0310077d53ae4ed9904df42e3f81c634['h002c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00161] =  I0310077d53ae4ed9904df42e3f81c634['h002c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00162] =  I0310077d53ae4ed9904df42e3f81c634['h002c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00163] =  I0310077d53ae4ed9904df42e3f81c634['h002c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00164] =  I0310077d53ae4ed9904df42e3f81c634['h002c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00165] =  I0310077d53ae4ed9904df42e3f81c634['h002ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00166] =  I0310077d53ae4ed9904df42e3f81c634['h002cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00167] =  I0310077d53ae4ed9904df42e3f81c634['h002ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00168] =  I0310077d53ae4ed9904df42e3f81c634['h002d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00169] =  I0310077d53ae4ed9904df42e3f81c634['h002d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0016a] =  I0310077d53ae4ed9904df42e3f81c634['h002d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0016b] =  I0310077d53ae4ed9904df42e3f81c634['h002d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0016c] =  I0310077d53ae4ed9904df42e3f81c634['h002d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0016d] =  I0310077d53ae4ed9904df42e3f81c634['h002da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0016e] =  I0310077d53ae4ed9904df42e3f81c634['h002dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0016f] =  I0310077d53ae4ed9904df42e3f81c634['h002de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00170] =  I0310077d53ae4ed9904df42e3f81c634['h002e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00171] =  I0310077d53ae4ed9904df42e3f81c634['h002e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00172] =  I0310077d53ae4ed9904df42e3f81c634['h002e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00173] =  I0310077d53ae4ed9904df42e3f81c634['h002e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00174] =  I0310077d53ae4ed9904df42e3f81c634['h002e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00175] =  I0310077d53ae4ed9904df42e3f81c634['h002ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00176] =  I0310077d53ae4ed9904df42e3f81c634['h002ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00177] =  I0310077d53ae4ed9904df42e3f81c634['h002ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00178] =  I0310077d53ae4ed9904df42e3f81c634['h002f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00179] =  I0310077d53ae4ed9904df42e3f81c634['h002f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0017a] =  I0310077d53ae4ed9904df42e3f81c634['h002f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0017b] =  I0310077d53ae4ed9904df42e3f81c634['h002f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0017c] =  I0310077d53ae4ed9904df42e3f81c634['h002f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0017d] =  I0310077d53ae4ed9904df42e3f81c634['h002fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0017e] =  I0310077d53ae4ed9904df42e3f81c634['h002fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0017f] =  I0310077d53ae4ed9904df42e3f81c634['h002fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00180] =  I0310077d53ae4ed9904df42e3f81c634['h00300] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00181] =  I0310077d53ae4ed9904df42e3f81c634['h00302] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00182] =  I0310077d53ae4ed9904df42e3f81c634['h00304] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00183] =  I0310077d53ae4ed9904df42e3f81c634['h00306] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00184] =  I0310077d53ae4ed9904df42e3f81c634['h00308] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00185] =  I0310077d53ae4ed9904df42e3f81c634['h0030a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00186] =  I0310077d53ae4ed9904df42e3f81c634['h0030c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00187] =  I0310077d53ae4ed9904df42e3f81c634['h0030e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00188] =  I0310077d53ae4ed9904df42e3f81c634['h00310] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00189] =  I0310077d53ae4ed9904df42e3f81c634['h00312] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0018a] =  I0310077d53ae4ed9904df42e3f81c634['h00314] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0018b] =  I0310077d53ae4ed9904df42e3f81c634['h00316] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0018c] =  I0310077d53ae4ed9904df42e3f81c634['h00318] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0018d] =  I0310077d53ae4ed9904df42e3f81c634['h0031a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0018e] =  I0310077d53ae4ed9904df42e3f81c634['h0031c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0018f] =  I0310077d53ae4ed9904df42e3f81c634['h0031e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00190] =  I0310077d53ae4ed9904df42e3f81c634['h00320] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00191] =  I0310077d53ae4ed9904df42e3f81c634['h00322] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00192] =  I0310077d53ae4ed9904df42e3f81c634['h00324] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00193] =  I0310077d53ae4ed9904df42e3f81c634['h00326] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00194] =  I0310077d53ae4ed9904df42e3f81c634['h00328] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00195] =  I0310077d53ae4ed9904df42e3f81c634['h0032a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00196] =  I0310077d53ae4ed9904df42e3f81c634['h0032c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00197] =  I0310077d53ae4ed9904df42e3f81c634['h0032e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00198] =  I0310077d53ae4ed9904df42e3f81c634['h00330] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00199] =  I0310077d53ae4ed9904df42e3f81c634['h00332] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0019a] =  I0310077d53ae4ed9904df42e3f81c634['h00334] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0019b] =  I0310077d53ae4ed9904df42e3f81c634['h00336] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0019c] =  I0310077d53ae4ed9904df42e3f81c634['h00338] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0019d] =  I0310077d53ae4ed9904df42e3f81c634['h0033a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0019e] =  I0310077d53ae4ed9904df42e3f81c634['h0033c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0019f] =  I0310077d53ae4ed9904df42e3f81c634['h0033e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a0] =  I0310077d53ae4ed9904df42e3f81c634['h00340] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a1] =  I0310077d53ae4ed9904df42e3f81c634['h00342] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a2] =  I0310077d53ae4ed9904df42e3f81c634['h00344] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a3] =  I0310077d53ae4ed9904df42e3f81c634['h00346] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a4] =  I0310077d53ae4ed9904df42e3f81c634['h00348] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a5] =  I0310077d53ae4ed9904df42e3f81c634['h0034a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a6] =  I0310077d53ae4ed9904df42e3f81c634['h0034c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a7] =  I0310077d53ae4ed9904df42e3f81c634['h0034e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a8] =  I0310077d53ae4ed9904df42e3f81c634['h00350] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001a9] =  I0310077d53ae4ed9904df42e3f81c634['h00352] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001aa] =  I0310077d53ae4ed9904df42e3f81c634['h00354] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ab] =  I0310077d53ae4ed9904df42e3f81c634['h00356] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ac] =  I0310077d53ae4ed9904df42e3f81c634['h00358] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ad] =  I0310077d53ae4ed9904df42e3f81c634['h0035a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ae] =  I0310077d53ae4ed9904df42e3f81c634['h0035c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001af] =  I0310077d53ae4ed9904df42e3f81c634['h0035e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b0] =  I0310077d53ae4ed9904df42e3f81c634['h00360] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b1] =  I0310077d53ae4ed9904df42e3f81c634['h00362] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b2] =  I0310077d53ae4ed9904df42e3f81c634['h00364] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b3] =  I0310077d53ae4ed9904df42e3f81c634['h00366] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b4] =  I0310077d53ae4ed9904df42e3f81c634['h00368] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b5] =  I0310077d53ae4ed9904df42e3f81c634['h0036a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b6] =  I0310077d53ae4ed9904df42e3f81c634['h0036c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b7] =  I0310077d53ae4ed9904df42e3f81c634['h0036e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b8] =  I0310077d53ae4ed9904df42e3f81c634['h00370] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001b9] =  I0310077d53ae4ed9904df42e3f81c634['h00372] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ba] =  I0310077d53ae4ed9904df42e3f81c634['h00374] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001bb] =  I0310077d53ae4ed9904df42e3f81c634['h00376] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001bc] =  I0310077d53ae4ed9904df42e3f81c634['h00378] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001bd] =  I0310077d53ae4ed9904df42e3f81c634['h0037a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001be] =  I0310077d53ae4ed9904df42e3f81c634['h0037c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001bf] =  I0310077d53ae4ed9904df42e3f81c634['h0037e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c0] =  I0310077d53ae4ed9904df42e3f81c634['h00380] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c1] =  I0310077d53ae4ed9904df42e3f81c634['h00382] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c2] =  I0310077d53ae4ed9904df42e3f81c634['h00384] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c3] =  I0310077d53ae4ed9904df42e3f81c634['h00386] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c4] =  I0310077d53ae4ed9904df42e3f81c634['h00388] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c5] =  I0310077d53ae4ed9904df42e3f81c634['h0038a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c6] =  I0310077d53ae4ed9904df42e3f81c634['h0038c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c7] =  I0310077d53ae4ed9904df42e3f81c634['h0038e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c8] =  I0310077d53ae4ed9904df42e3f81c634['h00390] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001c9] =  I0310077d53ae4ed9904df42e3f81c634['h00392] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ca] =  I0310077d53ae4ed9904df42e3f81c634['h00394] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001cb] =  I0310077d53ae4ed9904df42e3f81c634['h00396] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001cc] =  I0310077d53ae4ed9904df42e3f81c634['h00398] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001cd] =  I0310077d53ae4ed9904df42e3f81c634['h0039a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ce] =  I0310077d53ae4ed9904df42e3f81c634['h0039c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001cf] =  I0310077d53ae4ed9904df42e3f81c634['h0039e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d0] =  I0310077d53ae4ed9904df42e3f81c634['h003a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d1] =  I0310077d53ae4ed9904df42e3f81c634['h003a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d2] =  I0310077d53ae4ed9904df42e3f81c634['h003a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d3] =  I0310077d53ae4ed9904df42e3f81c634['h003a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d4] =  I0310077d53ae4ed9904df42e3f81c634['h003a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d5] =  I0310077d53ae4ed9904df42e3f81c634['h003aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d6] =  I0310077d53ae4ed9904df42e3f81c634['h003ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d7] =  I0310077d53ae4ed9904df42e3f81c634['h003ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d8] =  I0310077d53ae4ed9904df42e3f81c634['h003b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001d9] =  I0310077d53ae4ed9904df42e3f81c634['h003b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001da] =  I0310077d53ae4ed9904df42e3f81c634['h003b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001db] =  I0310077d53ae4ed9904df42e3f81c634['h003b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001dc] =  I0310077d53ae4ed9904df42e3f81c634['h003b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001dd] =  I0310077d53ae4ed9904df42e3f81c634['h003ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001de] =  I0310077d53ae4ed9904df42e3f81c634['h003bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001df] =  I0310077d53ae4ed9904df42e3f81c634['h003be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e0] =  I0310077d53ae4ed9904df42e3f81c634['h003c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e1] =  I0310077d53ae4ed9904df42e3f81c634['h003c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e2] =  I0310077d53ae4ed9904df42e3f81c634['h003c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e3] =  I0310077d53ae4ed9904df42e3f81c634['h003c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e4] =  I0310077d53ae4ed9904df42e3f81c634['h003c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e5] =  I0310077d53ae4ed9904df42e3f81c634['h003ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e6] =  I0310077d53ae4ed9904df42e3f81c634['h003cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e7] =  I0310077d53ae4ed9904df42e3f81c634['h003ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e8] =  I0310077d53ae4ed9904df42e3f81c634['h003d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001e9] =  I0310077d53ae4ed9904df42e3f81c634['h003d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ea] =  I0310077d53ae4ed9904df42e3f81c634['h003d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001eb] =  I0310077d53ae4ed9904df42e3f81c634['h003d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ec] =  I0310077d53ae4ed9904df42e3f81c634['h003d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ed] =  I0310077d53ae4ed9904df42e3f81c634['h003da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ee] =  I0310077d53ae4ed9904df42e3f81c634['h003dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ef] =  I0310077d53ae4ed9904df42e3f81c634['h003de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f0] =  I0310077d53ae4ed9904df42e3f81c634['h003e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f1] =  I0310077d53ae4ed9904df42e3f81c634['h003e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f2] =  I0310077d53ae4ed9904df42e3f81c634['h003e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f3] =  I0310077d53ae4ed9904df42e3f81c634['h003e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f4] =  I0310077d53ae4ed9904df42e3f81c634['h003e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f5] =  I0310077d53ae4ed9904df42e3f81c634['h003ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f6] =  I0310077d53ae4ed9904df42e3f81c634['h003ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f7] =  I0310077d53ae4ed9904df42e3f81c634['h003ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f8] =  I0310077d53ae4ed9904df42e3f81c634['h003f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001f9] =  I0310077d53ae4ed9904df42e3f81c634['h003f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001fa] =  I0310077d53ae4ed9904df42e3f81c634['h003f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001fb] =  I0310077d53ae4ed9904df42e3f81c634['h003f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001fc] =  I0310077d53ae4ed9904df42e3f81c634['h003f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001fd] =  I0310077d53ae4ed9904df42e3f81c634['h003fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001fe] =  I0310077d53ae4ed9904df42e3f81c634['h003fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h001ff] =  I0310077d53ae4ed9904df42e3f81c634['h003fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00200] =  I0310077d53ae4ed9904df42e3f81c634['h00400] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00201] =  I0310077d53ae4ed9904df42e3f81c634['h00402] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00202] =  I0310077d53ae4ed9904df42e3f81c634['h00404] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00203] =  I0310077d53ae4ed9904df42e3f81c634['h00406] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00204] =  I0310077d53ae4ed9904df42e3f81c634['h00408] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00205] =  I0310077d53ae4ed9904df42e3f81c634['h0040a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00206] =  I0310077d53ae4ed9904df42e3f81c634['h0040c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00207] =  I0310077d53ae4ed9904df42e3f81c634['h0040e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00208] =  I0310077d53ae4ed9904df42e3f81c634['h00410] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00209] =  I0310077d53ae4ed9904df42e3f81c634['h00412] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0020a] =  I0310077d53ae4ed9904df42e3f81c634['h00414] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0020b] =  I0310077d53ae4ed9904df42e3f81c634['h00416] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0020c] =  I0310077d53ae4ed9904df42e3f81c634['h00418] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0020d] =  I0310077d53ae4ed9904df42e3f81c634['h0041a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0020e] =  I0310077d53ae4ed9904df42e3f81c634['h0041c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0020f] =  I0310077d53ae4ed9904df42e3f81c634['h0041e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00210] =  I0310077d53ae4ed9904df42e3f81c634['h00420] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00211] =  I0310077d53ae4ed9904df42e3f81c634['h00422] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00212] =  I0310077d53ae4ed9904df42e3f81c634['h00424] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00213] =  I0310077d53ae4ed9904df42e3f81c634['h00426] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00214] =  I0310077d53ae4ed9904df42e3f81c634['h00428] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00215] =  I0310077d53ae4ed9904df42e3f81c634['h0042a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00216] =  I0310077d53ae4ed9904df42e3f81c634['h0042c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00217] =  I0310077d53ae4ed9904df42e3f81c634['h0042e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00218] =  I0310077d53ae4ed9904df42e3f81c634['h00430] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00219] =  I0310077d53ae4ed9904df42e3f81c634['h00432] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0021a] =  I0310077d53ae4ed9904df42e3f81c634['h00434] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0021b] =  I0310077d53ae4ed9904df42e3f81c634['h00436] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0021c] =  I0310077d53ae4ed9904df42e3f81c634['h00438] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0021d] =  I0310077d53ae4ed9904df42e3f81c634['h0043a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0021e] =  I0310077d53ae4ed9904df42e3f81c634['h0043c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0021f] =  I0310077d53ae4ed9904df42e3f81c634['h0043e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00220] =  I0310077d53ae4ed9904df42e3f81c634['h00440] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00221] =  I0310077d53ae4ed9904df42e3f81c634['h00442] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00222] =  I0310077d53ae4ed9904df42e3f81c634['h00444] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00223] =  I0310077d53ae4ed9904df42e3f81c634['h00446] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00224] =  I0310077d53ae4ed9904df42e3f81c634['h00448] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00225] =  I0310077d53ae4ed9904df42e3f81c634['h0044a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00226] =  I0310077d53ae4ed9904df42e3f81c634['h0044c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00227] =  I0310077d53ae4ed9904df42e3f81c634['h0044e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00228] =  I0310077d53ae4ed9904df42e3f81c634['h00450] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00229] =  I0310077d53ae4ed9904df42e3f81c634['h00452] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0022a] =  I0310077d53ae4ed9904df42e3f81c634['h00454] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0022b] =  I0310077d53ae4ed9904df42e3f81c634['h00456] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0022c] =  I0310077d53ae4ed9904df42e3f81c634['h00458] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0022d] =  I0310077d53ae4ed9904df42e3f81c634['h0045a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0022e] =  I0310077d53ae4ed9904df42e3f81c634['h0045c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0022f] =  I0310077d53ae4ed9904df42e3f81c634['h0045e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00230] =  I0310077d53ae4ed9904df42e3f81c634['h00460] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00231] =  I0310077d53ae4ed9904df42e3f81c634['h00462] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00232] =  I0310077d53ae4ed9904df42e3f81c634['h00464] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00233] =  I0310077d53ae4ed9904df42e3f81c634['h00466] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00234] =  I0310077d53ae4ed9904df42e3f81c634['h00468] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00235] =  I0310077d53ae4ed9904df42e3f81c634['h0046a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00236] =  I0310077d53ae4ed9904df42e3f81c634['h0046c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00237] =  I0310077d53ae4ed9904df42e3f81c634['h0046e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00238] =  I0310077d53ae4ed9904df42e3f81c634['h00470] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00239] =  I0310077d53ae4ed9904df42e3f81c634['h00472] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0023a] =  I0310077d53ae4ed9904df42e3f81c634['h00474] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0023b] =  I0310077d53ae4ed9904df42e3f81c634['h00476] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0023c] =  I0310077d53ae4ed9904df42e3f81c634['h00478] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0023d] =  I0310077d53ae4ed9904df42e3f81c634['h0047a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0023e] =  I0310077d53ae4ed9904df42e3f81c634['h0047c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0023f] =  I0310077d53ae4ed9904df42e3f81c634['h0047e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00240] =  I0310077d53ae4ed9904df42e3f81c634['h00480] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00241] =  I0310077d53ae4ed9904df42e3f81c634['h00482] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00242] =  I0310077d53ae4ed9904df42e3f81c634['h00484] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00243] =  I0310077d53ae4ed9904df42e3f81c634['h00486] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00244] =  I0310077d53ae4ed9904df42e3f81c634['h00488] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00245] =  I0310077d53ae4ed9904df42e3f81c634['h0048a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00246] =  I0310077d53ae4ed9904df42e3f81c634['h0048c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00247] =  I0310077d53ae4ed9904df42e3f81c634['h0048e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00248] =  I0310077d53ae4ed9904df42e3f81c634['h00490] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00249] =  I0310077d53ae4ed9904df42e3f81c634['h00492] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0024a] =  I0310077d53ae4ed9904df42e3f81c634['h00494] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0024b] =  I0310077d53ae4ed9904df42e3f81c634['h00496] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0024c] =  I0310077d53ae4ed9904df42e3f81c634['h00498] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0024d] =  I0310077d53ae4ed9904df42e3f81c634['h0049a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0024e] =  I0310077d53ae4ed9904df42e3f81c634['h0049c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0024f] =  I0310077d53ae4ed9904df42e3f81c634['h0049e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00250] =  I0310077d53ae4ed9904df42e3f81c634['h004a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00251] =  I0310077d53ae4ed9904df42e3f81c634['h004a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00252] =  I0310077d53ae4ed9904df42e3f81c634['h004a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00253] =  I0310077d53ae4ed9904df42e3f81c634['h004a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00254] =  I0310077d53ae4ed9904df42e3f81c634['h004a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00255] =  I0310077d53ae4ed9904df42e3f81c634['h004aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00256] =  I0310077d53ae4ed9904df42e3f81c634['h004ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00257] =  I0310077d53ae4ed9904df42e3f81c634['h004ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00258] =  I0310077d53ae4ed9904df42e3f81c634['h004b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00259] =  I0310077d53ae4ed9904df42e3f81c634['h004b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0025a] =  I0310077d53ae4ed9904df42e3f81c634['h004b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0025b] =  I0310077d53ae4ed9904df42e3f81c634['h004b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0025c] =  I0310077d53ae4ed9904df42e3f81c634['h004b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0025d] =  I0310077d53ae4ed9904df42e3f81c634['h004ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0025e] =  I0310077d53ae4ed9904df42e3f81c634['h004bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0025f] =  I0310077d53ae4ed9904df42e3f81c634['h004be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00260] =  I0310077d53ae4ed9904df42e3f81c634['h004c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00261] =  I0310077d53ae4ed9904df42e3f81c634['h004c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00262] =  I0310077d53ae4ed9904df42e3f81c634['h004c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00263] =  I0310077d53ae4ed9904df42e3f81c634['h004c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00264] =  I0310077d53ae4ed9904df42e3f81c634['h004c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00265] =  I0310077d53ae4ed9904df42e3f81c634['h004ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00266] =  I0310077d53ae4ed9904df42e3f81c634['h004cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00267] =  I0310077d53ae4ed9904df42e3f81c634['h004ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00268] =  I0310077d53ae4ed9904df42e3f81c634['h004d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00269] =  I0310077d53ae4ed9904df42e3f81c634['h004d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0026a] =  I0310077d53ae4ed9904df42e3f81c634['h004d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0026b] =  I0310077d53ae4ed9904df42e3f81c634['h004d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0026c] =  I0310077d53ae4ed9904df42e3f81c634['h004d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0026d] =  I0310077d53ae4ed9904df42e3f81c634['h004da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0026e] =  I0310077d53ae4ed9904df42e3f81c634['h004dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0026f] =  I0310077d53ae4ed9904df42e3f81c634['h004de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00270] =  I0310077d53ae4ed9904df42e3f81c634['h004e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00271] =  I0310077d53ae4ed9904df42e3f81c634['h004e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00272] =  I0310077d53ae4ed9904df42e3f81c634['h004e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00273] =  I0310077d53ae4ed9904df42e3f81c634['h004e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00274] =  I0310077d53ae4ed9904df42e3f81c634['h004e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00275] =  I0310077d53ae4ed9904df42e3f81c634['h004ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00276] =  I0310077d53ae4ed9904df42e3f81c634['h004ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00277] =  I0310077d53ae4ed9904df42e3f81c634['h004ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00278] =  I0310077d53ae4ed9904df42e3f81c634['h004f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00279] =  I0310077d53ae4ed9904df42e3f81c634['h004f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0027a] =  I0310077d53ae4ed9904df42e3f81c634['h004f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0027b] =  I0310077d53ae4ed9904df42e3f81c634['h004f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0027c] =  I0310077d53ae4ed9904df42e3f81c634['h004f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0027d] =  I0310077d53ae4ed9904df42e3f81c634['h004fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0027e] =  I0310077d53ae4ed9904df42e3f81c634['h004fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0027f] =  I0310077d53ae4ed9904df42e3f81c634['h004fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00280] =  I0310077d53ae4ed9904df42e3f81c634['h00500] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00281] =  I0310077d53ae4ed9904df42e3f81c634['h00502] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00282] =  I0310077d53ae4ed9904df42e3f81c634['h00504] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00283] =  I0310077d53ae4ed9904df42e3f81c634['h00506] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00284] =  I0310077d53ae4ed9904df42e3f81c634['h00508] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00285] =  I0310077d53ae4ed9904df42e3f81c634['h0050a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00286] =  I0310077d53ae4ed9904df42e3f81c634['h0050c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00287] =  I0310077d53ae4ed9904df42e3f81c634['h0050e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00288] =  I0310077d53ae4ed9904df42e3f81c634['h00510] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00289] =  I0310077d53ae4ed9904df42e3f81c634['h00512] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0028a] =  I0310077d53ae4ed9904df42e3f81c634['h00514] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0028b] =  I0310077d53ae4ed9904df42e3f81c634['h00516] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0028c] =  I0310077d53ae4ed9904df42e3f81c634['h00518] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0028d] =  I0310077d53ae4ed9904df42e3f81c634['h0051a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0028e] =  I0310077d53ae4ed9904df42e3f81c634['h0051c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0028f] =  I0310077d53ae4ed9904df42e3f81c634['h0051e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00290] =  I0310077d53ae4ed9904df42e3f81c634['h00520] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00291] =  I0310077d53ae4ed9904df42e3f81c634['h00522] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00292] =  I0310077d53ae4ed9904df42e3f81c634['h00524] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00293] =  I0310077d53ae4ed9904df42e3f81c634['h00526] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00294] =  I0310077d53ae4ed9904df42e3f81c634['h00528] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00295] =  I0310077d53ae4ed9904df42e3f81c634['h0052a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00296] =  I0310077d53ae4ed9904df42e3f81c634['h0052c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00297] =  I0310077d53ae4ed9904df42e3f81c634['h0052e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00298] =  I0310077d53ae4ed9904df42e3f81c634['h00530] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00299] =  I0310077d53ae4ed9904df42e3f81c634['h00532] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0029a] =  I0310077d53ae4ed9904df42e3f81c634['h00534] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0029b] =  I0310077d53ae4ed9904df42e3f81c634['h00536] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0029c] =  I0310077d53ae4ed9904df42e3f81c634['h00538] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0029d] =  I0310077d53ae4ed9904df42e3f81c634['h0053a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0029e] =  I0310077d53ae4ed9904df42e3f81c634['h0053c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0029f] =  I0310077d53ae4ed9904df42e3f81c634['h0053e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a0] =  I0310077d53ae4ed9904df42e3f81c634['h00540] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a1] =  I0310077d53ae4ed9904df42e3f81c634['h00542] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a2] =  I0310077d53ae4ed9904df42e3f81c634['h00544] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a3] =  I0310077d53ae4ed9904df42e3f81c634['h00546] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a4] =  I0310077d53ae4ed9904df42e3f81c634['h00548] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a5] =  I0310077d53ae4ed9904df42e3f81c634['h0054a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a6] =  I0310077d53ae4ed9904df42e3f81c634['h0054c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a7] =  I0310077d53ae4ed9904df42e3f81c634['h0054e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a8] =  I0310077d53ae4ed9904df42e3f81c634['h00550] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002a9] =  I0310077d53ae4ed9904df42e3f81c634['h00552] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002aa] =  I0310077d53ae4ed9904df42e3f81c634['h00554] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ab] =  I0310077d53ae4ed9904df42e3f81c634['h00556] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ac] =  I0310077d53ae4ed9904df42e3f81c634['h00558] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ad] =  I0310077d53ae4ed9904df42e3f81c634['h0055a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ae] =  I0310077d53ae4ed9904df42e3f81c634['h0055c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002af] =  I0310077d53ae4ed9904df42e3f81c634['h0055e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b0] =  I0310077d53ae4ed9904df42e3f81c634['h00560] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b1] =  I0310077d53ae4ed9904df42e3f81c634['h00562] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b2] =  I0310077d53ae4ed9904df42e3f81c634['h00564] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b3] =  I0310077d53ae4ed9904df42e3f81c634['h00566] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b4] =  I0310077d53ae4ed9904df42e3f81c634['h00568] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b5] =  I0310077d53ae4ed9904df42e3f81c634['h0056a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b6] =  I0310077d53ae4ed9904df42e3f81c634['h0056c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b7] =  I0310077d53ae4ed9904df42e3f81c634['h0056e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b8] =  I0310077d53ae4ed9904df42e3f81c634['h00570] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002b9] =  I0310077d53ae4ed9904df42e3f81c634['h00572] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ba] =  I0310077d53ae4ed9904df42e3f81c634['h00574] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002bb] =  I0310077d53ae4ed9904df42e3f81c634['h00576] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002bc] =  I0310077d53ae4ed9904df42e3f81c634['h00578] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002bd] =  I0310077d53ae4ed9904df42e3f81c634['h0057a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002be] =  I0310077d53ae4ed9904df42e3f81c634['h0057c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002bf] =  I0310077d53ae4ed9904df42e3f81c634['h0057e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c0] =  I0310077d53ae4ed9904df42e3f81c634['h00580] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c1] =  I0310077d53ae4ed9904df42e3f81c634['h00582] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c2] =  I0310077d53ae4ed9904df42e3f81c634['h00584] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c3] =  I0310077d53ae4ed9904df42e3f81c634['h00586] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c4] =  I0310077d53ae4ed9904df42e3f81c634['h00588] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c5] =  I0310077d53ae4ed9904df42e3f81c634['h0058a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c6] =  I0310077d53ae4ed9904df42e3f81c634['h0058c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c7] =  I0310077d53ae4ed9904df42e3f81c634['h0058e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c8] =  I0310077d53ae4ed9904df42e3f81c634['h00590] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002c9] =  I0310077d53ae4ed9904df42e3f81c634['h00592] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ca] =  I0310077d53ae4ed9904df42e3f81c634['h00594] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002cb] =  I0310077d53ae4ed9904df42e3f81c634['h00596] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002cc] =  I0310077d53ae4ed9904df42e3f81c634['h00598] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002cd] =  I0310077d53ae4ed9904df42e3f81c634['h0059a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ce] =  I0310077d53ae4ed9904df42e3f81c634['h0059c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002cf] =  I0310077d53ae4ed9904df42e3f81c634['h0059e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d0] =  I0310077d53ae4ed9904df42e3f81c634['h005a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d1] =  I0310077d53ae4ed9904df42e3f81c634['h005a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d2] =  I0310077d53ae4ed9904df42e3f81c634['h005a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d3] =  I0310077d53ae4ed9904df42e3f81c634['h005a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d4] =  I0310077d53ae4ed9904df42e3f81c634['h005a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d5] =  I0310077d53ae4ed9904df42e3f81c634['h005aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d6] =  I0310077d53ae4ed9904df42e3f81c634['h005ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d7] =  I0310077d53ae4ed9904df42e3f81c634['h005ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d8] =  I0310077d53ae4ed9904df42e3f81c634['h005b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002d9] =  I0310077d53ae4ed9904df42e3f81c634['h005b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002da] =  I0310077d53ae4ed9904df42e3f81c634['h005b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002db] =  I0310077d53ae4ed9904df42e3f81c634['h005b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002dc] =  I0310077d53ae4ed9904df42e3f81c634['h005b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002dd] =  I0310077d53ae4ed9904df42e3f81c634['h005ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002de] =  I0310077d53ae4ed9904df42e3f81c634['h005bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002df] =  I0310077d53ae4ed9904df42e3f81c634['h005be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e0] =  I0310077d53ae4ed9904df42e3f81c634['h005c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e1] =  I0310077d53ae4ed9904df42e3f81c634['h005c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e2] =  I0310077d53ae4ed9904df42e3f81c634['h005c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e3] =  I0310077d53ae4ed9904df42e3f81c634['h005c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e4] =  I0310077d53ae4ed9904df42e3f81c634['h005c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e5] =  I0310077d53ae4ed9904df42e3f81c634['h005ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e6] =  I0310077d53ae4ed9904df42e3f81c634['h005cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e7] =  I0310077d53ae4ed9904df42e3f81c634['h005ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e8] =  I0310077d53ae4ed9904df42e3f81c634['h005d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002e9] =  I0310077d53ae4ed9904df42e3f81c634['h005d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ea] =  I0310077d53ae4ed9904df42e3f81c634['h005d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002eb] =  I0310077d53ae4ed9904df42e3f81c634['h005d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ec] =  I0310077d53ae4ed9904df42e3f81c634['h005d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ed] =  I0310077d53ae4ed9904df42e3f81c634['h005da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ee] =  I0310077d53ae4ed9904df42e3f81c634['h005dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ef] =  I0310077d53ae4ed9904df42e3f81c634['h005de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f0] =  I0310077d53ae4ed9904df42e3f81c634['h005e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f1] =  I0310077d53ae4ed9904df42e3f81c634['h005e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f2] =  I0310077d53ae4ed9904df42e3f81c634['h005e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f3] =  I0310077d53ae4ed9904df42e3f81c634['h005e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f4] =  I0310077d53ae4ed9904df42e3f81c634['h005e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f5] =  I0310077d53ae4ed9904df42e3f81c634['h005ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f6] =  I0310077d53ae4ed9904df42e3f81c634['h005ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f7] =  I0310077d53ae4ed9904df42e3f81c634['h005ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f8] =  I0310077d53ae4ed9904df42e3f81c634['h005f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002f9] =  I0310077d53ae4ed9904df42e3f81c634['h005f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002fa] =  I0310077d53ae4ed9904df42e3f81c634['h005f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002fb] =  I0310077d53ae4ed9904df42e3f81c634['h005f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002fc] =  I0310077d53ae4ed9904df42e3f81c634['h005f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002fd] =  I0310077d53ae4ed9904df42e3f81c634['h005fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002fe] =  I0310077d53ae4ed9904df42e3f81c634['h005fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h002ff] =  I0310077d53ae4ed9904df42e3f81c634['h005fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00300] =  I0310077d53ae4ed9904df42e3f81c634['h00600] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00301] =  I0310077d53ae4ed9904df42e3f81c634['h00602] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00302] =  I0310077d53ae4ed9904df42e3f81c634['h00604] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00303] =  I0310077d53ae4ed9904df42e3f81c634['h00606] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00304] =  I0310077d53ae4ed9904df42e3f81c634['h00608] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00305] =  I0310077d53ae4ed9904df42e3f81c634['h0060a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00306] =  I0310077d53ae4ed9904df42e3f81c634['h0060c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00307] =  I0310077d53ae4ed9904df42e3f81c634['h0060e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00308] =  I0310077d53ae4ed9904df42e3f81c634['h00610] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00309] =  I0310077d53ae4ed9904df42e3f81c634['h00612] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0030a] =  I0310077d53ae4ed9904df42e3f81c634['h00614] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0030b] =  I0310077d53ae4ed9904df42e3f81c634['h00616] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0030c] =  I0310077d53ae4ed9904df42e3f81c634['h00618] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0030d] =  I0310077d53ae4ed9904df42e3f81c634['h0061a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0030e] =  I0310077d53ae4ed9904df42e3f81c634['h0061c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0030f] =  I0310077d53ae4ed9904df42e3f81c634['h0061e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00310] =  I0310077d53ae4ed9904df42e3f81c634['h00620] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00311] =  I0310077d53ae4ed9904df42e3f81c634['h00622] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00312] =  I0310077d53ae4ed9904df42e3f81c634['h00624] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00313] =  I0310077d53ae4ed9904df42e3f81c634['h00626] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00314] =  I0310077d53ae4ed9904df42e3f81c634['h00628] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00315] =  I0310077d53ae4ed9904df42e3f81c634['h0062a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00316] =  I0310077d53ae4ed9904df42e3f81c634['h0062c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00317] =  I0310077d53ae4ed9904df42e3f81c634['h0062e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00318] =  I0310077d53ae4ed9904df42e3f81c634['h00630] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00319] =  I0310077d53ae4ed9904df42e3f81c634['h00632] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0031a] =  I0310077d53ae4ed9904df42e3f81c634['h00634] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0031b] =  I0310077d53ae4ed9904df42e3f81c634['h00636] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0031c] =  I0310077d53ae4ed9904df42e3f81c634['h00638] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0031d] =  I0310077d53ae4ed9904df42e3f81c634['h0063a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0031e] =  I0310077d53ae4ed9904df42e3f81c634['h0063c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0031f] =  I0310077d53ae4ed9904df42e3f81c634['h0063e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00320] =  I0310077d53ae4ed9904df42e3f81c634['h00640] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00321] =  I0310077d53ae4ed9904df42e3f81c634['h00642] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00322] =  I0310077d53ae4ed9904df42e3f81c634['h00644] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00323] =  I0310077d53ae4ed9904df42e3f81c634['h00646] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00324] =  I0310077d53ae4ed9904df42e3f81c634['h00648] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00325] =  I0310077d53ae4ed9904df42e3f81c634['h0064a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00326] =  I0310077d53ae4ed9904df42e3f81c634['h0064c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00327] =  I0310077d53ae4ed9904df42e3f81c634['h0064e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00328] =  I0310077d53ae4ed9904df42e3f81c634['h00650] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00329] =  I0310077d53ae4ed9904df42e3f81c634['h00652] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0032a] =  I0310077d53ae4ed9904df42e3f81c634['h00654] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0032b] =  I0310077d53ae4ed9904df42e3f81c634['h00656] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0032c] =  I0310077d53ae4ed9904df42e3f81c634['h00658] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0032d] =  I0310077d53ae4ed9904df42e3f81c634['h0065a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0032e] =  I0310077d53ae4ed9904df42e3f81c634['h0065c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0032f] =  I0310077d53ae4ed9904df42e3f81c634['h0065e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00330] =  I0310077d53ae4ed9904df42e3f81c634['h00660] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00331] =  I0310077d53ae4ed9904df42e3f81c634['h00662] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00332] =  I0310077d53ae4ed9904df42e3f81c634['h00664] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00333] =  I0310077d53ae4ed9904df42e3f81c634['h00666] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00334] =  I0310077d53ae4ed9904df42e3f81c634['h00668] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00335] =  I0310077d53ae4ed9904df42e3f81c634['h0066a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00336] =  I0310077d53ae4ed9904df42e3f81c634['h0066c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00337] =  I0310077d53ae4ed9904df42e3f81c634['h0066e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00338] =  I0310077d53ae4ed9904df42e3f81c634['h00670] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00339] =  I0310077d53ae4ed9904df42e3f81c634['h00672] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0033a] =  I0310077d53ae4ed9904df42e3f81c634['h00674] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0033b] =  I0310077d53ae4ed9904df42e3f81c634['h00676] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0033c] =  I0310077d53ae4ed9904df42e3f81c634['h00678] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0033d] =  I0310077d53ae4ed9904df42e3f81c634['h0067a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0033e] =  I0310077d53ae4ed9904df42e3f81c634['h0067c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0033f] =  I0310077d53ae4ed9904df42e3f81c634['h0067e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00340] =  I0310077d53ae4ed9904df42e3f81c634['h00680] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00341] =  I0310077d53ae4ed9904df42e3f81c634['h00682] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00342] =  I0310077d53ae4ed9904df42e3f81c634['h00684] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00343] =  I0310077d53ae4ed9904df42e3f81c634['h00686] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00344] =  I0310077d53ae4ed9904df42e3f81c634['h00688] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00345] =  I0310077d53ae4ed9904df42e3f81c634['h0068a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00346] =  I0310077d53ae4ed9904df42e3f81c634['h0068c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00347] =  I0310077d53ae4ed9904df42e3f81c634['h0068e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00348] =  I0310077d53ae4ed9904df42e3f81c634['h00690] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00349] =  I0310077d53ae4ed9904df42e3f81c634['h00692] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0034a] =  I0310077d53ae4ed9904df42e3f81c634['h00694] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0034b] =  I0310077d53ae4ed9904df42e3f81c634['h00696] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0034c] =  I0310077d53ae4ed9904df42e3f81c634['h00698] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0034d] =  I0310077d53ae4ed9904df42e3f81c634['h0069a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0034e] =  I0310077d53ae4ed9904df42e3f81c634['h0069c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0034f] =  I0310077d53ae4ed9904df42e3f81c634['h0069e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00350] =  I0310077d53ae4ed9904df42e3f81c634['h006a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00351] =  I0310077d53ae4ed9904df42e3f81c634['h006a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00352] =  I0310077d53ae4ed9904df42e3f81c634['h006a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00353] =  I0310077d53ae4ed9904df42e3f81c634['h006a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00354] =  I0310077d53ae4ed9904df42e3f81c634['h006a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00355] =  I0310077d53ae4ed9904df42e3f81c634['h006aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00356] =  I0310077d53ae4ed9904df42e3f81c634['h006ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00357] =  I0310077d53ae4ed9904df42e3f81c634['h006ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00358] =  I0310077d53ae4ed9904df42e3f81c634['h006b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00359] =  I0310077d53ae4ed9904df42e3f81c634['h006b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0035a] =  I0310077d53ae4ed9904df42e3f81c634['h006b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0035b] =  I0310077d53ae4ed9904df42e3f81c634['h006b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0035c] =  I0310077d53ae4ed9904df42e3f81c634['h006b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0035d] =  I0310077d53ae4ed9904df42e3f81c634['h006ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0035e] =  I0310077d53ae4ed9904df42e3f81c634['h006bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0035f] =  I0310077d53ae4ed9904df42e3f81c634['h006be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00360] =  I0310077d53ae4ed9904df42e3f81c634['h006c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00361] =  I0310077d53ae4ed9904df42e3f81c634['h006c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00362] =  I0310077d53ae4ed9904df42e3f81c634['h006c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00363] =  I0310077d53ae4ed9904df42e3f81c634['h006c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00364] =  I0310077d53ae4ed9904df42e3f81c634['h006c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00365] =  I0310077d53ae4ed9904df42e3f81c634['h006ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00366] =  I0310077d53ae4ed9904df42e3f81c634['h006cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00367] =  I0310077d53ae4ed9904df42e3f81c634['h006ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00368] =  I0310077d53ae4ed9904df42e3f81c634['h006d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00369] =  I0310077d53ae4ed9904df42e3f81c634['h006d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0036a] =  I0310077d53ae4ed9904df42e3f81c634['h006d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0036b] =  I0310077d53ae4ed9904df42e3f81c634['h006d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0036c] =  I0310077d53ae4ed9904df42e3f81c634['h006d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0036d] =  I0310077d53ae4ed9904df42e3f81c634['h006da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0036e] =  I0310077d53ae4ed9904df42e3f81c634['h006dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0036f] =  I0310077d53ae4ed9904df42e3f81c634['h006de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00370] =  I0310077d53ae4ed9904df42e3f81c634['h006e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00371] =  I0310077d53ae4ed9904df42e3f81c634['h006e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00372] =  I0310077d53ae4ed9904df42e3f81c634['h006e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00373] =  I0310077d53ae4ed9904df42e3f81c634['h006e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00374] =  I0310077d53ae4ed9904df42e3f81c634['h006e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00375] =  I0310077d53ae4ed9904df42e3f81c634['h006ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00376] =  I0310077d53ae4ed9904df42e3f81c634['h006ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00377] =  I0310077d53ae4ed9904df42e3f81c634['h006ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00378] =  I0310077d53ae4ed9904df42e3f81c634['h006f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00379] =  I0310077d53ae4ed9904df42e3f81c634['h006f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0037a] =  I0310077d53ae4ed9904df42e3f81c634['h006f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0037b] =  I0310077d53ae4ed9904df42e3f81c634['h006f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0037c] =  I0310077d53ae4ed9904df42e3f81c634['h006f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0037d] =  I0310077d53ae4ed9904df42e3f81c634['h006fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0037e] =  I0310077d53ae4ed9904df42e3f81c634['h006fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0037f] =  I0310077d53ae4ed9904df42e3f81c634['h006fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00380] =  I0310077d53ae4ed9904df42e3f81c634['h00700] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00381] =  I0310077d53ae4ed9904df42e3f81c634['h00702] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00382] =  I0310077d53ae4ed9904df42e3f81c634['h00704] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00383] =  I0310077d53ae4ed9904df42e3f81c634['h00706] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00384] =  I0310077d53ae4ed9904df42e3f81c634['h00708] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00385] =  I0310077d53ae4ed9904df42e3f81c634['h0070a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00386] =  I0310077d53ae4ed9904df42e3f81c634['h0070c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00387] =  I0310077d53ae4ed9904df42e3f81c634['h0070e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00388] =  I0310077d53ae4ed9904df42e3f81c634['h00710] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00389] =  I0310077d53ae4ed9904df42e3f81c634['h00712] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0038a] =  I0310077d53ae4ed9904df42e3f81c634['h00714] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0038b] =  I0310077d53ae4ed9904df42e3f81c634['h00716] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0038c] =  I0310077d53ae4ed9904df42e3f81c634['h00718] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0038d] =  I0310077d53ae4ed9904df42e3f81c634['h0071a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0038e] =  I0310077d53ae4ed9904df42e3f81c634['h0071c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0038f] =  I0310077d53ae4ed9904df42e3f81c634['h0071e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00390] =  I0310077d53ae4ed9904df42e3f81c634['h00720] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00391] =  I0310077d53ae4ed9904df42e3f81c634['h00722] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00392] =  I0310077d53ae4ed9904df42e3f81c634['h00724] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00393] =  I0310077d53ae4ed9904df42e3f81c634['h00726] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00394] =  I0310077d53ae4ed9904df42e3f81c634['h00728] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00395] =  I0310077d53ae4ed9904df42e3f81c634['h0072a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00396] =  I0310077d53ae4ed9904df42e3f81c634['h0072c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00397] =  I0310077d53ae4ed9904df42e3f81c634['h0072e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00398] =  I0310077d53ae4ed9904df42e3f81c634['h00730] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00399] =  I0310077d53ae4ed9904df42e3f81c634['h00732] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0039a] =  I0310077d53ae4ed9904df42e3f81c634['h00734] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0039b] =  I0310077d53ae4ed9904df42e3f81c634['h00736] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0039c] =  I0310077d53ae4ed9904df42e3f81c634['h00738] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0039d] =  I0310077d53ae4ed9904df42e3f81c634['h0073a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0039e] =  I0310077d53ae4ed9904df42e3f81c634['h0073c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0039f] =  I0310077d53ae4ed9904df42e3f81c634['h0073e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a0] =  I0310077d53ae4ed9904df42e3f81c634['h00740] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a1] =  I0310077d53ae4ed9904df42e3f81c634['h00742] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a2] =  I0310077d53ae4ed9904df42e3f81c634['h00744] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a3] =  I0310077d53ae4ed9904df42e3f81c634['h00746] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a4] =  I0310077d53ae4ed9904df42e3f81c634['h00748] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a5] =  I0310077d53ae4ed9904df42e3f81c634['h0074a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a6] =  I0310077d53ae4ed9904df42e3f81c634['h0074c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a7] =  I0310077d53ae4ed9904df42e3f81c634['h0074e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a8] =  I0310077d53ae4ed9904df42e3f81c634['h00750] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003a9] =  I0310077d53ae4ed9904df42e3f81c634['h00752] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003aa] =  I0310077d53ae4ed9904df42e3f81c634['h00754] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ab] =  I0310077d53ae4ed9904df42e3f81c634['h00756] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ac] =  I0310077d53ae4ed9904df42e3f81c634['h00758] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ad] =  I0310077d53ae4ed9904df42e3f81c634['h0075a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ae] =  I0310077d53ae4ed9904df42e3f81c634['h0075c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003af] =  I0310077d53ae4ed9904df42e3f81c634['h0075e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b0] =  I0310077d53ae4ed9904df42e3f81c634['h00760] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b1] =  I0310077d53ae4ed9904df42e3f81c634['h00762] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b2] =  I0310077d53ae4ed9904df42e3f81c634['h00764] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b3] =  I0310077d53ae4ed9904df42e3f81c634['h00766] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b4] =  I0310077d53ae4ed9904df42e3f81c634['h00768] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b5] =  I0310077d53ae4ed9904df42e3f81c634['h0076a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b6] =  I0310077d53ae4ed9904df42e3f81c634['h0076c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b7] =  I0310077d53ae4ed9904df42e3f81c634['h0076e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b8] =  I0310077d53ae4ed9904df42e3f81c634['h00770] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003b9] =  I0310077d53ae4ed9904df42e3f81c634['h00772] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ba] =  I0310077d53ae4ed9904df42e3f81c634['h00774] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003bb] =  I0310077d53ae4ed9904df42e3f81c634['h00776] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003bc] =  I0310077d53ae4ed9904df42e3f81c634['h00778] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003bd] =  I0310077d53ae4ed9904df42e3f81c634['h0077a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003be] =  I0310077d53ae4ed9904df42e3f81c634['h0077c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003bf] =  I0310077d53ae4ed9904df42e3f81c634['h0077e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c0] =  I0310077d53ae4ed9904df42e3f81c634['h00780] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c1] =  I0310077d53ae4ed9904df42e3f81c634['h00782] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c2] =  I0310077d53ae4ed9904df42e3f81c634['h00784] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c3] =  I0310077d53ae4ed9904df42e3f81c634['h00786] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c4] =  I0310077d53ae4ed9904df42e3f81c634['h00788] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c5] =  I0310077d53ae4ed9904df42e3f81c634['h0078a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c6] =  I0310077d53ae4ed9904df42e3f81c634['h0078c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c7] =  I0310077d53ae4ed9904df42e3f81c634['h0078e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c8] =  I0310077d53ae4ed9904df42e3f81c634['h00790] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003c9] =  I0310077d53ae4ed9904df42e3f81c634['h00792] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ca] =  I0310077d53ae4ed9904df42e3f81c634['h00794] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003cb] =  I0310077d53ae4ed9904df42e3f81c634['h00796] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003cc] =  I0310077d53ae4ed9904df42e3f81c634['h00798] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003cd] =  I0310077d53ae4ed9904df42e3f81c634['h0079a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ce] =  I0310077d53ae4ed9904df42e3f81c634['h0079c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003cf] =  I0310077d53ae4ed9904df42e3f81c634['h0079e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d0] =  I0310077d53ae4ed9904df42e3f81c634['h007a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d1] =  I0310077d53ae4ed9904df42e3f81c634['h007a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d2] =  I0310077d53ae4ed9904df42e3f81c634['h007a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d3] =  I0310077d53ae4ed9904df42e3f81c634['h007a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d4] =  I0310077d53ae4ed9904df42e3f81c634['h007a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d5] =  I0310077d53ae4ed9904df42e3f81c634['h007aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d6] =  I0310077d53ae4ed9904df42e3f81c634['h007ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d7] =  I0310077d53ae4ed9904df42e3f81c634['h007ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d8] =  I0310077d53ae4ed9904df42e3f81c634['h007b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003d9] =  I0310077d53ae4ed9904df42e3f81c634['h007b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003da] =  I0310077d53ae4ed9904df42e3f81c634['h007b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003db] =  I0310077d53ae4ed9904df42e3f81c634['h007b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003dc] =  I0310077d53ae4ed9904df42e3f81c634['h007b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003dd] =  I0310077d53ae4ed9904df42e3f81c634['h007ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003de] =  I0310077d53ae4ed9904df42e3f81c634['h007bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003df] =  I0310077d53ae4ed9904df42e3f81c634['h007be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e0] =  I0310077d53ae4ed9904df42e3f81c634['h007c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e1] =  I0310077d53ae4ed9904df42e3f81c634['h007c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e2] =  I0310077d53ae4ed9904df42e3f81c634['h007c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e3] =  I0310077d53ae4ed9904df42e3f81c634['h007c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e4] =  I0310077d53ae4ed9904df42e3f81c634['h007c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e5] =  I0310077d53ae4ed9904df42e3f81c634['h007ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e6] =  I0310077d53ae4ed9904df42e3f81c634['h007cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e7] =  I0310077d53ae4ed9904df42e3f81c634['h007ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e8] =  I0310077d53ae4ed9904df42e3f81c634['h007d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003e9] =  I0310077d53ae4ed9904df42e3f81c634['h007d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ea] =  I0310077d53ae4ed9904df42e3f81c634['h007d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003eb] =  I0310077d53ae4ed9904df42e3f81c634['h007d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ec] =  I0310077d53ae4ed9904df42e3f81c634['h007d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ed] =  I0310077d53ae4ed9904df42e3f81c634['h007da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ee] =  I0310077d53ae4ed9904df42e3f81c634['h007dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ef] =  I0310077d53ae4ed9904df42e3f81c634['h007de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f0] =  I0310077d53ae4ed9904df42e3f81c634['h007e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f1] =  I0310077d53ae4ed9904df42e3f81c634['h007e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f2] =  I0310077d53ae4ed9904df42e3f81c634['h007e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f3] =  I0310077d53ae4ed9904df42e3f81c634['h007e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f4] =  I0310077d53ae4ed9904df42e3f81c634['h007e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f5] =  I0310077d53ae4ed9904df42e3f81c634['h007ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f6] =  I0310077d53ae4ed9904df42e3f81c634['h007ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f7] =  I0310077d53ae4ed9904df42e3f81c634['h007ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f8] =  I0310077d53ae4ed9904df42e3f81c634['h007f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003f9] =  I0310077d53ae4ed9904df42e3f81c634['h007f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003fa] =  I0310077d53ae4ed9904df42e3f81c634['h007f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003fb] =  I0310077d53ae4ed9904df42e3f81c634['h007f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003fc] =  I0310077d53ae4ed9904df42e3f81c634['h007f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003fd] =  I0310077d53ae4ed9904df42e3f81c634['h007fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003fe] =  I0310077d53ae4ed9904df42e3f81c634['h007fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h003ff] =  I0310077d53ae4ed9904df42e3f81c634['h007fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00400] =  I0310077d53ae4ed9904df42e3f81c634['h00800] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00401] =  I0310077d53ae4ed9904df42e3f81c634['h00802] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00402] =  I0310077d53ae4ed9904df42e3f81c634['h00804] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00403] =  I0310077d53ae4ed9904df42e3f81c634['h00806] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00404] =  I0310077d53ae4ed9904df42e3f81c634['h00808] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00405] =  I0310077d53ae4ed9904df42e3f81c634['h0080a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00406] =  I0310077d53ae4ed9904df42e3f81c634['h0080c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00407] =  I0310077d53ae4ed9904df42e3f81c634['h0080e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00408] =  I0310077d53ae4ed9904df42e3f81c634['h00810] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00409] =  I0310077d53ae4ed9904df42e3f81c634['h00812] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0040a] =  I0310077d53ae4ed9904df42e3f81c634['h00814] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0040b] =  I0310077d53ae4ed9904df42e3f81c634['h00816] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0040c] =  I0310077d53ae4ed9904df42e3f81c634['h00818] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0040d] =  I0310077d53ae4ed9904df42e3f81c634['h0081a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0040e] =  I0310077d53ae4ed9904df42e3f81c634['h0081c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0040f] =  I0310077d53ae4ed9904df42e3f81c634['h0081e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00410] =  I0310077d53ae4ed9904df42e3f81c634['h00820] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00411] =  I0310077d53ae4ed9904df42e3f81c634['h00822] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00412] =  I0310077d53ae4ed9904df42e3f81c634['h00824] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00413] =  I0310077d53ae4ed9904df42e3f81c634['h00826] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00414] =  I0310077d53ae4ed9904df42e3f81c634['h00828] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00415] =  I0310077d53ae4ed9904df42e3f81c634['h0082a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00416] =  I0310077d53ae4ed9904df42e3f81c634['h0082c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00417] =  I0310077d53ae4ed9904df42e3f81c634['h0082e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00418] =  I0310077d53ae4ed9904df42e3f81c634['h00830] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00419] =  I0310077d53ae4ed9904df42e3f81c634['h00832] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0041a] =  I0310077d53ae4ed9904df42e3f81c634['h00834] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0041b] =  I0310077d53ae4ed9904df42e3f81c634['h00836] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0041c] =  I0310077d53ae4ed9904df42e3f81c634['h00838] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0041d] =  I0310077d53ae4ed9904df42e3f81c634['h0083a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0041e] =  I0310077d53ae4ed9904df42e3f81c634['h0083c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0041f] =  I0310077d53ae4ed9904df42e3f81c634['h0083e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00420] =  I0310077d53ae4ed9904df42e3f81c634['h00840] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00421] =  I0310077d53ae4ed9904df42e3f81c634['h00842] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00422] =  I0310077d53ae4ed9904df42e3f81c634['h00844] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00423] =  I0310077d53ae4ed9904df42e3f81c634['h00846] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00424] =  I0310077d53ae4ed9904df42e3f81c634['h00848] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00425] =  I0310077d53ae4ed9904df42e3f81c634['h0084a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00426] =  I0310077d53ae4ed9904df42e3f81c634['h0084c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00427] =  I0310077d53ae4ed9904df42e3f81c634['h0084e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00428] =  I0310077d53ae4ed9904df42e3f81c634['h00850] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00429] =  I0310077d53ae4ed9904df42e3f81c634['h00852] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0042a] =  I0310077d53ae4ed9904df42e3f81c634['h00854] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0042b] =  I0310077d53ae4ed9904df42e3f81c634['h00856] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0042c] =  I0310077d53ae4ed9904df42e3f81c634['h00858] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0042d] =  I0310077d53ae4ed9904df42e3f81c634['h0085a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0042e] =  I0310077d53ae4ed9904df42e3f81c634['h0085c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0042f] =  I0310077d53ae4ed9904df42e3f81c634['h0085e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00430] =  I0310077d53ae4ed9904df42e3f81c634['h00860] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00431] =  I0310077d53ae4ed9904df42e3f81c634['h00862] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00432] =  I0310077d53ae4ed9904df42e3f81c634['h00864] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00433] =  I0310077d53ae4ed9904df42e3f81c634['h00866] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00434] =  I0310077d53ae4ed9904df42e3f81c634['h00868] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00435] =  I0310077d53ae4ed9904df42e3f81c634['h0086a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00436] =  I0310077d53ae4ed9904df42e3f81c634['h0086c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00437] =  I0310077d53ae4ed9904df42e3f81c634['h0086e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00438] =  I0310077d53ae4ed9904df42e3f81c634['h00870] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00439] =  I0310077d53ae4ed9904df42e3f81c634['h00872] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0043a] =  I0310077d53ae4ed9904df42e3f81c634['h00874] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0043b] =  I0310077d53ae4ed9904df42e3f81c634['h00876] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0043c] =  I0310077d53ae4ed9904df42e3f81c634['h00878] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0043d] =  I0310077d53ae4ed9904df42e3f81c634['h0087a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0043e] =  I0310077d53ae4ed9904df42e3f81c634['h0087c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0043f] =  I0310077d53ae4ed9904df42e3f81c634['h0087e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00440] =  I0310077d53ae4ed9904df42e3f81c634['h00880] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00441] =  I0310077d53ae4ed9904df42e3f81c634['h00882] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00442] =  I0310077d53ae4ed9904df42e3f81c634['h00884] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00443] =  I0310077d53ae4ed9904df42e3f81c634['h00886] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00444] =  I0310077d53ae4ed9904df42e3f81c634['h00888] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00445] =  I0310077d53ae4ed9904df42e3f81c634['h0088a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00446] =  I0310077d53ae4ed9904df42e3f81c634['h0088c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00447] =  I0310077d53ae4ed9904df42e3f81c634['h0088e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00448] =  I0310077d53ae4ed9904df42e3f81c634['h00890] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00449] =  I0310077d53ae4ed9904df42e3f81c634['h00892] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0044a] =  I0310077d53ae4ed9904df42e3f81c634['h00894] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0044b] =  I0310077d53ae4ed9904df42e3f81c634['h00896] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0044c] =  I0310077d53ae4ed9904df42e3f81c634['h00898] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0044d] =  I0310077d53ae4ed9904df42e3f81c634['h0089a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0044e] =  I0310077d53ae4ed9904df42e3f81c634['h0089c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0044f] =  I0310077d53ae4ed9904df42e3f81c634['h0089e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00450] =  I0310077d53ae4ed9904df42e3f81c634['h008a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00451] =  I0310077d53ae4ed9904df42e3f81c634['h008a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00452] =  I0310077d53ae4ed9904df42e3f81c634['h008a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00453] =  I0310077d53ae4ed9904df42e3f81c634['h008a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00454] =  I0310077d53ae4ed9904df42e3f81c634['h008a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00455] =  I0310077d53ae4ed9904df42e3f81c634['h008aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00456] =  I0310077d53ae4ed9904df42e3f81c634['h008ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00457] =  I0310077d53ae4ed9904df42e3f81c634['h008ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00458] =  I0310077d53ae4ed9904df42e3f81c634['h008b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00459] =  I0310077d53ae4ed9904df42e3f81c634['h008b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0045a] =  I0310077d53ae4ed9904df42e3f81c634['h008b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0045b] =  I0310077d53ae4ed9904df42e3f81c634['h008b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0045c] =  I0310077d53ae4ed9904df42e3f81c634['h008b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0045d] =  I0310077d53ae4ed9904df42e3f81c634['h008ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0045e] =  I0310077d53ae4ed9904df42e3f81c634['h008bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0045f] =  I0310077d53ae4ed9904df42e3f81c634['h008be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00460] =  I0310077d53ae4ed9904df42e3f81c634['h008c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00461] =  I0310077d53ae4ed9904df42e3f81c634['h008c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00462] =  I0310077d53ae4ed9904df42e3f81c634['h008c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00463] =  I0310077d53ae4ed9904df42e3f81c634['h008c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00464] =  I0310077d53ae4ed9904df42e3f81c634['h008c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00465] =  I0310077d53ae4ed9904df42e3f81c634['h008ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00466] =  I0310077d53ae4ed9904df42e3f81c634['h008cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00467] =  I0310077d53ae4ed9904df42e3f81c634['h008ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00468] =  I0310077d53ae4ed9904df42e3f81c634['h008d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00469] =  I0310077d53ae4ed9904df42e3f81c634['h008d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0046a] =  I0310077d53ae4ed9904df42e3f81c634['h008d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0046b] =  I0310077d53ae4ed9904df42e3f81c634['h008d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0046c] =  I0310077d53ae4ed9904df42e3f81c634['h008d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0046d] =  I0310077d53ae4ed9904df42e3f81c634['h008da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0046e] =  I0310077d53ae4ed9904df42e3f81c634['h008dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0046f] =  I0310077d53ae4ed9904df42e3f81c634['h008de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00470] =  I0310077d53ae4ed9904df42e3f81c634['h008e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00471] =  I0310077d53ae4ed9904df42e3f81c634['h008e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00472] =  I0310077d53ae4ed9904df42e3f81c634['h008e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00473] =  I0310077d53ae4ed9904df42e3f81c634['h008e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00474] =  I0310077d53ae4ed9904df42e3f81c634['h008e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00475] =  I0310077d53ae4ed9904df42e3f81c634['h008ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00476] =  I0310077d53ae4ed9904df42e3f81c634['h008ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00477] =  I0310077d53ae4ed9904df42e3f81c634['h008ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00478] =  I0310077d53ae4ed9904df42e3f81c634['h008f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00479] =  I0310077d53ae4ed9904df42e3f81c634['h008f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0047a] =  I0310077d53ae4ed9904df42e3f81c634['h008f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0047b] =  I0310077d53ae4ed9904df42e3f81c634['h008f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0047c] =  I0310077d53ae4ed9904df42e3f81c634['h008f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0047d] =  I0310077d53ae4ed9904df42e3f81c634['h008fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0047e] =  I0310077d53ae4ed9904df42e3f81c634['h008fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0047f] =  I0310077d53ae4ed9904df42e3f81c634['h008fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00480] =  I0310077d53ae4ed9904df42e3f81c634['h00900] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00481] =  I0310077d53ae4ed9904df42e3f81c634['h00902] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00482] =  I0310077d53ae4ed9904df42e3f81c634['h00904] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00483] =  I0310077d53ae4ed9904df42e3f81c634['h00906] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00484] =  I0310077d53ae4ed9904df42e3f81c634['h00908] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00485] =  I0310077d53ae4ed9904df42e3f81c634['h0090a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00486] =  I0310077d53ae4ed9904df42e3f81c634['h0090c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00487] =  I0310077d53ae4ed9904df42e3f81c634['h0090e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00488] =  I0310077d53ae4ed9904df42e3f81c634['h00910] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00489] =  I0310077d53ae4ed9904df42e3f81c634['h00912] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0048a] =  I0310077d53ae4ed9904df42e3f81c634['h00914] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0048b] =  I0310077d53ae4ed9904df42e3f81c634['h00916] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0048c] =  I0310077d53ae4ed9904df42e3f81c634['h00918] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0048d] =  I0310077d53ae4ed9904df42e3f81c634['h0091a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0048e] =  I0310077d53ae4ed9904df42e3f81c634['h0091c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0048f] =  I0310077d53ae4ed9904df42e3f81c634['h0091e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00490] =  I0310077d53ae4ed9904df42e3f81c634['h00920] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00491] =  I0310077d53ae4ed9904df42e3f81c634['h00922] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00492] =  I0310077d53ae4ed9904df42e3f81c634['h00924] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00493] =  I0310077d53ae4ed9904df42e3f81c634['h00926] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00494] =  I0310077d53ae4ed9904df42e3f81c634['h00928] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00495] =  I0310077d53ae4ed9904df42e3f81c634['h0092a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00496] =  I0310077d53ae4ed9904df42e3f81c634['h0092c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00497] =  I0310077d53ae4ed9904df42e3f81c634['h0092e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00498] =  I0310077d53ae4ed9904df42e3f81c634['h00930] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00499] =  I0310077d53ae4ed9904df42e3f81c634['h00932] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0049a] =  I0310077d53ae4ed9904df42e3f81c634['h00934] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0049b] =  I0310077d53ae4ed9904df42e3f81c634['h00936] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0049c] =  I0310077d53ae4ed9904df42e3f81c634['h00938] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0049d] =  I0310077d53ae4ed9904df42e3f81c634['h0093a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0049e] =  I0310077d53ae4ed9904df42e3f81c634['h0093c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0049f] =  I0310077d53ae4ed9904df42e3f81c634['h0093e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a0] =  I0310077d53ae4ed9904df42e3f81c634['h00940] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a1] =  I0310077d53ae4ed9904df42e3f81c634['h00942] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a2] =  I0310077d53ae4ed9904df42e3f81c634['h00944] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a3] =  I0310077d53ae4ed9904df42e3f81c634['h00946] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a4] =  I0310077d53ae4ed9904df42e3f81c634['h00948] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a5] =  I0310077d53ae4ed9904df42e3f81c634['h0094a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a6] =  I0310077d53ae4ed9904df42e3f81c634['h0094c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a7] =  I0310077d53ae4ed9904df42e3f81c634['h0094e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a8] =  I0310077d53ae4ed9904df42e3f81c634['h00950] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004a9] =  I0310077d53ae4ed9904df42e3f81c634['h00952] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004aa] =  I0310077d53ae4ed9904df42e3f81c634['h00954] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ab] =  I0310077d53ae4ed9904df42e3f81c634['h00956] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ac] =  I0310077d53ae4ed9904df42e3f81c634['h00958] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ad] =  I0310077d53ae4ed9904df42e3f81c634['h0095a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ae] =  I0310077d53ae4ed9904df42e3f81c634['h0095c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004af] =  I0310077d53ae4ed9904df42e3f81c634['h0095e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b0] =  I0310077d53ae4ed9904df42e3f81c634['h00960] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b1] =  I0310077d53ae4ed9904df42e3f81c634['h00962] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b2] =  I0310077d53ae4ed9904df42e3f81c634['h00964] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b3] =  I0310077d53ae4ed9904df42e3f81c634['h00966] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b4] =  I0310077d53ae4ed9904df42e3f81c634['h00968] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b5] =  I0310077d53ae4ed9904df42e3f81c634['h0096a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b6] =  I0310077d53ae4ed9904df42e3f81c634['h0096c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b7] =  I0310077d53ae4ed9904df42e3f81c634['h0096e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b8] =  I0310077d53ae4ed9904df42e3f81c634['h00970] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004b9] =  I0310077d53ae4ed9904df42e3f81c634['h00972] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ba] =  I0310077d53ae4ed9904df42e3f81c634['h00974] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004bb] =  I0310077d53ae4ed9904df42e3f81c634['h00976] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004bc] =  I0310077d53ae4ed9904df42e3f81c634['h00978] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004bd] =  I0310077d53ae4ed9904df42e3f81c634['h0097a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004be] =  I0310077d53ae4ed9904df42e3f81c634['h0097c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004bf] =  I0310077d53ae4ed9904df42e3f81c634['h0097e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c0] =  I0310077d53ae4ed9904df42e3f81c634['h00980] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c1] =  I0310077d53ae4ed9904df42e3f81c634['h00982] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c2] =  I0310077d53ae4ed9904df42e3f81c634['h00984] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c3] =  I0310077d53ae4ed9904df42e3f81c634['h00986] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c4] =  I0310077d53ae4ed9904df42e3f81c634['h00988] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c5] =  I0310077d53ae4ed9904df42e3f81c634['h0098a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c6] =  I0310077d53ae4ed9904df42e3f81c634['h0098c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c7] =  I0310077d53ae4ed9904df42e3f81c634['h0098e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c8] =  I0310077d53ae4ed9904df42e3f81c634['h00990] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004c9] =  I0310077d53ae4ed9904df42e3f81c634['h00992] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ca] =  I0310077d53ae4ed9904df42e3f81c634['h00994] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004cb] =  I0310077d53ae4ed9904df42e3f81c634['h00996] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004cc] =  I0310077d53ae4ed9904df42e3f81c634['h00998] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004cd] =  I0310077d53ae4ed9904df42e3f81c634['h0099a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ce] =  I0310077d53ae4ed9904df42e3f81c634['h0099c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004cf] =  I0310077d53ae4ed9904df42e3f81c634['h0099e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d0] =  I0310077d53ae4ed9904df42e3f81c634['h009a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d1] =  I0310077d53ae4ed9904df42e3f81c634['h009a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d2] =  I0310077d53ae4ed9904df42e3f81c634['h009a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d3] =  I0310077d53ae4ed9904df42e3f81c634['h009a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d4] =  I0310077d53ae4ed9904df42e3f81c634['h009a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d5] =  I0310077d53ae4ed9904df42e3f81c634['h009aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d6] =  I0310077d53ae4ed9904df42e3f81c634['h009ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d7] =  I0310077d53ae4ed9904df42e3f81c634['h009ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d8] =  I0310077d53ae4ed9904df42e3f81c634['h009b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004d9] =  I0310077d53ae4ed9904df42e3f81c634['h009b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004da] =  I0310077d53ae4ed9904df42e3f81c634['h009b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004db] =  I0310077d53ae4ed9904df42e3f81c634['h009b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004dc] =  I0310077d53ae4ed9904df42e3f81c634['h009b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004dd] =  I0310077d53ae4ed9904df42e3f81c634['h009ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004de] =  I0310077d53ae4ed9904df42e3f81c634['h009bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004df] =  I0310077d53ae4ed9904df42e3f81c634['h009be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e0] =  I0310077d53ae4ed9904df42e3f81c634['h009c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e1] =  I0310077d53ae4ed9904df42e3f81c634['h009c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e2] =  I0310077d53ae4ed9904df42e3f81c634['h009c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e3] =  I0310077d53ae4ed9904df42e3f81c634['h009c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e4] =  I0310077d53ae4ed9904df42e3f81c634['h009c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e5] =  I0310077d53ae4ed9904df42e3f81c634['h009ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e6] =  I0310077d53ae4ed9904df42e3f81c634['h009cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e7] =  I0310077d53ae4ed9904df42e3f81c634['h009ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e8] =  I0310077d53ae4ed9904df42e3f81c634['h009d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004e9] =  I0310077d53ae4ed9904df42e3f81c634['h009d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ea] =  I0310077d53ae4ed9904df42e3f81c634['h009d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004eb] =  I0310077d53ae4ed9904df42e3f81c634['h009d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ec] =  I0310077d53ae4ed9904df42e3f81c634['h009d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ed] =  I0310077d53ae4ed9904df42e3f81c634['h009da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ee] =  I0310077d53ae4ed9904df42e3f81c634['h009dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ef] =  I0310077d53ae4ed9904df42e3f81c634['h009de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f0] =  I0310077d53ae4ed9904df42e3f81c634['h009e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f1] =  I0310077d53ae4ed9904df42e3f81c634['h009e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f2] =  I0310077d53ae4ed9904df42e3f81c634['h009e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f3] =  I0310077d53ae4ed9904df42e3f81c634['h009e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f4] =  I0310077d53ae4ed9904df42e3f81c634['h009e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f5] =  I0310077d53ae4ed9904df42e3f81c634['h009ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f6] =  I0310077d53ae4ed9904df42e3f81c634['h009ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f7] =  I0310077d53ae4ed9904df42e3f81c634['h009ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f8] =  I0310077d53ae4ed9904df42e3f81c634['h009f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004f9] =  I0310077d53ae4ed9904df42e3f81c634['h009f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004fa] =  I0310077d53ae4ed9904df42e3f81c634['h009f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004fb] =  I0310077d53ae4ed9904df42e3f81c634['h009f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004fc] =  I0310077d53ae4ed9904df42e3f81c634['h009f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004fd] =  I0310077d53ae4ed9904df42e3f81c634['h009fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004fe] =  I0310077d53ae4ed9904df42e3f81c634['h009fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h004ff] =  I0310077d53ae4ed9904df42e3f81c634['h009fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00500] =  I0310077d53ae4ed9904df42e3f81c634['h00a00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00501] =  I0310077d53ae4ed9904df42e3f81c634['h00a02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00502] =  I0310077d53ae4ed9904df42e3f81c634['h00a04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00503] =  I0310077d53ae4ed9904df42e3f81c634['h00a06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00504] =  I0310077d53ae4ed9904df42e3f81c634['h00a08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00505] =  I0310077d53ae4ed9904df42e3f81c634['h00a0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00506] =  I0310077d53ae4ed9904df42e3f81c634['h00a0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00507] =  I0310077d53ae4ed9904df42e3f81c634['h00a0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00508] =  I0310077d53ae4ed9904df42e3f81c634['h00a10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00509] =  I0310077d53ae4ed9904df42e3f81c634['h00a12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0050a] =  I0310077d53ae4ed9904df42e3f81c634['h00a14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0050b] =  I0310077d53ae4ed9904df42e3f81c634['h00a16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0050c] =  I0310077d53ae4ed9904df42e3f81c634['h00a18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0050d] =  I0310077d53ae4ed9904df42e3f81c634['h00a1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0050e] =  I0310077d53ae4ed9904df42e3f81c634['h00a1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0050f] =  I0310077d53ae4ed9904df42e3f81c634['h00a1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00510] =  I0310077d53ae4ed9904df42e3f81c634['h00a20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00511] =  I0310077d53ae4ed9904df42e3f81c634['h00a22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00512] =  I0310077d53ae4ed9904df42e3f81c634['h00a24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00513] =  I0310077d53ae4ed9904df42e3f81c634['h00a26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00514] =  I0310077d53ae4ed9904df42e3f81c634['h00a28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00515] =  I0310077d53ae4ed9904df42e3f81c634['h00a2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00516] =  I0310077d53ae4ed9904df42e3f81c634['h00a2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00517] =  I0310077d53ae4ed9904df42e3f81c634['h00a2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00518] =  I0310077d53ae4ed9904df42e3f81c634['h00a30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00519] =  I0310077d53ae4ed9904df42e3f81c634['h00a32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0051a] =  I0310077d53ae4ed9904df42e3f81c634['h00a34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0051b] =  I0310077d53ae4ed9904df42e3f81c634['h00a36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0051c] =  I0310077d53ae4ed9904df42e3f81c634['h00a38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0051d] =  I0310077d53ae4ed9904df42e3f81c634['h00a3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0051e] =  I0310077d53ae4ed9904df42e3f81c634['h00a3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0051f] =  I0310077d53ae4ed9904df42e3f81c634['h00a3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00520] =  I0310077d53ae4ed9904df42e3f81c634['h00a40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00521] =  I0310077d53ae4ed9904df42e3f81c634['h00a42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00522] =  I0310077d53ae4ed9904df42e3f81c634['h00a44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00523] =  I0310077d53ae4ed9904df42e3f81c634['h00a46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00524] =  I0310077d53ae4ed9904df42e3f81c634['h00a48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00525] =  I0310077d53ae4ed9904df42e3f81c634['h00a4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00526] =  I0310077d53ae4ed9904df42e3f81c634['h00a4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00527] =  I0310077d53ae4ed9904df42e3f81c634['h00a4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00528] =  I0310077d53ae4ed9904df42e3f81c634['h00a50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00529] =  I0310077d53ae4ed9904df42e3f81c634['h00a52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0052a] =  I0310077d53ae4ed9904df42e3f81c634['h00a54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0052b] =  I0310077d53ae4ed9904df42e3f81c634['h00a56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0052c] =  I0310077d53ae4ed9904df42e3f81c634['h00a58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0052d] =  I0310077d53ae4ed9904df42e3f81c634['h00a5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0052e] =  I0310077d53ae4ed9904df42e3f81c634['h00a5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0052f] =  I0310077d53ae4ed9904df42e3f81c634['h00a5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00530] =  I0310077d53ae4ed9904df42e3f81c634['h00a60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00531] =  I0310077d53ae4ed9904df42e3f81c634['h00a62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00532] =  I0310077d53ae4ed9904df42e3f81c634['h00a64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00533] =  I0310077d53ae4ed9904df42e3f81c634['h00a66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00534] =  I0310077d53ae4ed9904df42e3f81c634['h00a68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00535] =  I0310077d53ae4ed9904df42e3f81c634['h00a6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00536] =  I0310077d53ae4ed9904df42e3f81c634['h00a6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00537] =  I0310077d53ae4ed9904df42e3f81c634['h00a6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00538] =  I0310077d53ae4ed9904df42e3f81c634['h00a70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00539] =  I0310077d53ae4ed9904df42e3f81c634['h00a72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0053a] =  I0310077d53ae4ed9904df42e3f81c634['h00a74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0053b] =  I0310077d53ae4ed9904df42e3f81c634['h00a76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0053c] =  I0310077d53ae4ed9904df42e3f81c634['h00a78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0053d] =  I0310077d53ae4ed9904df42e3f81c634['h00a7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0053e] =  I0310077d53ae4ed9904df42e3f81c634['h00a7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0053f] =  I0310077d53ae4ed9904df42e3f81c634['h00a7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00540] =  I0310077d53ae4ed9904df42e3f81c634['h00a80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00541] =  I0310077d53ae4ed9904df42e3f81c634['h00a82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00542] =  I0310077d53ae4ed9904df42e3f81c634['h00a84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00543] =  I0310077d53ae4ed9904df42e3f81c634['h00a86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00544] =  I0310077d53ae4ed9904df42e3f81c634['h00a88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00545] =  I0310077d53ae4ed9904df42e3f81c634['h00a8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00546] =  I0310077d53ae4ed9904df42e3f81c634['h00a8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00547] =  I0310077d53ae4ed9904df42e3f81c634['h00a8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00548] =  I0310077d53ae4ed9904df42e3f81c634['h00a90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00549] =  I0310077d53ae4ed9904df42e3f81c634['h00a92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0054a] =  I0310077d53ae4ed9904df42e3f81c634['h00a94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0054b] =  I0310077d53ae4ed9904df42e3f81c634['h00a96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0054c] =  I0310077d53ae4ed9904df42e3f81c634['h00a98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0054d] =  I0310077d53ae4ed9904df42e3f81c634['h00a9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0054e] =  I0310077d53ae4ed9904df42e3f81c634['h00a9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0054f] =  I0310077d53ae4ed9904df42e3f81c634['h00a9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00550] =  I0310077d53ae4ed9904df42e3f81c634['h00aa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00551] =  I0310077d53ae4ed9904df42e3f81c634['h00aa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00552] =  I0310077d53ae4ed9904df42e3f81c634['h00aa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00553] =  I0310077d53ae4ed9904df42e3f81c634['h00aa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00554] =  I0310077d53ae4ed9904df42e3f81c634['h00aa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00555] =  I0310077d53ae4ed9904df42e3f81c634['h00aaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00556] =  I0310077d53ae4ed9904df42e3f81c634['h00aac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00557] =  I0310077d53ae4ed9904df42e3f81c634['h00aae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00558] =  I0310077d53ae4ed9904df42e3f81c634['h00ab0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00559] =  I0310077d53ae4ed9904df42e3f81c634['h00ab2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0055a] =  I0310077d53ae4ed9904df42e3f81c634['h00ab4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0055b] =  I0310077d53ae4ed9904df42e3f81c634['h00ab6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0055c] =  I0310077d53ae4ed9904df42e3f81c634['h00ab8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0055d] =  I0310077d53ae4ed9904df42e3f81c634['h00aba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0055e] =  I0310077d53ae4ed9904df42e3f81c634['h00abc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0055f] =  I0310077d53ae4ed9904df42e3f81c634['h00abe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00560] =  I0310077d53ae4ed9904df42e3f81c634['h00ac0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00561] =  I0310077d53ae4ed9904df42e3f81c634['h00ac2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00562] =  I0310077d53ae4ed9904df42e3f81c634['h00ac4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00563] =  I0310077d53ae4ed9904df42e3f81c634['h00ac6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00564] =  I0310077d53ae4ed9904df42e3f81c634['h00ac8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00565] =  I0310077d53ae4ed9904df42e3f81c634['h00aca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00566] =  I0310077d53ae4ed9904df42e3f81c634['h00acc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00567] =  I0310077d53ae4ed9904df42e3f81c634['h00ace] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00568] =  I0310077d53ae4ed9904df42e3f81c634['h00ad0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00569] =  I0310077d53ae4ed9904df42e3f81c634['h00ad2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0056a] =  I0310077d53ae4ed9904df42e3f81c634['h00ad4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0056b] =  I0310077d53ae4ed9904df42e3f81c634['h00ad6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0056c] =  I0310077d53ae4ed9904df42e3f81c634['h00ad8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0056d] =  I0310077d53ae4ed9904df42e3f81c634['h00ada] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0056e] =  I0310077d53ae4ed9904df42e3f81c634['h00adc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0056f] =  I0310077d53ae4ed9904df42e3f81c634['h00ade] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00570] =  I0310077d53ae4ed9904df42e3f81c634['h00ae0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00571] =  I0310077d53ae4ed9904df42e3f81c634['h00ae2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00572] =  I0310077d53ae4ed9904df42e3f81c634['h00ae4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00573] =  I0310077d53ae4ed9904df42e3f81c634['h00ae6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00574] =  I0310077d53ae4ed9904df42e3f81c634['h00ae8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00575] =  I0310077d53ae4ed9904df42e3f81c634['h00aea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00576] =  I0310077d53ae4ed9904df42e3f81c634['h00aec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00577] =  I0310077d53ae4ed9904df42e3f81c634['h00aee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00578] =  I0310077d53ae4ed9904df42e3f81c634['h00af0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00579] =  I0310077d53ae4ed9904df42e3f81c634['h00af2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0057a] =  I0310077d53ae4ed9904df42e3f81c634['h00af4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0057b] =  I0310077d53ae4ed9904df42e3f81c634['h00af6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0057c] =  I0310077d53ae4ed9904df42e3f81c634['h00af8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0057d] =  I0310077d53ae4ed9904df42e3f81c634['h00afa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0057e] =  I0310077d53ae4ed9904df42e3f81c634['h00afc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0057f] =  I0310077d53ae4ed9904df42e3f81c634['h00afe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00580] =  I0310077d53ae4ed9904df42e3f81c634['h00b00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00581] =  I0310077d53ae4ed9904df42e3f81c634['h00b02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00582] =  I0310077d53ae4ed9904df42e3f81c634['h00b04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00583] =  I0310077d53ae4ed9904df42e3f81c634['h00b06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00584] =  I0310077d53ae4ed9904df42e3f81c634['h00b08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00585] =  I0310077d53ae4ed9904df42e3f81c634['h00b0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00586] =  I0310077d53ae4ed9904df42e3f81c634['h00b0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00587] =  I0310077d53ae4ed9904df42e3f81c634['h00b0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00588] =  I0310077d53ae4ed9904df42e3f81c634['h00b10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00589] =  I0310077d53ae4ed9904df42e3f81c634['h00b12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0058a] =  I0310077d53ae4ed9904df42e3f81c634['h00b14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0058b] =  I0310077d53ae4ed9904df42e3f81c634['h00b16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0058c] =  I0310077d53ae4ed9904df42e3f81c634['h00b18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0058d] =  I0310077d53ae4ed9904df42e3f81c634['h00b1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0058e] =  I0310077d53ae4ed9904df42e3f81c634['h00b1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0058f] =  I0310077d53ae4ed9904df42e3f81c634['h00b1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00590] =  I0310077d53ae4ed9904df42e3f81c634['h00b20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00591] =  I0310077d53ae4ed9904df42e3f81c634['h00b22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00592] =  I0310077d53ae4ed9904df42e3f81c634['h00b24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00593] =  I0310077d53ae4ed9904df42e3f81c634['h00b26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00594] =  I0310077d53ae4ed9904df42e3f81c634['h00b28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00595] =  I0310077d53ae4ed9904df42e3f81c634['h00b2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00596] =  I0310077d53ae4ed9904df42e3f81c634['h00b2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00597] =  I0310077d53ae4ed9904df42e3f81c634['h00b2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00598] =  I0310077d53ae4ed9904df42e3f81c634['h00b30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00599] =  I0310077d53ae4ed9904df42e3f81c634['h00b32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0059a] =  I0310077d53ae4ed9904df42e3f81c634['h00b34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0059b] =  I0310077d53ae4ed9904df42e3f81c634['h00b36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0059c] =  I0310077d53ae4ed9904df42e3f81c634['h00b38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0059d] =  I0310077d53ae4ed9904df42e3f81c634['h00b3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0059e] =  I0310077d53ae4ed9904df42e3f81c634['h00b3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0059f] =  I0310077d53ae4ed9904df42e3f81c634['h00b3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a0] =  I0310077d53ae4ed9904df42e3f81c634['h00b40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a1] =  I0310077d53ae4ed9904df42e3f81c634['h00b42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a2] =  I0310077d53ae4ed9904df42e3f81c634['h00b44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a3] =  I0310077d53ae4ed9904df42e3f81c634['h00b46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a4] =  I0310077d53ae4ed9904df42e3f81c634['h00b48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a5] =  I0310077d53ae4ed9904df42e3f81c634['h00b4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a6] =  I0310077d53ae4ed9904df42e3f81c634['h00b4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a7] =  I0310077d53ae4ed9904df42e3f81c634['h00b4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a8] =  I0310077d53ae4ed9904df42e3f81c634['h00b50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005a9] =  I0310077d53ae4ed9904df42e3f81c634['h00b52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005aa] =  I0310077d53ae4ed9904df42e3f81c634['h00b54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ab] =  I0310077d53ae4ed9904df42e3f81c634['h00b56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ac] =  I0310077d53ae4ed9904df42e3f81c634['h00b58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ad] =  I0310077d53ae4ed9904df42e3f81c634['h00b5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ae] =  I0310077d53ae4ed9904df42e3f81c634['h00b5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005af] =  I0310077d53ae4ed9904df42e3f81c634['h00b5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b0] =  I0310077d53ae4ed9904df42e3f81c634['h00b60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b1] =  I0310077d53ae4ed9904df42e3f81c634['h00b62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b2] =  I0310077d53ae4ed9904df42e3f81c634['h00b64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b3] =  I0310077d53ae4ed9904df42e3f81c634['h00b66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b4] =  I0310077d53ae4ed9904df42e3f81c634['h00b68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b5] =  I0310077d53ae4ed9904df42e3f81c634['h00b6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b6] =  I0310077d53ae4ed9904df42e3f81c634['h00b6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b7] =  I0310077d53ae4ed9904df42e3f81c634['h00b6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b8] =  I0310077d53ae4ed9904df42e3f81c634['h00b70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005b9] =  I0310077d53ae4ed9904df42e3f81c634['h00b72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ba] =  I0310077d53ae4ed9904df42e3f81c634['h00b74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005bb] =  I0310077d53ae4ed9904df42e3f81c634['h00b76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005bc] =  I0310077d53ae4ed9904df42e3f81c634['h00b78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005bd] =  I0310077d53ae4ed9904df42e3f81c634['h00b7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005be] =  I0310077d53ae4ed9904df42e3f81c634['h00b7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005bf] =  I0310077d53ae4ed9904df42e3f81c634['h00b7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c0] =  I0310077d53ae4ed9904df42e3f81c634['h00b80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c1] =  I0310077d53ae4ed9904df42e3f81c634['h00b82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c2] =  I0310077d53ae4ed9904df42e3f81c634['h00b84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c3] =  I0310077d53ae4ed9904df42e3f81c634['h00b86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c4] =  I0310077d53ae4ed9904df42e3f81c634['h00b88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c5] =  I0310077d53ae4ed9904df42e3f81c634['h00b8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c6] =  I0310077d53ae4ed9904df42e3f81c634['h00b8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c7] =  I0310077d53ae4ed9904df42e3f81c634['h00b8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c8] =  I0310077d53ae4ed9904df42e3f81c634['h00b90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005c9] =  I0310077d53ae4ed9904df42e3f81c634['h00b92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ca] =  I0310077d53ae4ed9904df42e3f81c634['h00b94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005cb] =  I0310077d53ae4ed9904df42e3f81c634['h00b96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005cc] =  I0310077d53ae4ed9904df42e3f81c634['h00b98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005cd] =  I0310077d53ae4ed9904df42e3f81c634['h00b9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ce] =  I0310077d53ae4ed9904df42e3f81c634['h00b9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005cf] =  I0310077d53ae4ed9904df42e3f81c634['h00b9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d0] =  I0310077d53ae4ed9904df42e3f81c634['h00ba0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d1] =  I0310077d53ae4ed9904df42e3f81c634['h00ba2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d2] =  I0310077d53ae4ed9904df42e3f81c634['h00ba4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d3] =  I0310077d53ae4ed9904df42e3f81c634['h00ba6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d4] =  I0310077d53ae4ed9904df42e3f81c634['h00ba8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d5] =  I0310077d53ae4ed9904df42e3f81c634['h00baa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d6] =  I0310077d53ae4ed9904df42e3f81c634['h00bac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d7] =  I0310077d53ae4ed9904df42e3f81c634['h00bae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d8] =  I0310077d53ae4ed9904df42e3f81c634['h00bb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005d9] =  I0310077d53ae4ed9904df42e3f81c634['h00bb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005da] =  I0310077d53ae4ed9904df42e3f81c634['h00bb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005db] =  I0310077d53ae4ed9904df42e3f81c634['h00bb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005dc] =  I0310077d53ae4ed9904df42e3f81c634['h00bb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005dd] =  I0310077d53ae4ed9904df42e3f81c634['h00bba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005de] =  I0310077d53ae4ed9904df42e3f81c634['h00bbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005df] =  I0310077d53ae4ed9904df42e3f81c634['h00bbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e0] =  I0310077d53ae4ed9904df42e3f81c634['h00bc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e1] =  I0310077d53ae4ed9904df42e3f81c634['h00bc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e2] =  I0310077d53ae4ed9904df42e3f81c634['h00bc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e3] =  I0310077d53ae4ed9904df42e3f81c634['h00bc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e4] =  I0310077d53ae4ed9904df42e3f81c634['h00bc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e5] =  I0310077d53ae4ed9904df42e3f81c634['h00bca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e6] =  I0310077d53ae4ed9904df42e3f81c634['h00bcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e7] =  I0310077d53ae4ed9904df42e3f81c634['h00bce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e8] =  I0310077d53ae4ed9904df42e3f81c634['h00bd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005e9] =  I0310077d53ae4ed9904df42e3f81c634['h00bd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ea] =  I0310077d53ae4ed9904df42e3f81c634['h00bd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005eb] =  I0310077d53ae4ed9904df42e3f81c634['h00bd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ec] =  I0310077d53ae4ed9904df42e3f81c634['h00bd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ed] =  I0310077d53ae4ed9904df42e3f81c634['h00bda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ee] =  I0310077d53ae4ed9904df42e3f81c634['h00bdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ef] =  I0310077d53ae4ed9904df42e3f81c634['h00bde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f0] =  I0310077d53ae4ed9904df42e3f81c634['h00be0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f1] =  I0310077d53ae4ed9904df42e3f81c634['h00be2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f2] =  I0310077d53ae4ed9904df42e3f81c634['h00be4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f3] =  I0310077d53ae4ed9904df42e3f81c634['h00be6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f4] =  I0310077d53ae4ed9904df42e3f81c634['h00be8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f5] =  I0310077d53ae4ed9904df42e3f81c634['h00bea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f6] =  I0310077d53ae4ed9904df42e3f81c634['h00bec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f7] =  I0310077d53ae4ed9904df42e3f81c634['h00bee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f8] =  I0310077d53ae4ed9904df42e3f81c634['h00bf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005f9] =  I0310077d53ae4ed9904df42e3f81c634['h00bf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005fa] =  I0310077d53ae4ed9904df42e3f81c634['h00bf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005fb] =  I0310077d53ae4ed9904df42e3f81c634['h00bf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005fc] =  I0310077d53ae4ed9904df42e3f81c634['h00bf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005fd] =  I0310077d53ae4ed9904df42e3f81c634['h00bfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005fe] =  I0310077d53ae4ed9904df42e3f81c634['h00bfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h005ff] =  I0310077d53ae4ed9904df42e3f81c634['h00bfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00600] =  I0310077d53ae4ed9904df42e3f81c634['h00c00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00601] =  I0310077d53ae4ed9904df42e3f81c634['h00c02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00602] =  I0310077d53ae4ed9904df42e3f81c634['h00c04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00603] =  I0310077d53ae4ed9904df42e3f81c634['h00c06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00604] =  I0310077d53ae4ed9904df42e3f81c634['h00c08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00605] =  I0310077d53ae4ed9904df42e3f81c634['h00c0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00606] =  I0310077d53ae4ed9904df42e3f81c634['h00c0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00607] =  I0310077d53ae4ed9904df42e3f81c634['h00c0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00608] =  I0310077d53ae4ed9904df42e3f81c634['h00c10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00609] =  I0310077d53ae4ed9904df42e3f81c634['h00c12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0060a] =  I0310077d53ae4ed9904df42e3f81c634['h00c14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0060b] =  I0310077d53ae4ed9904df42e3f81c634['h00c16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0060c] =  I0310077d53ae4ed9904df42e3f81c634['h00c18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0060d] =  I0310077d53ae4ed9904df42e3f81c634['h00c1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0060e] =  I0310077d53ae4ed9904df42e3f81c634['h00c1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0060f] =  I0310077d53ae4ed9904df42e3f81c634['h00c1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00610] =  I0310077d53ae4ed9904df42e3f81c634['h00c20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00611] =  I0310077d53ae4ed9904df42e3f81c634['h00c22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00612] =  I0310077d53ae4ed9904df42e3f81c634['h00c24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00613] =  I0310077d53ae4ed9904df42e3f81c634['h00c26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00614] =  I0310077d53ae4ed9904df42e3f81c634['h00c28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00615] =  I0310077d53ae4ed9904df42e3f81c634['h00c2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00616] =  I0310077d53ae4ed9904df42e3f81c634['h00c2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00617] =  I0310077d53ae4ed9904df42e3f81c634['h00c2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00618] =  I0310077d53ae4ed9904df42e3f81c634['h00c30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00619] =  I0310077d53ae4ed9904df42e3f81c634['h00c32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0061a] =  I0310077d53ae4ed9904df42e3f81c634['h00c34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0061b] =  I0310077d53ae4ed9904df42e3f81c634['h00c36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0061c] =  I0310077d53ae4ed9904df42e3f81c634['h00c38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0061d] =  I0310077d53ae4ed9904df42e3f81c634['h00c3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0061e] =  I0310077d53ae4ed9904df42e3f81c634['h00c3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0061f] =  I0310077d53ae4ed9904df42e3f81c634['h00c3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00620] =  I0310077d53ae4ed9904df42e3f81c634['h00c40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00621] =  I0310077d53ae4ed9904df42e3f81c634['h00c42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00622] =  I0310077d53ae4ed9904df42e3f81c634['h00c44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00623] =  I0310077d53ae4ed9904df42e3f81c634['h00c46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00624] =  I0310077d53ae4ed9904df42e3f81c634['h00c48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00625] =  I0310077d53ae4ed9904df42e3f81c634['h00c4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00626] =  I0310077d53ae4ed9904df42e3f81c634['h00c4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00627] =  I0310077d53ae4ed9904df42e3f81c634['h00c4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00628] =  I0310077d53ae4ed9904df42e3f81c634['h00c50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00629] =  I0310077d53ae4ed9904df42e3f81c634['h00c52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0062a] =  I0310077d53ae4ed9904df42e3f81c634['h00c54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0062b] =  I0310077d53ae4ed9904df42e3f81c634['h00c56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0062c] =  I0310077d53ae4ed9904df42e3f81c634['h00c58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0062d] =  I0310077d53ae4ed9904df42e3f81c634['h00c5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0062e] =  I0310077d53ae4ed9904df42e3f81c634['h00c5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0062f] =  I0310077d53ae4ed9904df42e3f81c634['h00c5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00630] =  I0310077d53ae4ed9904df42e3f81c634['h00c60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00631] =  I0310077d53ae4ed9904df42e3f81c634['h00c62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00632] =  I0310077d53ae4ed9904df42e3f81c634['h00c64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00633] =  I0310077d53ae4ed9904df42e3f81c634['h00c66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00634] =  I0310077d53ae4ed9904df42e3f81c634['h00c68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00635] =  I0310077d53ae4ed9904df42e3f81c634['h00c6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00636] =  I0310077d53ae4ed9904df42e3f81c634['h00c6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00637] =  I0310077d53ae4ed9904df42e3f81c634['h00c6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00638] =  I0310077d53ae4ed9904df42e3f81c634['h00c70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00639] =  I0310077d53ae4ed9904df42e3f81c634['h00c72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0063a] =  I0310077d53ae4ed9904df42e3f81c634['h00c74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0063b] =  I0310077d53ae4ed9904df42e3f81c634['h00c76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0063c] =  I0310077d53ae4ed9904df42e3f81c634['h00c78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0063d] =  I0310077d53ae4ed9904df42e3f81c634['h00c7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0063e] =  I0310077d53ae4ed9904df42e3f81c634['h00c7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0063f] =  I0310077d53ae4ed9904df42e3f81c634['h00c7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00640] =  I0310077d53ae4ed9904df42e3f81c634['h00c80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00641] =  I0310077d53ae4ed9904df42e3f81c634['h00c82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00642] =  I0310077d53ae4ed9904df42e3f81c634['h00c84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00643] =  I0310077d53ae4ed9904df42e3f81c634['h00c86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00644] =  I0310077d53ae4ed9904df42e3f81c634['h00c88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00645] =  I0310077d53ae4ed9904df42e3f81c634['h00c8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00646] =  I0310077d53ae4ed9904df42e3f81c634['h00c8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00647] =  I0310077d53ae4ed9904df42e3f81c634['h00c8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00648] =  I0310077d53ae4ed9904df42e3f81c634['h00c90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00649] =  I0310077d53ae4ed9904df42e3f81c634['h00c92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0064a] =  I0310077d53ae4ed9904df42e3f81c634['h00c94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0064b] =  I0310077d53ae4ed9904df42e3f81c634['h00c96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0064c] =  I0310077d53ae4ed9904df42e3f81c634['h00c98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0064d] =  I0310077d53ae4ed9904df42e3f81c634['h00c9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0064e] =  I0310077d53ae4ed9904df42e3f81c634['h00c9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0064f] =  I0310077d53ae4ed9904df42e3f81c634['h00c9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00650] =  I0310077d53ae4ed9904df42e3f81c634['h00ca0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00651] =  I0310077d53ae4ed9904df42e3f81c634['h00ca2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00652] =  I0310077d53ae4ed9904df42e3f81c634['h00ca4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00653] =  I0310077d53ae4ed9904df42e3f81c634['h00ca6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00654] =  I0310077d53ae4ed9904df42e3f81c634['h00ca8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00655] =  I0310077d53ae4ed9904df42e3f81c634['h00caa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00656] =  I0310077d53ae4ed9904df42e3f81c634['h00cac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00657] =  I0310077d53ae4ed9904df42e3f81c634['h00cae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00658] =  I0310077d53ae4ed9904df42e3f81c634['h00cb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00659] =  I0310077d53ae4ed9904df42e3f81c634['h00cb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0065a] =  I0310077d53ae4ed9904df42e3f81c634['h00cb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0065b] =  I0310077d53ae4ed9904df42e3f81c634['h00cb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0065c] =  I0310077d53ae4ed9904df42e3f81c634['h00cb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0065d] =  I0310077d53ae4ed9904df42e3f81c634['h00cba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0065e] =  I0310077d53ae4ed9904df42e3f81c634['h00cbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0065f] =  I0310077d53ae4ed9904df42e3f81c634['h00cbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00660] =  I0310077d53ae4ed9904df42e3f81c634['h00cc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00661] =  I0310077d53ae4ed9904df42e3f81c634['h00cc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00662] =  I0310077d53ae4ed9904df42e3f81c634['h00cc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00663] =  I0310077d53ae4ed9904df42e3f81c634['h00cc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00664] =  I0310077d53ae4ed9904df42e3f81c634['h00cc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00665] =  I0310077d53ae4ed9904df42e3f81c634['h00cca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00666] =  I0310077d53ae4ed9904df42e3f81c634['h00ccc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00667] =  I0310077d53ae4ed9904df42e3f81c634['h00cce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00668] =  I0310077d53ae4ed9904df42e3f81c634['h00cd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00669] =  I0310077d53ae4ed9904df42e3f81c634['h00cd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0066a] =  I0310077d53ae4ed9904df42e3f81c634['h00cd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0066b] =  I0310077d53ae4ed9904df42e3f81c634['h00cd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0066c] =  I0310077d53ae4ed9904df42e3f81c634['h00cd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0066d] =  I0310077d53ae4ed9904df42e3f81c634['h00cda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0066e] =  I0310077d53ae4ed9904df42e3f81c634['h00cdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0066f] =  I0310077d53ae4ed9904df42e3f81c634['h00cde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00670] =  I0310077d53ae4ed9904df42e3f81c634['h00ce0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00671] =  I0310077d53ae4ed9904df42e3f81c634['h00ce2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00672] =  I0310077d53ae4ed9904df42e3f81c634['h00ce4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00673] =  I0310077d53ae4ed9904df42e3f81c634['h00ce6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00674] =  I0310077d53ae4ed9904df42e3f81c634['h00ce8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00675] =  I0310077d53ae4ed9904df42e3f81c634['h00cea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00676] =  I0310077d53ae4ed9904df42e3f81c634['h00cec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00677] =  I0310077d53ae4ed9904df42e3f81c634['h00cee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00678] =  I0310077d53ae4ed9904df42e3f81c634['h00cf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00679] =  I0310077d53ae4ed9904df42e3f81c634['h00cf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0067a] =  I0310077d53ae4ed9904df42e3f81c634['h00cf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0067b] =  I0310077d53ae4ed9904df42e3f81c634['h00cf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0067c] =  I0310077d53ae4ed9904df42e3f81c634['h00cf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0067d] =  I0310077d53ae4ed9904df42e3f81c634['h00cfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0067e] =  I0310077d53ae4ed9904df42e3f81c634['h00cfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0067f] =  I0310077d53ae4ed9904df42e3f81c634['h00cfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00680] =  I0310077d53ae4ed9904df42e3f81c634['h00d00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00681] =  I0310077d53ae4ed9904df42e3f81c634['h00d02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00682] =  I0310077d53ae4ed9904df42e3f81c634['h00d04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00683] =  I0310077d53ae4ed9904df42e3f81c634['h00d06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00684] =  I0310077d53ae4ed9904df42e3f81c634['h00d08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00685] =  I0310077d53ae4ed9904df42e3f81c634['h00d0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00686] =  I0310077d53ae4ed9904df42e3f81c634['h00d0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00687] =  I0310077d53ae4ed9904df42e3f81c634['h00d0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00688] =  I0310077d53ae4ed9904df42e3f81c634['h00d10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00689] =  I0310077d53ae4ed9904df42e3f81c634['h00d12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0068a] =  I0310077d53ae4ed9904df42e3f81c634['h00d14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0068b] =  I0310077d53ae4ed9904df42e3f81c634['h00d16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0068c] =  I0310077d53ae4ed9904df42e3f81c634['h00d18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0068d] =  I0310077d53ae4ed9904df42e3f81c634['h00d1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0068e] =  I0310077d53ae4ed9904df42e3f81c634['h00d1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0068f] =  I0310077d53ae4ed9904df42e3f81c634['h00d1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00690] =  I0310077d53ae4ed9904df42e3f81c634['h00d20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00691] =  I0310077d53ae4ed9904df42e3f81c634['h00d22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00692] =  I0310077d53ae4ed9904df42e3f81c634['h00d24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00693] =  I0310077d53ae4ed9904df42e3f81c634['h00d26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00694] =  I0310077d53ae4ed9904df42e3f81c634['h00d28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00695] =  I0310077d53ae4ed9904df42e3f81c634['h00d2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00696] =  I0310077d53ae4ed9904df42e3f81c634['h00d2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00697] =  I0310077d53ae4ed9904df42e3f81c634['h00d2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00698] =  I0310077d53ae4ed9904df42e3f81c634['h00d30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00699] =  I0310077d53ae4ed9904df42e3f81c634['h00d32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0069a] =  I0310077d53ae4ed9904df42e3f81c634['h00d34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0069b] =  I0310077d53ae4ed9904df42e3f81c634['h00d36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0069c] =  I0310077d53ae4ed9904df42e3f81c634['h00d38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0069d] =  I0310077d53ae4ed9904df42e3f81c634['h00d3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0069e] =  I0310077d53ae4ed9904df42e3f81c634['h00d3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0069f] =  I0310077d53ae4ed9904df42e3f81c634['h00d3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a0] =  I0310077d53ae4ed9904df42e3f81c634['h00d40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a1] =  I0310077d53ae4ed9904df42e3f81c634['h00d42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a2] =  I0310077d53ae4ed9904df42e3f81c634['h00d44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a3] =  I0310077d53ae4ed9904df42e3f81c634['h00d46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a4] =  I0310077d53ae4ed9904df42e3f81c634['h00d48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a5] =  I0310077d53ae4ed9904df42e3f81c634['h00d4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a6] =  I0310077d53ae4ed9904df42e3f81c634['h00d4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a7] =  I0310077d53ae4ed9904df42e3f81c634['h00d4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a8] =  I0310077d53ae4ed9904df42e3f81c634['h00d50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006a9] =  I0310077d53ae4ed9904df42e3f81c634['h00d52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006aa] =  I0310077d53ae4ed9904df42e3f81c634['h00d54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ab] =  I0310077d53ae4ed9904df42e3f81c634['h00d56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ac] =  I0310077d53ae4ed9904df42e3f81c634['h00d58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ad] =  I0310077d53ae4ed9904df42e3f81c634['h00d5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ae] =  I0310077d53ae4ed9904df42e3f81c634['h00d5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006af] =  I0310077d53ae4ed9904df42e3f81c634['h00d5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b0] =  I0310077d53ae4ed9904df42e3f81c634['h00d60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b1] =  I0310077d53ae4ed9904df42e3f81c634['h00d62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b2] =  I0310077d53ae4ed9904df42e3f81c634['h00d64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b3] =  I0310077d53ae4ed9904df42e3f81c634['h00d66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b4] =  I0310077d53ae4ed9904df42e3f81c634['h00d68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b5] =  I0310077d53ae4ed9904df42e3f81c634['h00d6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b6] =  I0310077d53ae4ed9904df42e3f81c634['h00d6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b7] =  I0310077d53ae4ed9904df42e3f81c634['h00d6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b8] =  I0310077d53ae4ed9904df42e3f81c634['h00d70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006b9] =  I0310077d53ae4ed9904df42e3f81c634['h00d72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ba] =  I0310077d53ae4ed9904df42e3f81c634['h00d74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006bb] =  I0310077d53ae4ed9904df42e3f81c634['h00d76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006bc] =  I0310077d53ae4ed9904df42e3f81c634['h00d78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006bd] =  I0310077d53ae4ed9904df42e3f81c634['h00d7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006be] =  I0310077d53ae4ed9904df42e3f81c634['h00d7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006bf] =  I0310077d53ae4ed9904df42e3f81c634['h00d7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c0] =  I0310077d53ae4ed9904df42e3f81c634['h00d80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c1] =  I0310077d53ae4ed9904df42e3f81c634['h00d82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c2] =  I0310077d53ae4ed9904df42e3f81c634['h00d84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c3] =  I0310077d53ae4ed9904df42e3f81c634['h00d86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c4] =  I0310077d53ae4ed9904df42e3f81c634['h00d88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c5] =  I0310077d53ae4ed9904df42e3f81c634['h00d8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c6] =  I0310077d53ae4ed9904df42e3f81c634['h00d8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c7] =  I0310077d53ae4ed9904df42e3f81c634['h00d8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c8] =  I0310077d53ae4ed9904df42e3f81c634['h00d90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006c9] =  I0310077d53ae4ed9904df42e3f81c634['h00d92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ca] =  I0310077d53ae4ed9904df42e3f81c634['h00d94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006cb] =  I0310077d53ae4ed9904df42e3f81c634['h00d96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006cc] =  I0310077d53ae4ed9904df42e3f81c634['h00d98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006cd] =  I0310077d53ae4ed9904df42e3f81c634['h00d9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ce] =  I0310077d53ae4ed9904df42e3f81c634['h00d9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006cf] =  I0310077d53ae4ed9904df42e3f81c634['h00d9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d0] =  I0310077d53ae4ed9904df42e3f81c634['h00da0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d1] =  I0310077d53ae4ed9904df42e3f81c634['h00da2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d2] =  I0310077d53ae4ed9904df42e3f81c634['h00da4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d3] =  I0310077d53ae4ed9904df42e3f81c634['h00da6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d4] =  I0310077d53ae4ed9904df42e3f81c634['h00da8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d5] =  I0310077d53ae4ed9904df42e3f81c634['h00daa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d6] =  I0310077d53ae4ed9904df42e3f81c634['h00dac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d7] =  I0310077d53ae4ed9904df42e3f81c634['h00dae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d8] =  I0310077d53ae4ed9904df42e3f81c634['h00db0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006d9] =  I0310077d53ae4ed9904df42e3f81c634['h00db2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006da] =  I0310077d53ae4ed9904df42e3f81c634['h00db4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006db] =  I0310077d53ae4ed9904df42e3f81c634['h00db6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006dc] =  I0310077d53ae4ed9904df42e3f81c634['h00db8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006dd] =  I0310077d53ae4ed9904df42e3f81c634['h00dba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006de] =  I0310077d53ae4ed9904df42e3f81c634['h00dbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006df] =  I0310077d53ae4ed9904df42e3f81c634['h00dbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e0] =  I0310077d53ae4ed9904df42e3f81c634['h00dc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e1] =  I0310077d53ae4ed9904df42e3f81c634['h00dc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e2] =  I0310077d53ae4ed9904df42e3f81c634['h00dc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e3] =  I0310077d53ae4ed9904df42e3f81c634['h00dc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e4] =  I0310077d53ae4ed9904df42e3f81c634['h00dc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e5] =  I0310077d53ae4ed9904df42e3f81c634['h00dca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e6] =  I0310077d53ae4ed9904df42e3f81c634['h00dcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e7] =  I0310077d53ae4ed9904df42e3f81c634['h00dce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e8] =  I0310077d53ae4ed9904df42e3f81c634['h00dd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006e9] =  I0310077d53ae4ed9904df42e3f81c634['h00dd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ea] =  I0310077d53ae4ed9904df42e3f81c634['h00dd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006eb] =  I0310077d53ae4ed9904df42e3f81c634['h00dd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ec] =  I0310077d53ae4ed9904df42e3f81c634['h00dd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ed] =  I0310077d53ae4ed9904df42e3f81c634['h00dda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ee] =  I0310077d53ae4ed9904df42e3f81c634['h00ddc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ef] =  I0310077d53ae4ed9904df42e3f81c634['h00dde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f0] =  I0310077d53ae4ed9904df42e3f81c634['h00de0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f1] =  I0310077d53ae4ed9904df42e3f81c634['h00de2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f2] =  I0310077d53ae4ed9904df42e3f81c634['h00de4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f3] =  I0310077d53ae4ed9904df42e3f81c634['h00de6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f4] =  I0310077d53ae4ed9904df42e3f81c634['h00de8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f5] =  I0310077d53ae4ed9904df42e3f81c634['h00dea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f6] =  I0310077d53ae4ed9904df42e3f81c634['h00dec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f7] =  I0310077d53ae4ed9904df42e3f81c634['h00dee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f8] =  I0310077d53ae4ed9904df42e3f81c634['h00df0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006f9] =  I0310077d53ae4ed9904df42e3f81c634['h00df2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006fa] =  I0310077d53ae4ed9904df42e3f81c634['h00df4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006fb] =  I0310077d53ae4ed9904df42e3f81c634['h00df6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006fc] =  I0310077d53ae4ed9904df42e3f81c634['h00df8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006fd] =  I0310077d53ae4ed9904df42e3f81c634['h00dfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006fe] =  I0310077d53ae4ed9904df42e3f81c634['h00dfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h006ff] =  I0310077d53ae4ed9904df42e3f81c634['h00dfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00700] =  I0310077d53ae4ed9904df42e3f81c634['h00e00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00701] =  I0310077d53ae4ed9904df42e3f81c634['h00e02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00702] =  I0310077d53ae4ed9904df42e3f81c634['h00e04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00703] =  I0310077d53ae4ed9904df42e3f81c634['h00e06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00704] =  I0310077d53ae4ed9904df42e3f81c634['h00e08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00705] =  I0310077d53ae4ed9904df42e3f81c634['h00e0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00706] =  I0310077d53ae4ed9904df42e3f81c634['h00e0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00707] =  I0310077d53ae4ed9904df42e3f81c634['h00e0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00708] =  I0310077d53ae4ed9904df42e3f81c634['h00e10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00709] =  I0310077d53ae4ed9904df42e3f81c634['h00e12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0070a] =  I0310077d53ae4ed9904df42e3f81c634['h00e14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0070b] =  I0310077d53ae4ed9904df42e3f81c634['h00e16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0070c] =  I0310077d53ae4ed9904df42e3f81c634['h00e18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0070d] =  I0310077d53ae4ed9904df42e3f81c634['h00e1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0070e] =  I0310077d53ae4ed9904df42e3f81c634['h00e1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0070f] =  I0310077d53ae4ed9904df42e3f81c634['h00e1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00710] =  I0310077d53ae4ed9904df42e3f81c634['h00e20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00711] =  I0310077d53ae4ed9904df42e3f81c634['h00e22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00712] =  I0310077d53ae4ed9904df42e3f81c634['h00e24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00713] =  I0310077d53ae4ed9904df42e3f81c634['h00e26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00714] =  I0310077d53ae4ed9904df42e3f81c634['h00e28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00715] =  I0310077d53ae4ed9904df42e3f81c634['h00e2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00716] =  I0310077d53ae4ed9904df42e3f81c634['h00e2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00717] =  I0310077d53ae4ed9904df42e3f81c634['h00e2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00718] =  I0310077d53ae4ed9904df42e3f81c634['h00e30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00719] =  I0310077d53ae4ed9904df42e3f81c634['h00e32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0071a] =  I0310077d53ae4ed9904df42e3f81c634['h00e34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0071b] =  I0310077d53ae4ed9904df42e3f81c634['h00e36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0071c] =  I0310077d53ae4ed9904df42e3f81c634['h00e38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0071d] =  I0310077d53ae4ed9904df42e3f81c634['h00e3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0071e] =  I0310077d53ae4ed9904df42e3f81c634['h00e3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0071f] =  I0310077d53ae4ed9904df42e3f81c634['h00e3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00720] =  I0310077d53ae4ed9904df42e3f81c634['h00e40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00721] =  I0310077d53ae4ed9904df42e3f81c634['h00e42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00722] =  I0310077d53ae4ed9904df42e3f81c634['h00e44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00723] =  I0310077d53ae4ed9904df42e3f81c634['h00e46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00724] =  I0310077d53ae4ed9904df42e3f81c634['h00e48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00725] =  I0310077d53ae4ed9904df42e3f81c634['h00e4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00726] =  I0310077d53ae4ed9904df42e3f81c634['h00e4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00727] =  I0310077d53ae4ed9904df42e3f81c634['h00e4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00728] =  I0310077d53ae4ed9904df42e3f81c634['h00e50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00729] =  I0310077d53ae4ed9904df42e3f81c634['h00e52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0072a] =  I0310077d53ae4ed9904df42e3f81c634['h00e54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0072b] =  I0310077d53ae4ed9904df42e3f81c634['h00e56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0072c] =  I0310077d53ae4ed9904df42e3f81c634['h00e58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0072d] =  I0310077d53ae4ed9904df42e3f81c634['h00e5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0072e] =  I0310077d53ae4ed9904df42e3f81c634['h00e5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0072f] =  I0310077d53ae4ed9904df42e3f81c634['h00e5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00730] =  I0310077d53ae4ed9904df42e3f81c634['h00e60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00731] =  I0310077d53ae4ed9904df42e3f81c634['h00e62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00732] =  I0310077d53ae4ed9904df42e3f81c634['h00e64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00733] =  I0310077d53ae4ed9904df42e3f81c634['h00e66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00734] =  I0310077d53ae4ed9904df42e3f81c634['h00e68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00735] =  I0310077d53ae4ed9904df42e3f81c634['h00e6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00736] =  I0310077d53ae4ed9904df42e3f81c634['h00e6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00737] =  I0310077d53ae4ed9904df42e3f81c634['h00e6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00738] =  I0310077d53ae4ed9904df42e3f81c634['h00e70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00739] =  I0310077d53ae4ed9904df42e3f81c634['h00e72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0073a] =  I0310077d53ae4ed9904df42e3f81c634['h00e74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0073b] =  I0310077d53ae4ed9904df42e3f81c634['h00e76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0073c] =  I0310077d53ae4ed9904df42e3f81c634['h00e78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0073d] =  I0310077d53ae4ed9904df42e3f81c634['h00e7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0073e] =  I0310077d53ae4ed9904df42e3f81c634['h00e7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0073f] =  I0310077d53ae4ed9904df42e3f81c634['h00e7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00740] =  I0310077d53ae4ed9904df42e3f81c634['h00e80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00741] =  I0310077d53ae4ed9904df42e3f81c634['h00e82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00742] =  I0310077d53ae4ed9904df42e3f81c634['h00e84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00743] =  I0310077d53ae4ed9904df42e3f81c634['h00e86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00744] =  I0310077d53ae4ed9904df42e3f81c634['h00e88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00745] =  I0310077d53ae4ed9904df42e3f81c634['h00e8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00746] =  I0310077d53ae4ed9904df42e3f81c634['h00e8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00747] =  I0310077d53ae4ed9904df42e3f81c634['h00e8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00748] =  I0310077d53ae4ed9904df42e3f81c634['h00e90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00749] =  I0310077d53ae4ed9904df42e3f81c634['h00e92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0074a] =  I0310077d53ae4ed9904df42e3f81c634['h00e94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0074b] =  I0310077d53ae4ed9904df42e3f81c634['h00e96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0074c] =  I0310077d53ae4ed9904df42e3f81c634['h00e98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0074d] =  I0310077d53ae4ed9904df42e3f81c634['h00e9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0074e] =  I0310077d53ae4ed9904df42e3f81c634['h00e9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0074f] =  I0310077d53ae4ed9904df42e3f81c634['h00e9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00750] =  I0310077d53ae4ed9904df42e3f81c634['h00ea0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00751] =  I0310077d53ae4ed9904df42e3f81c634['h00ea2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00752] =  I0310077d53ae4ed9904df42e3f81c634['h00ea4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00753] =  I0310077d53ae4ed9904df42e3f81c634['h00ea6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00754] =  I0310077d53ae4ed9904df42e3f81c634['h00ea8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00755] =  I0310077d53ae4ed9904df42e3f81c634['h00eaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00756] =  I0310077d53ae4ed9904df42e3f81c634['h00eac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00757] =  I0310077d53ae4ed9904df42e3f81c634['h00eae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00758] =  I0310077d53ae4ed9904df42e3f81c634['h00eb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00759] =  I0310077d53ae4ed9904df42e3f81c634['h00eb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0075a] =  I0310077d53ae4ed9904df42e3f81c634['h00eb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0075b] =  I0310077d53ae4ed9904df42e3f81c634['h00eb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0075c] =  I0310077d53ae4ed9904df42e3f81c634['h00eb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0075d] =  I0310077d53ae4ed9904df42e3f81c634['h00eba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0075e] =  I0310077d53ae4ed9904df42e3f81c634['h00ebc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0075f] =  I0310077d53ae4ed9904df42e3f81c634['h00ebe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00760] =  I0310077d53ae4ed9904df42e3f81c634['h00ec0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00761] =  I0310077d53ae4ed9904df42e3f81c634['h00ec2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00762] =  I0310077d53ae4ed9904df42e3f81c634['h00ec4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00763] =  I0310077d53ae4ed9904df42e3f81c634['h00ec6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00764] =  I0310077d53ae4ed9904df42e3f81c634['h00ec8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00765] =  I0310077d53ae4ed9904df42e3f81c634['h00eca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00766] =  I0310077d53ae4ed9904df42e3f81c634['h00ecc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00767] =  I0310077d53ae4ed9904df42e3f81c634['h00ece] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00768] =  I0310077d53ae4ed9904df42e3f81c634['h00ed0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00769] =  I0310077d53ae4ed9904df42e3f81c634['h00ed2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0076a] =  I0310077d53ae4ed9904df42e3f81c634['h00ed4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0076b] =  I0310077d53ae4ed9904df42e3f81c634['h00ed6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0076c] =  I0310077d53ae4ed9904df42e3f81c634['h00ed8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0076d] =  I0310077d53ae4ed9904df42e3f81c634['h00eda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0076e] =  I0310077d53ae4ed9904df42e3f81c634['h00edc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0076f] =  I0310077d53ae4ed9904df42e3f81c634['h00ede] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00770] =  I0310077d53ae4ed9904df42e3f81c634['h00ee0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00771] =  I0310077d53ae4ed9904df42e3f81c634['h00ee2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00772] =  I0310077d53ae4ed9904df42e3f81c634['h00ee4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00773] =  I0310077d53ae4ed9904df42e3f81c634['h00ee6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00774] =  I0310077d53ae4ed9904df42e3f81c634['h00ee8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00775] =  I0310077d53ae4ed9904df42e3f81c634['h00eea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00776] =  I0310077d53ae4ed9904df42e3f81c634['h00eec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00777] =  I0310077d53ae4ed9904df42e3f81c634['h00eee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00778] =  I0310077d53ae4ed9904df42e3f81c634['h00ef0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00779] =  I0310077d53ae4ed9904df42e3f81c634['h00ef2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0077a] =  I0310077d53ae4ed9904df42e3f81c634['h00ef4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0077b] =  I0310077d53ae4ed9904df42e3f81c634['h00ef6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0077c] =  I0310077d53ae4ed9904df42e3f81c634['h00ef8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0077d] =  I0310077d53ae4ed9904df42e3f81c634['h00efa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0077e] =  I0310077d53ae4ed9904df42e3f81c634['h00efc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0077f] =  I0310077d53ae4ed9904df42e3f81c634['h00efe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00780] =  I0310077d53ae4ed9904df42e3f81c634['h00f00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00781] =  I0310077d53ae4ed9904df42e3f81c634['h00f02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00782] =  I0310077d53ae4ed9904df42e3f81c634['h00f04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00783] =  I0310077d53ae4ed9904df42e3f81c634['h00f06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00784] =  I0310077d53ae4ed9904df42e3f81c634['h00f08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00785] =  I0310077d53ae4ed9904df42e3f81c634['h00f0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00786] =  I0310077d53ae4ed9904df42e3f81c634['h00f0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00787] =  I0310077d53ae4ed9904df42e3f81c634['h00f0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00788] =  I0310077d53ae4ed9904df42e3f81c634['h00f10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00789] =  I0310077d53ae4ed9904df42e3f81c634['h00f12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0078a] =  I0310077d53ae4ed9904df42e3f81c634['h00f14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0078b] =  I0310077d53ae4ed9904df42e3f81c634['h00f16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0078c] =  I0310077d53ae4ed9904df42e3f81c634['h00f18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0078d] =  I0310077d53ae4ed9904df42e3f81c634['h00f1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0078e] =  I0310077d53ae4ed9904df42e3f81c634['h00f1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0078f] =  I0310077d53ae4ed9904df42e3f81c634['h00f1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00790] =  I0310077d53ae4ed9904df42e3f81c634['h00f20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00791] =  I0310077d53ae4ed9904df42e3f81c634['h00f22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00792] =  I0310077d53ae4ed9904df42e3f81c634['h00f24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00793] =  I0310077d53ae4ed9904df42e3f81c634['h00f26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00794] =  I0310077d53ae4ed9904df42e3f81c634['h00f28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00795] =  I0310077d53ae4ed9904df42e3f81c634['h00f2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00796] =  I0310077d53ae4ed9904df42e3f81c634['h00f2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00797] =  I0310077d53ae4ed9904df42e3f81c634['h00f2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00798] =  I0310077d53ae4ed9904df42e3f81c634['h00f30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00799] =  I0310077d53ae4ed9904df42e3f81c634['h00f32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0079a] =  I0310077d53ae4ed9904df42e3f81c634['h00f34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0079b] =  I0310077d53ae4ed9904df42e3f81c634['h00f36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0079c] =  I0310077d53ae4ed9904df42e3f81c634['h00f38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0079d] =  I0310077d53ae4ed9904df42e3f81c634['h00f3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0079e] =  I0310077d53ae4ed9904df42e3f81c634['h00f3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0079f] =  I0310077d53ae4ed9904df42e3f81c634['h00f3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a0] =  I0310077d53ae4ed9904df42e3f81c634['h00f40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a1] =  I0310077d53ae4ed9904df42e3f81c634['h00f42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a2] =  I0310077d53ae4ed9904df42e3f81c634['h00f44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a3] =  I0310077d53ae4ed9904df42e3f81c634['h00f46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a4] =  I0310077d53ae4ed9904df42e3f81c634['h00f48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a5] =  I0310077d53ae4ed9904df42e3f81c634['h00f4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a6] =  I0310077d53ae4ed9904df42e3f81c634['h00f4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a7] =  I0310077d53ae4ed9904df42e3f81c634['h00f4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a8] =  I0310077d53ae4ed9904df42e3f81c634['h00f50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007a9] =  I0310077d53ae4ed9904df42e3f81c634['h00f52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007aa] =  I0310077d53ae4ed9904df42e3f81c634['h00f54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ab] =  I0310077d53ae4ed9904df42e3f81c634['h00f56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ac] =  I0310077d53ae4ed9904df42e3f81c634['h00f58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ad] =  I0310077d53ae4ed9904df42e3f81c634['h00f5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ae] =  I0310077d53ae4ed9904df42e3f81c634['h00f5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007af] =  I0310077d53ae4ed9904df42e3f81c634['h00f5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b0] =  I0310077d53ae4ed9904df42e3f81c634['h00f60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b1] =  I0310077d53ae4ed9904df42e3f81c634['h00f62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b2] =  I0310077d53ae4ed9904df42e3f81c634['h00f64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b3] =  I0310077d53ae4ed9904df42e3f81c634['h00f66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b4] =  I0310077d53ae4ed9904df42e3f81c634['h00f68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b5] =  I0310077d53ae4ed9904df42e3f81c634['h00f6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b6] =  I0310077d53ae4ed9904df42e3f81c634['h00f6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b7] =  I0310077d53ae4ed9904df42e3f81c634['h00f6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b8] =  I0310077d53ae4ed9904df42e3f81c634['h00f70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007b9] =  I0310077d53ae4ed9904df42e3f81c634['h00f72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ba] =  I0310077d53ae4ed9904df42e3f81c634['h00f74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007bb] =  I0310077d53ae4ed9904df42e3f81c634['h00f76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007bc] =  I0310077d53ae4ed9904df42e3f81c634['h00f78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007bd] =  I0310077d53ae4ed9904df42e3f81c634['h00f7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007be] =  I0310077d53ae4ed9904df42e3f81c634['h00f7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007bf] =  I0310077d53ae4ed9904df42e3f81c634['h00f7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c0] =  I0310077d53ae4ed9904df42e3f81c634['h00f80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c1] =  I0310077d53ae4ed9904df42e3f81c634['h00f82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c2] =  I0310077d53ae4ed9904df42e3f81c634['h00f84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c3] =  I0310077d53ae4ed9904df42e3f81c634['h00f86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c4] =  I0310077d53ae4ed9904df42e3f81c634['h00f88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c5] =  I0310077d53ae4ed9904df42e3f81c634['h00f8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c6] =  I0310077d53ae4ed9904df42e3f81c634['h00f8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c7] =  I0310077d53ae4ed9904df42e3f81c634['h00f8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c8] =  I0310077d53ae4ed9904df42e3f81c634['h00f90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007c9] =  I0310077d53ae4ed9904df42e3f81c634['h00f92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ca] =  I0310077d53ae4ed9904df42e3f81c634['h00f94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007cb] =  I0310077d53ae4ed9904df42e3f81c634['h00f96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007cc] =  I0310077d53ae4ed9904df42e3f81c634['h00f98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007cd] =  I0310077d53ae4ed9904df42e3f81c634['h00f9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ce] =  I0310077d53ae4ed9904df42e3f81c634['h00f9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007cf] =  I0310077d53ae4ed9904df42e3f81c634['h00f9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d0] =  I0310077d53ae4ed9904df42e3f81c634['h00fa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d1] =  I0310077d53ae4ed9904df42e3f81c634['h00fa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d2] =  I0310077d53ae4ed9904df42e3f81c634['h00fa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d3] =  I0310077d53ae4ed9904df42e3f81c634['h00fa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d4] =  I0310077d53ae4ed9904df42e3f81c634['h00fa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d5] =  I0310077d53ae4ed9904df42e3f81c634['h00faa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d6] =  I0310077d53ae4ed9904df42e3f81c634['h00fac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d7] =  I0310077d53ae4ed9904df42e3f81c634['h00fae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d8] =  I0310077d53ae4ed9904df42e3f81c634['h00fb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007d9] =  I0310077d53ae4ed9904df42e3f81c634['h00fb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007da] =  I0310077d53ae4ed9904df42e3f81c634['h00fb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007db] =  I0310077d53ae4ed9904df42e3f81c634['h00fb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007dc] =  I0310077d53ae4ed9904df42e3f81c634['h00fb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007dd] =  I0310077d53ae4ed9904df42e3f81c634['h00fba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007de] =  I0310077d53ae4ed9904df42e3f81c634['h00fbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007df] =  I0310077d53ae4ed9904df42e3f81c634['h00fbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e0] =  I0310077d53ae4ed9904df42e3f81c634['h00fc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e1] =  I0310077d53ae4ed9904df42e3f81c634['h00fc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e2] =  I0310077d53ae4ed9904df42e3f81c634['h00fc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e3] =  I0310077d53ae4ed9904df42e3f81c634['h00fc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e4] =  I0310077d53ae4ed9904df42e3f81c634['h00fc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e5] =  I0310077d53ae4ed9904df42e3f81c634['h00fca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e6] =  I0310077d53ae4ed9904df42e3f81c634['h00fcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e7] =  I0310077d53ae4ed9904df42e3f81c634['h00fce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e8] =  I0310077d53ae4ed9904df42e3f81c634['h00fd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007e9] =  I0310077d53ae4ed9904df42e3f81c634['h00fd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ea] =  I0310077d53ae4ed9904df42e3f81c634['h00fd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007eb] =  I0310077d53ae4ed9904df42e3f81c634['h00fd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ec] =  I0310077d53ae4ed9904df42e3f81c634['h00fd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ed] =  I0310077d53ae4ed9904df42e3f81c634['h00fda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ee] =  I0310077d53ae4ed9904df42e3f81c634['h00fdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ef] =  I0310077d53ae4ed9904df42e3f81c634['h00fde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f0] =  I0310077d53ae4ed9904df42e3f81c634['h00fe0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f1] =  I0310077d53ae4ed9904df42e3f81c634['h00fe2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f2] =  I0310077d53ae4ed9904df42e3f81c634['h00fe4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f3] =  I0310077d53ae4ed9904df42e3f81c634['h00fe6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f4] =  I0310077d53ae4ed9904df42e3f81c634['h00fe8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f5] =  I0310077d53ae4ed9904df42e3f81c634['h00fea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f6] =  I0310077d53ae4ed9904df42e3f81c634['h00fec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f7] =  I0310077d53ae4ed9904df42e3f81c634['h00fee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f8] =  I0310077d53ae4ed9904df42e3f81c634['h00ff0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007f9] =  I0310077d53ae4ed9904df42e3f81c634['h00ff2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007fa] =  I0310077d53ae4ed9904df42e3f81c634['h00ff4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007fb] =  I0310077d53ae4ed9904df42e3f81c634['h00ff6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007fc] =  I0310077d53ae4ed9904df42e3f81c634['h00ff8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007fd] =  I0310077d53ae4ed9904df42e3f81c634['h00ffa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007fe] =  I0310077d53ae4ed9904df42e3f81c634['h00ffc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h007ff] =  I0310077d53ae4ed9904df42e3f81c634['h00ffe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00800] =  I0310077d53ae4ed9904df42e3f81c634['h01000] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00801] =  I0310077d53ae4ed9904df42e3f81c634['h01002] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00802] =  I0310077d53ae4ed9904df42e3f81c634['h01004] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00803] =  I0310077d53ae4ed9904df42e3f81c634['h01006] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00804] =  I0310077d53ae4ed9904df42e3f81c634['h01008] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00805] =  I0310077d53ae4ed9904df42e3f81c634['h0100a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00806] =  I0310077d53ae4ed9904df42e3f81c634['h0100c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00807] =  I0310077d53ae4ed9904df42e3f81c634['h0100e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00808] =  I0310077d53ae4ed9904df42e3f81c634['h01010] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00809] =  I0310077d53ae4ed9904df42e3f81c634['h01012] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0080a] =  I0310077d53ae4ed9904df42e3f81c634['h01014] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0080b] =  I0310077d53ae4ed9904df42e3f81c634['h01016] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0080c] =  I0310077d53ae4ed9904df42e3f81c634['h01018] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0080d] =  I0310077d53ae4ed9904df42e3f81c634['h0101a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0080e] =  I0310077d53ae4ed9904df42e3f81c634['h0101c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0080f] =  I0310077d53ae4ed9904df42e3f81c634['h0101e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00810] =  I0310077d53ae4ed9904df42e3f81c634['h01020] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00811] =  I0310077d53ae4ed9904df42e3f81c634['h01022] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00812] =  I0310077d53ae4ed9904df42e3f81c634['h01024] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00813] =  I0310077d53ae4ed9904df42e3f81c634['h01026] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00814] =  I0310077d53ae4ed9904df42e3f81c634['h01028] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00815] =  I0310077d53ae4ed9904df42e3f81c634['h0102a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00816] =  I0310077d53ae4ed9904df42e3f81c634['h0102c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00817] =  I0310077d53ae4ed9904df42e3f81c634['h0102e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00818] =  I0310077d53ae4ed9904df42e3f81c634['h01030] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00819] =  I0310077d53ae4ed9904df42e3f81c634['h01032] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0081a] =  I0310077d53ae4ed9904df42e3f81c634['h01034] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0081b] =  I0310077d53ae4ed9904df42e3f81c634['h01036] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0081c] =  I0310077d53ae4ed9904df42e3f81c634['h01038] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0081d] =  I0310077d53ae4ed9904df42e3f81c634['h0103a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0081e] =  I0310077d53ae4ed9904df42e3f81c634['h0103c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0081f] =  I0310077d53ae4ed9904df42e3f81c634['h0103e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00820] =  I0310077d53ae4ed9904df42e3f81c634['h01040] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00821] =  I0310077d53ae4ed9904df42e3f81c634['h01042] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00822] =  I0310077d53ae4ed9904df42e3f81c634['h01044] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00823] =  I0310077d53ae4ed9904df42e3f81c634['h01046] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00824] =  I0310077d53ae4ed9904df42e3f81c634['h01048] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00825] =  I0310077d53ae4ed9904df42e3f81c634['h0104a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00826] =  I0310077d53ae4ed9904df42e3f81c634['h0104c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00827] =  I0310077d53ae4ed9904df42e3f81c634['h0104e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00828] =  I0310077d53ae4ed9904df42e3f81c634['h01050] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00829] =  I0310077d53ae4ed9904df42e3f81c634['h01052] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0082a] =  I0310077d53ae4ed9904df42e3f81c634['h01054] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0082b] =  I0310077d53ae4ed9904df42e3f81c634['h01056] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0082c] =  I0310077d53ae4ed9904df42e3f81c634['h01058] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0082d] =  I0310077d53ae4ed9904df42e3f81c634['h0105a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0082e] =  I0310077d53ae4ed9904df42e3f81c634['h0105c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0082f] =  I0310077d53ae4ed9904df42e3f81c634['h0105e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00830] =  I0310077d53ae4ed9904df42e3f81c634['h01060] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00831] =  I0310077d53ae4ed9904df42e3f81c634['h01062] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00832] =  I0310077d53ae4ed9904df42e3f81c634['h01064] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00833] =  I0310077d53ae4ed9904df42e3f81c634['h01066] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00834] =  I0310077d53ae4ed9904df42e3f81c634['h01068] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00835] =  I0310077d53ae4ed9904df42e3f81c634['h0106a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00836] =  I0310077d53ae4ed9904df42e3f81c634['h0106c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00837] =  I0310077d53ae4ed9904df42e3f81c634['h0106e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00838] =  I0310077d53ae4ed9904df42e3f81c634['h01070] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00839] =  I0310077d53ae4ed9904df42e3f81c634['h01072] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0083a] =  I0310077d53ae4ed9904df42e3f81c634['h01074] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0083b] =  I0310077d53ae4ed9904df42e3f81c634['h01076] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0083c] =  I0310077d53ae4ed9904df42e3f81c634['h01078] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0083d] =  I0310077d53ae4ed9904df42e3f81c634['h0107a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0083e] =  I0310077d53ae4ed9904df42e3f81c634['h0107c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0083f] =  I0310077d53ae4ed9904df42e3f81c634['h0107e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00840] =  I0310077d53ae4ed9904df42e3f81c634['h01080] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00841] =  I0310077d53ae4ed9904df42e3f81c634['h01082] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00842] =  I0310077d53ae4ed9904df42e3f81c634['h01084] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00843] =  I0310077d53ae4ed9904df42e3f81c634['h01086] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00844] =  I0310077d53ae4ed9904df42e3f81c634['h01088] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00845] =  I0310077d53ae4ed9904df42e3f81c634['h0108a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00846] =  I0310077d53ae4ed9904df42e3f81c634['h0108c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00847] =  I0310077d53ae4ed9904df42e3f81c634['h0108e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00848] =  I0310077d53ae4ed9904df42e3f81c634['h01090] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00849] =  I0310077d53ae4ed9904df42e3f81c634['h01092] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0084a] =  I0310077d53ae4ed9904df42e3f81c634['h01094] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0084b] =  I0310077d53ae4ed9904df42e3f81c634['h01096] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0084c] =  I0310077d53ae4ed9904df42e3f81c634['h01098] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0084d] =  I0310077d53ae4ed9904df42e3f81c634['h0109a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0084e] =  I0310077d53ae4ed9904df42e3f81c634['h0109c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0084f] =  I0310077d53ae4ed9904df42e3f81c634['h0109e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00850] =  I0310077d53ae4ed9904df42e3f81c634['h010a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00851] =  I0310077d53ae4ed9904df42e3f81c634['h010a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00852] =  I0310077d53ae4ed9904df42e3f81c634['h010a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00853] =  I0310077d53ae4ed9904df42e3f81c634['h010a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00854] =  I0310077d53ae4ed9904df42e3f81c634['h010a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00855] =  I0310077d53ae4ed9904df42e3f81c634['h010aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00856] =  I0310077d53ae4ed9904df42e3f81c634['h010ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00857] =  I0310077d53ae4ed9904df42e3f81c634['h010ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00858] =  I0310077d53ae4ed9904df42e3f81c634['h010b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00859] =  I0310077d53ae4ed9904df42e3f81c634['h010b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0085a] =  I0310077d53ae4ed9904df42e3f81c634['h010b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0085b] =  I0310077d53ae4ed9904df42e3f81c634['h010b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0085c] =  I0310077d53ae4ed9904df42e3f81c634['h010b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0085d] =  I0310077d53ae4ed9904df42e3f81c634['h010ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0085e] =  I0310077d53ae4ed9904df42e3f81c634['h010bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0085f] =  I0310077d53ae4ed9904df42e3f81c634['h010be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00860] =  I0310077d53ae4ed9904df42e3f81c634['h010c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00861] =  I0310077d53ae4ed9904df42e3f81c634['h010c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00862] =  I0310077d53ae4ed9904df42e3f81c634['h010c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00863] =  I0310077d53ae4ed9904df42e3f81c634['h010c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00864] =  I0310077d53ae4ed9904df42e3f81c634['h010c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00865] =  I0310077d53ae4ed9904df42e3f81c634['h010ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00866] =  I0310077d53ae4ed9904df42e3f81c634['h010cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00867] =  I0310077d53ae4ed9904df42e3f81c634['h010ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00868] =  I0310077d53ae4ed9904df42e3f81c634['h010d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00869] =  I0310077d53ae4ed9904df42e3f81c634['h010d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0086a] =  I0310077d53ae4ed9904df42e3f81c634['h010d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0086b] =  I0310077d53ae4ed9904df42e3f81c634['h010d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0086c] =  I0310077d53ae4ed9904df42e3f81c634['h010d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0086d] =  I0310077d53ae4ed9904df42e3f81c634['h010da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0086e] =  I0310077d53ae4ed9904df42e3f81c634['h010dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0086f] =  I0310077d53ae4ed9904df42e3f81c634['h010de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00870] =  I0310077d53ae4ed9904df42e3f81c634['h010e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00871] =  I0310077d53ae4ed9904df42e3f81c634['h010e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00872] =  I0310077d53ae4ed9904df42e3f81c634['h010e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00873] =  I0310077d53ae4ed9904df42e3f81c634['h010e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00874] =  I0310077d53ae4ed9904df42e3f81c634['h010e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00875] =  I0310077d53ae4ed9904df42e3f81c634['h010ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00876] =  I0310077d53ae4ed9904df42e3f81c634['h010ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00877] =  I0310077d53ae4ed9904df42e3f81c634['h010ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00878] =  I0310077d53ae4ed9904df42e3f81c634['h010f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00879] =  I0310077d53ae4ed9904df42e3f81c634['h010f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0087a] =  I0310077d53ae4ed9904df42e3f81c634['h010f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0087b] =  I0310077d53ae4ed9904df42e3f81c634['h010f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0087c] =  I0310077d53ae4ed9904df42e3f81c634['h010f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0087d] =  I0310077d53ae4ed9904df42e3f81c634['h010fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0087e] =  I0310077d53ae4ed9904df42e3f81c634['h010fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0087f] =  I0310077d53ae4ed9904df42e3f81c634['h010fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00880] =  I0310077d53ae4ed9904df42e3f81c634['h01100] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00881] =  I0310077d53ae4ed9904df42e3f81c634['h01102] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00882] =  I0310077d53ae4ed9904df42e3f81c634['h01104] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00883] =  I0310077d53ae4ed9904df42e3f81c634['h01106] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00884] =  I0310077d53ae4ed9904df42e3f81c634['h01108] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00885] =  I0310077d53ae4ed9904df42e3f81c634['h0110a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00886] =  I0310077d53ae4ed9904df42e3f81c634['h0110c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00887] =  I0310077d53ae4ed9904df42e3f81c634['h0110e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00888] =  I0310077d53ae4ed9904df42e3f81c634['h01110] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00889] =  I0310077d53ae4ed9904df42e3f81c634['h01112] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0088a] =  I0310077d53ae4ed9904df42e3f81c634['h01114] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0088b] =  I0310077d53ae4ed9904df42e3f81c634['h01116] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0088c] =  I0310077d53ae4ed9904df42e3f81c634['h01118] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0088d] =  I0310077d53ae4ed9904df42e3f81c634['h0111a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0088e] =  I0310077d53ae4ed9904df42e3f81c634['h0111c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0088f] =  I0310077d53ae4ed9904df42e3f81c634['h0111e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00890] =  I0310077d53ae4ed9904df42e3f81c634['h01120] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00891] =  I0310077d53ae4ed9904df42e3f81c634['h01122] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00892] =  I0310077d53ae4ed9904df42e3f81c634['h01124] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00893] =  I0310077d53ae4ed9904df42e3f81c634['h01126] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00894] =  I0310077d53ae4ed9904df42e3f81c634['h01128] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00895] =  I0310077d53ae4ed9904df42e3f81c634['h0112a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00896] =  I0310077d53ae4ed9904df42e3f81c634['h0112c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00897] =  I0310077d53ae4ed9904df42e3f81c634['h0112e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00898] =  I0310077d53ae4ed9904df42e3f81c634['h01130] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00899] =  I0310077d53ae4ed9904df42e3f81c634['h01132] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0089a] =  I0310077d53ae4ed9904df42e3f81c634['h01134] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0089b] =  I0310077d53ae4ed9904df42e3f81c634['h01136] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0089c] =  I0310077d53ae4ed9904df42e3f81c634['h01138] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0089d] =  I0310077d53ae4ed9904df42e3f81c634['h0113a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0089e] =  I0310077d53ae4ed9904df42e3f81c634['h0113c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0089f] =  I0310077d53ae4ed9904df42e3f81c634['h0113e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a0] =  I0310077d53ae4ed9904df42e3f81c634['h01140] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a1] =  I0310077d53ae4ed9904df42e3f81c634['h01142] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a2] =  I0310077d53ae4ed9904df42e3f81c634['h01144] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a3] =  I0310077d53ae4ed9904df42e3f81c634['h01146] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a4] =  I0310077d53ae4ed9904df42e3f81c634['h01148] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a5] =  I0310077d53ae4ed9904df42e3f81c634['h0114a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a6] =  I0310077d53ae4ed9904df42e3f81c634['h0114c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a7] =  I0310077d53ae4ed9904df42e3f81c634['h0114e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a8] =  I0310077d53ae4ed9904df42e3f81c634['h01150] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008a9] =  I0310077d53ae4ed9904df42e3f81c634['h01152] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008aa] =  I0310077d53ae4ed9904df42e3f81c634['h01154] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ab] =  I0310077d53ae4ed9904df42e3f81c634['h01156] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ac] =  I0310077d53ae4ed9904df42e3f81c634['h01158] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ad] =  I0310077d53ae4ed9904df42e3f81c634['h0115a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ae] =  I0310077d53ae4ed9904df42e3f81c634['h0115c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008af] =  I0310077d53ae4ed9904df42e3f81c634['h0115e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b0] =  I0310077d53ae4ed9904df42e3f81c634['h01160] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b1] =  I0310077d53ae4ed9904df42e3f81c634['h01162] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b2] =  I0310077d53ae4ed9904df42e3f81c634['h01164] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b3] =  I0310077d53ae4ed9904df42e3f81c634['h01166] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b4] =  I0310077d53ae4ed9904df42e3f81c634['h01168] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b5] =  I0310077d53ae4ed9904df42e3f81c634['h0116a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b6] =  I0310077d53ae4ed9904df42e3f81c634['h0116c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b7] =  I0310077d53ae4ed9904df42e3f81c634['h0116e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b8] =  I0310077d53ae4ed9904df42e3f81c634['h01170] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008b9] =  I0310077d53ae4ed9904df42e3f81c634['h01172] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ba] =  I0310077d53ae4ed9904df42e3f81c634['h01174] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008bb] =  I0310077d53ae4ed9904df42e3f81c634['h01176] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008bc] =  I0310077d53ae4ed9904df42e3f81c634['h01178] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008bd] =  I0310077d53ae4ed9904df42e3f81c634['h0117a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008be] =  I0310077d53ae4ed9904df42e3f81c634['h0117c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008bf] =  I0310077d53ae4ed9904df42e3f81c634['h0117e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c0] =  I0310077d53ae4ed9904df42e3f81c634['h01180] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c1] =  I0310077d53ae4ed9904df42e3f81c634['h01182] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c2] =  I0310077d53ae4ed9904df42e3f81c634['h01184] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c3] =  I0310077d53ae4ed9904df42e3f81c634['h01186] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c4] =  I0310077d53ae4ed9904df42e3f81c634['h01188] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c5] =  I0310077d53ae4ed9904df42e3f81c634['h0118a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c6] =  I0310077d53ae4ed9904df42e3f81c634['h0118c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c7] =  I0310077d53ae4ed9904df42e3f81c634['h0118e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c8] =  I0310077d53ae4ed9904df42e3f81c634['h01190] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008c9] =  I0310077d53ae4ed9904df42e3f81c634['h01192] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ca] =  I0310077d53ae4ed9904df42e3f81c634['h01194] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008cb] =  I0310077d53ae4ed9904df42e3f81c634['h01196] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008cc] =  I0310077d53ae4ed9904df42e3f81c634['h01198] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008cd] =  I0310077d53ae4ed9904df42e3f81c634['h0119a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ce] =  I0310077d53ae4ed9904df42e3f81c634['h0119c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008cf] =  I0310077d53ae4ed9904df42e3f81c634['h0119e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d0] =  I0310077d53ae4ed9904df42e3f81c634['h011a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d1] =  I0310077d53ae4ed9904df42e3f81c634['h011a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d2] =  I0310077d53ae4ed9904df42e3f81c634['h011a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d3] =  I0310077d53ae4ed9904df42e3f81c634['h011a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d4] =  I0310077d53ae4ed9904df42e3f81c634['h011a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d5] =  I0310077d53ae4ed9904df42e3f81c634['h011aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d6] =  I0310077d53ae4ed9904df42e3f81c634['h011ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d7] =  I0310077d53ae4ed9904df42e3f81c634['h011ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d8] =  I0310077d53ae4ed9904df42e3f81c634['h011b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008d9] =  I0310077d53ae4ed9904df42e3f81c634['h011b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008da] =  I0310077d53ae4ed9904df42e3f81c634['h011b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008db] =  I0310077d53ae4ed9904df42e3f81c634['h011b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008dc] =  I0310077d53ae4ed9904df42e3f81c634['h011b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008dd] =  I0310077d53ae4ed9904df42e3f81c634['h011ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008de] =  I0310077d53ae4ed9904df42e3f81c634['h011bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008df] =  I0310077d53ae4ed9904df42e3f81c634['h011be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e0] =  I0310077d53ae4ed9904df42e3f81c634['h011c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e1] =  I0310077d53ae4ed9904df42e3f81c634['h011c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e2] =  I0310077d53ae4ed9904df42e3f81c634['h011c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e3] =  I0310077d53ae4ed9904df42e3f81c634['h011c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e4] =  I0310077d53ae4ed9904df42e3f81c634['h011c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e5] =  I0310077d53ae4ed9904df42e3f81c634['h011ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e6] =  I0310077d53ae4ed9904df42e3f81c634['h011cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e7] =  I0310077d53ae4ed9904df42e3f81c634['h011ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e8] =  I0310077d53ae4ed9904df42e3f81c634['h011d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008e9] =  I0310077d53ae4ed9904df42e3f81c634['h011d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ea] =  I0310077d53ae4ed9904df42e3f81c634['h011d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008eb] =  I0310077d53ae4ed9904df42e3f81c634['h011d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ec] =  I0310077d53ae4ed9904df42e3f81c634['h011d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ed] =  I0310077d53ae4ed9904df42e3f81c634['h011da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ee] =  I0310077d53ae4ed9904df42e3f81c634['h011dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ef] =  I0310077d53ae4ed9904df42e3f81c634['h011de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f0] =  I0310077d53ae4ed9904df42e3f81c634['h011e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f1] =  I0310077d53ae4ed9904df42e3f81c634['h011e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f2] =  I0310077d53ae4ed9904df42e3f81c634['h011e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f3] =  I0310077d53ae4ed9904df42e3f81c634['h011e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f4] =  I0310077d53ae4ed9904df42e3f81c634['h011e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f5] =  I0310077d53ae4ed9904df42e3f81c634['h011ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f6] =  I0310077d53ae4ed9904df42e3f81c634['h011ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f7] =  I0310077d53ae4ed9904df42e3f81c634['h011ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f8] =  I0310077d53ae4ed9904df42e3f81c634['h011f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008f9] =  I0310077d53ae4ed9904df42e3f81c634['h011f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008fa] =  I0310077d53ae4ed9904df42e3f81c634['h011f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008fb] =  I0310077d53ae4ed9904df42e3f81c634['h011f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008fc] =  I0310077d53ae4ed9904df42e3f81c634['h011f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008fd] =  I0310077d53ae4ed9904df42e3f81c634['h011fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008fe] =  I0310077d53ae4ed9904df42e3f81c634['h011fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h008ff] =  I0310077d53ae4ed9904df42e3f81c634['h011fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00900] =  I0310077d53ae4ed9904df42e3f81c634['h01200] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00901] =  I0310077d53ae4ed9904df42e3f81c634['h01202] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00902] =  I0310077d53ae4ed9904df42e3f81c634['h01204] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00903] =  I0310077d53ae4ed9904df42e3f81c634['h01206] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00904] =  I0310077d53ae4ed9904df42e3f81c634['h01208] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00905] =  I0310077d53ae4ed9904df42e3f81c634['h0120a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00906] =  I0310077d53ae4ed9904df42e3f81c634['h0120c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00907] =  I0310077d53ae4ed9904df42e3f81c634['h0120e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00908] =  I0310077d53ae4ed9904df42e3f81c634['h01210] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00909] =  I0310077d53ae4ed9904df42e3f81c634['h01212] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0090a] =  I0310077d53ae4ed9904df42e3f81c634['h01214] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0090b] =  I0310077d53ae4ed9904df42e3f81c634['h01216] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0090c] =  I0310077d53ae4ed9904df42e3f81c634['h01218] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0090d] =  I0310077d53ae4ed9904df42e3f81c634['h0121a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0090e] =  I0310077d53ae4ed9904df42e3f81c634['h0121c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0090f] =  I0310077d53ae4ed9904df42e3f81c634['h0121e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00910] =  I0310077d53ae4ed9904df42e3f81c634['h01220] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00911] =  I0310077d53ae4ed9904df42e3f81c634['h01222] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00912] =  I0310077d53ae4ed9904df42e3f81c634['h01224] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00913] =  I0310077d53ae4ed9904df42e3f81c634['h01226] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00914] =  I0310077d53ae4ed9904df42e3f81c634['h01228] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00915] =  I0310077d53ae4ed9904df42e3f81c634['h0122a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00916] =  I0310077d53ae4ed9904df42e3f81c634['h0122c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00917] =  I0310077d53ae4ed9904df42e3f81c634['h0122e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00918] =  I0310077d53ae4ed9904df42e3f81c634['h01230] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00919] =  I0310077d53ae4ed9904df42e3f81c634['h01232] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0091a] =  I0310077d53ae4ed9904df42e3f81c634['h01234] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0091b] =  I0310077d53ae4ed9904df42e3f81c634['h01236] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0091c] =  I0310077d53ae4ed9904df42e3f81c634['h01238] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0091d] =  I0310077d53ae4ed9904df42e3f81c634['h0123a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0091e] =  I0310077d53ae4ed9904df42e3f81c634['h0123c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0091f] =  I0310077d53ae4ed9904df42e3f81c634['h0123e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00920] =  I0310077d53ae4ed9904df42e3f81c634['h01240] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00921] =  I0310077d53ae4ed9904df42e3f81c634['h01242] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00922] =  I0310077d53ae4ed9904df42e3f81c634['h01244] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00923] =  I0310077d53ae4ed9904df42e3f81c634['h01246] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00924] =  I0310077d53ae4ed9904df42e3f81c634['h01248] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00925] =  I0310077d53ae4ed9904df42e3f81c634['h0124a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00926] =  I0310077d53ae4ed9904df42e3f81c634['h0124c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00927] =  I0310077d53ae4ed9904df42e3f81c634['h0124e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00928] =  I0310077d53ae4ed9904df42e3f81c634['h01250] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00929] =  I0310077d53ae4ed9904df42e3f81c634['h01252] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0092a] =  I0310077d53ae4ed9904df42e3f81c634['h01254] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0092b] =  I0310077d53ae4ed9904df42e3f81c634['h01256] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0092c] =  I0310077d53ae4ed9904df42e3f81c634['h01258] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0092d] =  I0310077d53ae4ed9904df42e3f81c634['h0125a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0092e] =  I0310077d53ae4ed9904df42e3f81c634['h0125c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0092f] =  I0310077d53ae4ed9904df42e3f81c634['h0125e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00930] =  I0310077d53ae4ed9904df42e3f81c634['h01260] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00931] =  I0310077d53ae4ed9904df42e3f81c634['h01262] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00932] =  I0310077d53ae4ed9904df42e3f81c634['h01264] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00933] =  I0310077d53ae4ed9904df42e3f81c634['h01266] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00934] =  I0310077d53ae4ed9904df42e3f81c634['h01268] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00935] =  I0310077d53ae4ed9904df42e3f81c634['h0126a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00936] =  I0310077d53ae4ed9904df42e3f81c634['h0126c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00937] =  I0310077d53ae4ed9904df42e3f81c634['h0126e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00938] =  I0310077d53ae4ed9904df42e3f81c634['h01270] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00939] =  I0310077d53ae4ed9904df42e3f81c634['h01272] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0093a] =  I0310077d53ae4ed9904df42e3f81c634['h01274] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0093b] =  I0310077d53ae4ed9904df42e3f81c634['h01276] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0093c] =  I0310077d53ae4ed9904df42e3f81c634['h01278] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0093d] =  I0310077d53ae4ed9904df42e3f81c634['h0127a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0093e] =  I0310077d53ae4ed9904df42e3f81c634['h0127c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0093f] =  I0310077d53ae4ed9904df42e3f81c634['h0127e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00940] =  I0310077d53ae4ed9904df42e3f81c634['h01280] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00941] =  I0310077d53ae4ed9904df42e3f81c634['h01282] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00942] =  I0310077d53ae4ed9904df42e3f81c634['h01284] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00943] =  I0310077d53ae4ed9904df42e3f81c634['h01286] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00944] =  I0310077d53ae4ed9904df42e3f81c634['h01288] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00945] =  I0310077d53ae4ed9904df42e3f81c634['h0128a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00946] =  I0310077d53ae4ed9904df42e3f81c634['h0128c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00947] =  I0310077d53ae4ed9904df42e3f81c634['h0128e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00948] =  I0310077d53ae4ed9904df42e3f81c634['h01290] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00949] =  I0310077d53ae4ed9904df42e3f81c634['h01292] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0094a] =  I0310077d53ae4ed9904df42e3f81c634['h01294] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0094b] =  I0310077d53ae4ed9904df42e3f81c634['h01296] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0094c] =  I0310077d53ae4ed9904df42e3f81c634['h01298] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0094d] =  I0310077d53ae4ed9904df42e3f81c634['h0129a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0094e] =  I0310077d53ae4ed9904df42e3f81c634['h0129c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0094f] =  I0310077d53ae4ed9904df42e3f81c634['h0129e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00950] =  I0310077d53ae4ed9904df42e3f81c634['h012a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00951] =  I0310077d53ae4ed9904df42e3f81c634['h012a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00952] =  I0310077d53ae4ed9904df42e3f81c634['h012a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00953] =  I0310077d53ae4ed9904df42e3f81c634['h012a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00954] =  I0310077d53ae4ed9904df42e3f81c634['h012a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00955] =  I0310077d53ae4ed9904df42e3f81c634['h012aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00956] =  I0310077d53ae4ed9904df42e3f81c634['h012ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00957] =  I0310077d53ae4ed9904df42e3f81c634['h012ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00958] =  I0310077d53ae4ed9904df42e3f81c634['h012b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00959] =  I0310077d53ae4ed9904df42e3f81c634['h012b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0095a] =  I0310077d53ae4ed9904df42e3f81c634['h012b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0095b] =  I0310077d53ae4ed9904df42e3f81c634['h012b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0095c] =  I0310077d53ae4ed9904df42e3f81c634['h012b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0095d] =  I0310077d53ae4ed9904df42e3f81c634['h012ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0095e] =  I0310077d53ae4ed9904df42e3f81c634['h012bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0095f] =  I0310077d53ae4ed9904df42e3f81c634['h012be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00960] =  I0310077d53ae4ed9904df42e3f81c634['h012c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00961] =  I0310077d53ae4ed9904df42e3f81c634['h012c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00962] =  I0310077d53ae4ed9904df42e3f81c634['h012c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00963] =  I0310077d53ae4ed9904df42e3f81c634['h012c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00964] =  I0310077d53ae4ed9904df42e3f81c634['h012c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00965] =  I0310077d53ae4ed9904df42e3f81c634['h012ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00966] =  I0310077d53ae4ed9904df42e3f81c634['h012cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00967] =  I0310077d53ae4ed9904df42e3f81c634['h012ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00968] =  I0310077d53ae4ed9904df42e3f81c634['h012d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00969] =  I0310077d53ae4ed9904df42e3f81c634['h012d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0096a] =  I0310077d53ae4ed9904df42e3f81c634['h012d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0096b] =  I0310077d53ae4ed9904df42e3f81c634['h012d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0096c] =  I0310077d53ae4ed9904df42e3f81c634['h012d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0096d] =  I0310077d53ae4ed9904df42e3f81c634['h012da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0096e] =  I0310077d53ae4ed9904df42e3f81c634['h012dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0096f] =  I0310077d53ae4ed9904df42e3f81c634['h012de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00970] =  I0310077d53ae4ed9904df42e3f81c634['h012e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00971] =  I0310077d53ae4ed9904df42e3f81c634['h012e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00972] =  I0310077d53ae4ed9904df42e3f81c634['h012e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00973] =  I0310077d53ae4ed9904df42e3f81c634['h012e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00974] =  I0310077d53ae4ed9904df42e3f81c634['h012e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00975] =  I0310077d53ae4ed9904df42e3f81c634['h012ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00976] =  I0310077d53ae4ed9904df42e3f81c634['h012ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00977] =  I0310077d53ae4ed9904df42e3f81c634['h012ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00978] =  I0310077d53ae4ed9904df42e3f81c634['h012f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00979] =  I0310077d53ae4ed9904df42e3f81c634['h012f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0097a] =  I0310077d53ae4ed9904df42e3f81c634['h012f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0097b] =  I0310077d53ae4ed9904df42e3f81c634['h012f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0097c] =  I0310077d53ae4ed9904df42e3f81c634['h012f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0097d] =  I0310077d53ae4ed9904df42e3f81c634['h012fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0097e] =  I0310077d53ae4ed9904df42e3f81c634['h012fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0097f] =  I0310077d53ae4ed9904df42e3f81c634['h012fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00980] =  I0310077d53ae4ed9904df42e3f81c634['h01300] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00981] =  I0310077d53ae4ed9904df42e3f81c634['h01302] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00982] =  I0310077d53ae4ed9904df42e3f81c634['h01304] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00983] =  I0310077d53ae4ed9904df42e3f81c634['h01306] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00984] =  I0310077d53ae4ed9904df42e3f81c634['h01308] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00985] =  I0310077d53ae4ed9904df42e3f81c634['h0130a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00986] =  I0310077d53ae4ed9904df42e3f81c634['h0130c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00987] =  I0310077d53ae4ed9904df42e3f81c634['h0130e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00988] =  I0310077d53ae4ed9904df42e3f81c634['h01310] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00989] =  I0310077d53ae4ed9904df42e3f81c634['h01312] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0098a] =  I0310077d53ae4ed9904df42e3f81c634['h01314] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0098b] =  I0310077d53ae4ed9904df42e3f81c634['h01316] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0098c] =  I0310077d53ae4ed9904df42e3f81c634['h01318] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0098d] =  I0310077d53ae4ed9904df42e3f81c634['h0131a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0098e] =  I0310077d53ae4ed9904df42e3f81c634['h0131c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0098f] =  I0310077d53ae4ed9904df42e3f81c634['h0131e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00990] =  I0310077d53ae4ed9904df42e3f81c634['h01320] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00991] =  I0310077d53ae4ed9904df42e3f81c634['h01322] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00992] =  I0310077d53ae4ed9904df42e3f81c634['h01324] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00993] =  I0310077d53ae4ed9904df42e3f81c634['h01326] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00994] =  I0310077d53ae4ed9904df42e3f81c634['h01328] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00995] =  I0310077d53ae4ed9904df42e3f81c634['h0132a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00996] =  I0310077d53ae4ed9904df42e3f81c634['h0132c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00997] =  I0310077d53ae4ed9904df42e3f81c634['h0132e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00998] =  I0310077d53ae4ed9904df42e3f81c634['h01330] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00999] =  I0310077d53ae4ed9904df42e3f81c634['h01332] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0099a] =  I0310077d53ae4ed9904df42e3f81c634['h01334] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0099b] =  I0310077d53ae4ed9904df42e3f81c634['h01336] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0099c] =  I0310077d53ae4ed9904df42e3f81c634['h01338] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0099d] =  I0310077d53ae4ed9904df42e3f81c634['h0133a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0099e] =  I0310077d53ae4ed9904df42e3f81c634['h0133c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0099f] =  I0310077d53ae4ed9904df42e3f81c634['h0133e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a0] =  I0310077d53ae4ed9904df42e3f81c634['h01340] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a1] =  I0310077d53ae4ed9904df42e3f81c634['h01342] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a2] =  I0310077d53ae4ed9904df42e3f81c634['h01344] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a3] =  I0310077d53ae4ed9904df42e3f81c634['h01346] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a4] =  I0310077d53ae4ed9904df42e3f81c634['h01348] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a5] =  I0310077d53ae4ed9904df42e3f81c634['h0134a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a6] =  I0310077d53ae4ed9904df42e3f81c634['h0134c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a7] =  I0310077d53ae4ed9904df42e3f81c634['h0134e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a8] =  I0310077d53ae4ed9904df42e3f81c634['h01350] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009a9] =  I0310077d53ae4ed9904df42e3f81c634['h01352] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009aa] =  I0310077d53ae4ed9904df42e3f81c634['h01354] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ab] =  I0310077d53ae4ed9904df42e3f81c634['h01356] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ac] =  I0310077d53ae4ed9904df42e3f81c634['h01358] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ad] =  I0310077d53ae4ed9904df42e3f81c634['h0135a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ae] =  I0310077d53ae4ed9904df42e3f81c634['h0135c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009af] =  I0310077d53ae4ed9904df42e3f81c634['h0135e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b0] =  I0310077d53ae4ed9904df42e3f81c634['h01360] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b1] =  I0310077d53ae4ed9904df42e3f81c634['h01362] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b2] =  I0310077d53ae4ed9904df42e3f81c634['h01364] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b3] =  I0310077d53ae4ed9904df42e3f81c634['h01366] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b4] =  I0310077d53ae4ed9904df42e3f81c634['h01368] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b5] =  I0310077d53ae4ed9904df42e3f81c634['h0136a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b6] =  I0310077d53ae4ed9904df42e3f81c634['h0136c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b7] =  I0310077d53ae4ed9904df42e3f81c634['h0136e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b8] =  I0310077d53ae4ed9904df42e3f81c634['h01370] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009b9] =  I0310077d53ae4ed9904df42e3f81c634['h01372] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ba] =  I0310077d53ae4ed9904df42e3f81c634['h01374] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009bb] =  I0310077d53ae4ed9904df42e3f81c634['h01376] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009bc] =  I0310077d53ae4ed9904df42e3f81c634['h01378] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009bd] =  I0310077d53ae4ed9904df42e3f81c634['h0137a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009be] =  I0310077d53ae4ed9904df42e3f81c634['h0137c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009bf] =  I0310077d53ae4ed9904df42e3f81c634['h0137e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c0] =  I0310077d53ae4ed9904df42e3f81c634['h01380] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c1] =  I0310077d53ae4ed9904df42e3f81c634['h01382] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c2] =  I0310077d53ae4ed9904df42e3f81c634['h01384] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c3] =  I0310077d53ae4ed9904df42e3f81c634['h01386] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c4] =  I0310077d53ae4ed9904df42e3f81c634['h01388] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c5] =  I0310077d53ae4ed9904df42e3f81c634['h0138a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c6] =  I0310077d53ae4ed9904df42e3f81c634['h0138c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c7] =  I0310077d53ae4ed9904df42e3f81c634['h0138e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c8] =  I0310077d53ae4ed9904df42e3f81c634['h01390] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009c9] =  I0310077d53ae4ed9904df42e3f81c634['h01392] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ca] =  I0310077d53ae4ed9904df42e3f81c634['h01394] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009cb] =  I0310077d53ae4ed9904df42e3f81c634['h01396] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009cc] =  I0310077d53ae4ed9904df42e3f81c634['h01398] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009cd] =  I0310077d53ae4ed9904df42e3f81c634['h0139a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ce] =  I0310077d53ae4ed9904df42e3f81c634['h0139c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009cf] =  I0310077d53ae4ed9904df42e3f81c634['h0139e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d0] =  I0310077d53ae4ed9904df42e3f81c634['h013a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d1] =  I0310077d53ae4ed9904df42e3f81c634['h013a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d2] =  I0310077d53ae4ed9904df42e3f81c634['h013a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d3] =  I0310077d53ae4ed9904df42e3f81c634['h013a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d4] =  I0310077d53ae4ed9904df42e3f81c634['h013a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d5] =  I0310077d53ae4ed9904df42e3f81c634['h013aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d6] =  I0310077d53ae4ed9904df42e3f81c634['h013ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d7] =  I0310077d53ae4ed9904df42e3f81c634['h013ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d8] =  I0310077d53ae4ed9904df42e3f81c634['h013b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009d9] =  I0310077d53ae4ed9904df42e3f81c634['h013b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009da] =  I0310077d53ae4ed9904df42e3f81c634['h013b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009db] =  I0310077d53ae4ed9904df42e3f81c634['h013b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009dc] =  I0310077d53ae4ed9904df42e3f81c634['h013b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009dd] =  I0310077d53ae4ed9904df42e3f81c634['h013ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009de] =  I0310077d53ae4ed9904df42e3f81c634['h013bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009df] =  I0310077d53ae4ed9904df42e3f81c634['h013be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e0] =  I0310077d53ae4ed9904df42e3f81c634['h013c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e1] =  I0310077d53ae4ed9904df42e3f81c634['h013c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e2] =  I0310077d53ae4ed9904df42e3f81c634['h013c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e3] =  I0310077d53ae4ed9904df42e3f81c634['h013c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e4] =  I0310077d53ae4ed9904df42e3f81c634['h013c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e5] =  I0310077d53ae4ed9904df42e3f81c634['h013ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e6] =  I0310077d53ae4ed9904df42e3f81c634['h013cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e7] =  I0310077d53ae4ed9904df42e3f81c634['h013ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e8] =  I0310077d53ae4ed9904df42e3f81c634['h013d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009e9] =  I0310077d53ae4ed9904df42e3f81c634['h013d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ea] =  I0310077d53ae4ed9904df42e3f81c634['h013d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009eb] =  I0310077d53ae4ed9904df42e3f81c634['h013d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ec] =  I0310077d53ae4ed9904df42e3f81c634['h013d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ed] =  I0310077d53ae4ed9904df42e3f81c634['h013da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ee] =  I0310077d53ae4ed9904df42e3f81c634['h013dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ef] =  I0310077d53ae4ed9904df42e3f81c634['h013de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f0] =  I0310077d53ae4ed9904df42e3f81c634['h013e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f1] =  I0310077d53ae4ed9904df42e3f81c634['h013e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f2] =  I0310077d53ae4ed9904df42e3f81c634['h013e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f3] =  I0310077d53ae4ed9904df42e3f81c634['h013e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f4] =  I0310077d53ae4ed9904df42e3f81c634['h013e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f5] =  I0310077d53ae4ed9904df42e3f81c634['h013ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f6] =  I0310077d53ae4ed9904df42e3f81c634['h013ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f7] =  I0310077d53ae4ed9904df42e3f81c634['h013ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f8] =  I0310077d53ae4ed9904df42e3f81c634['h013f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009f9] =  I0310077d53ae4ed9904df42e3f81c634['h013f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009fa] =  I0310077d53ae4ed9904df42e3f81c634['h013f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009fb] =  I0310077d53ae4ed9904df42e3f81c634['h013f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009fc] =  I0310077d53ae4ed9904df42e3f81c634['h013f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009fd] =  I0310077d53ae4ed9904df42e3f81c634['h013fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009fe] =  I0310077d53ae4ed9904df42e3f81c634['h013fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h009ff] =  I0310077d53ae4ed9904df42e3f81c634['h013fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a00] =  I0310077d53ae4ed9904df42e3f81c634['h01400] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a01] =  I0310077d53ae4ed9904df42e3f81c634['h01402] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a02] =  I0310077d53ae4ed9904df42e3f81c634['h01404] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a03] =  I0310077d53ae4ed9904df42e3f81c634['h01406] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a04] =  I0310077d53ae4ed9904df42e3f81c634['h01408] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a05] =  I0310077d53ae4ed9904df42e3f81c634['h0140a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a06] =  I0310077d53ae4ed9904df42e3f81c634['h0140c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a07] =  I0310077d53ae4ed9904df42e3f81c634['h0140e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a08] =  I0310077d53ae4ed9904df42e3f81c634['h01410] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a09] =  I0310077d53ae4ed9904df42e3f81c634['h01412] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a0a] =  I0310077d53ae4ed9904df42e3f81c634['h01414] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a0b] =  I0310077d53ae4ed9904df42e3f81c634['h01416] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a0c] =  I0310077d53ae4ed9904df42e3f81c634['h01418] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a0d] =  I0310077d53ae4ed9904df42e3f81c634['h0141a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a0e] =  I0310077d53ae4ed9904df42e3f81c634['h0141c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a0f] =  I0310077d53ae4ed9904df42e3f81c634['h0141e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a10] =  I0310077d53ae4ed9904df42e3f81c634['h01420] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a11] =  I0310077d53ae4ed9904df42e3f81c634['h01422] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a12] =  I0310077d53ae4ed9904df42e3f81c634['h01424] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a13] =  I0310077d53ae4ed9904df42e3f81c634['h01426] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a14] =  I0310077d53ae4ed9904df42e3f81c634['h01428] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a15] =  I0310077d53ae4ed9904df42e3f81c634['h0142a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a16] =  I0310077d53ae4ed9904df42e3f81c634['h0142c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a17] =  I0310077d53ae4ed9904df42e3f81c634['h0142e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a18] =  I0310077d53ae4ed9904df42e3f81c634['h01430] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a19] =  I0310077d53ae4ed9904df42e3f81c634['h01432] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a1a] =  I0310077d53ae4ed9904df42e3f81c634['h01434] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a1b] =  I0310077d53ae4ed9904df42e3f81c634['h01436] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a1c] =  I0310077d53ae4ed9904df42e3f81c634['h01438] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a1d] =  I0310077d53ae4ed9904df42e3f81c634['h0143a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a1e] =  I0310077d53ae4ed9904df42e3f81c634['h0143c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a1f] =  I0310077d53ae4ed9904df42e3f81c634['h0143e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a20] =  I0310077d53ae4ed9904df42e3f81c634['h01440] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a21] =  I0310077d53ae4ed9904df42e3f81c634['h01442] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a22] =  I0310077d53ae4ed9904df42e3f81c634['h01444] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a23] =  I0310077d53ae4ed9904df42e3f81c634['h01446] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a24] =  I0310077d53ae4ed9904df42e3f81c634['h01448] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a25] =  I0310077d53ae4ed9904df42e3f81c634['h0144a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a26] =  I0310077d53ae4ed9904df42e3f81c634['h0144c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a27] =  I0310077d53ae4ed9904df42e3f81c634['h0144e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a28] =  I0310077d53ae4ed9904df42e3f81c634['h01450] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a29] =  I0310077d53ae4ed9904df42e3f81c634['h01452] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a2a] =  I0310077d53ae4ed9904df42e3f81c634['h01454] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a2b] =  I0310077d53ae4ed9904df42e3f81c634['h01456] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a2c] =  I0310077d53ae4ed9904df42e3f81c634['h01458] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a2d] =  I0310077d53ae4ed9904df42e3f81c634['h0145a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a2e] =  I0310077d53ae4ed9904df42e3f81c634['h0145c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a2f] =  I0310077d53ae4ed9904df42e3f81c634['h0145e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a30] =  I0310077d53ae4ed9904df42e3f81c634['h01460] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a31] =  I0310077d53ae4ed9904df42e3f81c634['h01462] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a32] =  I0310077d53ae4ed9904df42e3f81c634['h01464] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a33] =  I0310077d53ae4ed9904df42e3f81c634['h01466] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a34] =  I0310077d53ae4ed9904df42e3f81c634['h01468] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a35] =  I0310077d53ae4ed9904df42e3f81c634['h0146a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a36] =  I0310077d53ae4ed9904df42e3f81c634['h0146c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a37] =  I0310077d53ae4ed9904df42e3f81c634['h0146e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a38] =  I0310077d53ae4ed9904df42e3f81c634['h01470] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a39] =  I0310077d53ae4ed9904df42e3f81c634['h01472] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a3a] =  I0310077d53ae4ed9904df42e3f81c634['h01474] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a3b] =  I0310077d53ae4ed9904df42e3f81c634['h01476] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a3c] =  I0310077d53ae4ed9904df42e3f81c634['h01478] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a3d] =  I0310077d53ae4ed9904df42e3f81c634['h0147a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a3e] =  I0310077d53ae4ed9904df42e3f81c634['h0147c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a3f] =  I0310077d53ae4ed9904df42e3f81c634['h0147e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a40] =  I0310077d53ae4ed9904df42e3f81c634['h01480] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a41] =  I0310077d53ae4ed9904df42e3f81c634['h01482] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a42] =  I0310077d53ae4ed9904df42e3f81c634['h01484] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a43] =  I0310077d53ae4ed9904df42e3f81c634['h01486] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a44] =  I0310077d53ae4ed9904df42e3f81c634['h01488] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a45] =  I0310077d53ae4ed9904df42e3f81c634['h0148a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a46] =  I0310077d53ae4ed9904df42e3f81c634['h0148c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a47] =  I0310077d53ae4ed9904df42e3f81c634['h0148e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a48] =  I0310077d53ae4ed9904df42e3f81c634['h01490] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a49] =  I0310077d53ae4ed9904df42e3f81c634['h01492] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a4a] =  I0310077d53ae4ed9904df42e3f81c634['h01494] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a4b] =  I0310077d53ae4ed9904df42e3f81c634['h01496] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a4c] =  I0310077d53ae4ed9904df42e3f81c634['h01498] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a4d] =  I0310077d53ae4ed9904df42e3f81c634['h0149a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a4e] =  I0310077d53ae4ed9904df42e3f81c634['h0149c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a4f] =  I0310077d53ae4ed9904df42e3f81c634['h0149e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a50] =  I0310077d53ae4ed9904df42e3f81c634['h014a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a51] =  I0310077d53ae4ed9904df42e3f81c634['h014a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a52] =  I0310077d53ae4ed9904df42e3f81c634['h014a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a53] =  I0310077d53ae4ed9904df42e3f81c634['h014a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a54] =  I0310077d53ae4ed9904df42e3f81c634['h014a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a55] =  I0310077d53ae4ed9904df42e3f81c634['h014aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a56] =  I0310077d53ae4ed9904df42e3f81c634['h014ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a57] =  I0310077d53ae4ed9904df42e3f81c634['h014ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a58] =  I0310077d53ae4ed9904df42e3f81c634['h014b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a59] =  I0310077d53ae4ed9904df42e3f81c634['h014b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a5a] =  I0310077d53ae4ed9904df42e3f81c634['h014b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a5b] =  I0310077d53ae4ed9904df42e3f81c634['h014b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a5c] =  I0310077d53ae4ed9904df42e3f81c634['h014b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a5d] =  I0310077d53ae4ed9904df42e3f81c634['h014ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a5e] =  I0310077d53ae4ed9904df42e3f81c634['h014bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a5f] =  I0310077d53ae4ed9904df42e3f81c634['h014be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a60] =  I0310077d53ae4ed9904df42e3f81c634['h014c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a61] =  I0310077d53ae4ed9904df42e3f81c634['h014c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a62] =  I0310077d53ae4ed9904df42e3f81c634['h014c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a63] =  I0310077d53ae4ed9904df42e3f81c634['h014c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a64] =  I0310077d53ae4ed9904df42e3f81c634['h014c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a65] =  I0310077d53ae4ed9904df42e3f81c634['h014ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a66] =  I0310077d53ae4ed9904df42e3f81c634['h014cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a67] =  I0310077d53ae4ed9904df42e3f81c634['h014ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a68] =  I0310077d53ae4ed9904df42e3f81c634['h014d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a69] =  I0310077d53ae4ed9904df42e3f81c634['h014d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a6a] =  I0310077d53ae4ed9904df42e3f81c634['h014d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a6b] =  I0310077d53ae4ed9904df42e3f81c634['h014d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a6c] =  I0310077d53ae4ed9904df42e3f81c634['h014d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a6d] =  I0310077d53ae4ed9904df42e3f81c634['h014da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a6e] =  I0310077d53ae4ed9904df42e3f81c634['h014dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a6f] =  I0310077d53ae4ed9904df42e3f81c634['h014de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a70] =  I0310077d53ae4ed9904df42e3f81c634['h014e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a71] =  I0310077d53ae4ed9904df42e3f81c634['h014e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a72] =  I0310077d53ae4ed9904df42e3f81c634['h014e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a73] =  I0310077d53ae4ed9904df42e3f81c634['h014e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a74] =  I0310077d53ae4ed9904df42e3f81c634['h014e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a75] =  I0310077d53ae4ed9904df42e3f81c634['h014ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a76] =  I0310077d53ae4ed9904df42e3f81c634['h014ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a77] =  I0310077d53ae4ed9904df42e3f81c634['h014ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a78] =  I0310077d53ae4ed9904df42e3f81c634['h014f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a79] =  I0310077d53ae4ed9904df42e3f81c634['h014f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a7a] =  I0310077d53ae4ed9904df42e3f81c634['h014f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a7b] =  I0310077d53ae4ed9904df42e3f81c634['h014f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a7c] =  I0310077d53ae4ed9904df42e3f81c634['h014f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a7d] =  I0310077d53ae4ed9904df42e3f81c634['h014fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a7e] =  I0310077d53ae4ed9904df42e3f81c634['h014fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a7f] =  I0310077d53ae4ed9904df42e3f81c634['h014fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a80] =  I0310077d53ae4ed9904df42e3f81c634['h01500] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a81] =  I0310077d53ae4ed9904df42e3f81c634['h01502] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a82] =  I0310077d53ae4ed9904df42e3f81c634['h01504] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a83] =  I0310077d53ae4ed9904df42e3f81c634['h01506] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a84] =  I0310077d53ae4ed9904df42e3f81c634['h01508] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a85] =  I0310077d53ae4ed9904df42e3f81c634['h0150a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a86] =  I0310077d53ae4ed9904df42e3f81c634['h0150c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a87] =  I0310077d53ae4ed9904df42e3f81c634['h0150e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a88] =  I0310077d53ae4ed9904df42e3f81c634['h01510] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a89] =  I0310077d53ae4ed9904df42e3f81c634['h01512] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a8a] =  I0310077d53ae4ed9904df42e3f81c634['h01514] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a8b] =  I0310077d53ae4ed9904df42e3f81c634['h01516] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a8c] =  I0310077d53ae4ed9904df42e3f81c634['h01518] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a8d] =  I0310077d53ae4ed9904df42e3f81c634['h0151a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a8e] =  I0310077d53ae4ed9904df42e3f81c634['h0151c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a8f] =  I0310077d53ae4ed9904df42e3f81c634['h0151e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a90] =  I0310077d53ae4ed9904df42e3f81c634['h01520] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a91] =  I0310077d53ae4ed9904df42e3f81c634['h01522] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a92] =  I0310077d53ae4ed9904df42e3f81c634['h01524] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a93] =  I0310077d53ae4ed9904df42e3f81c634['h01526] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a94] =  I0310077d53ae4ed9904df42e3f81c634['h01528] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a95] =  I0310077d53ae4ed9904df42e3f81c634['h0152a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a96] =  I0310077d53ae4ed9904df42e3f81c634['h0152c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a97] =  I0310077d53ae4ed9904df42e3f81c634['h0152e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a98] =  I0310077d53ae4ed9904df42e3f81c634['h01530] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a99] =  I0310077d53ae4ed9904df42e3f81c634['h01532] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a9a] =  I0310077d53ae4ed9904df42e3f81c634['h01534] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a9b] =  I0310077d53ae4ed9904df42e3f81c634['h01536] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a9c] =  I0310077d53ae4ed9904df42e3f81c634['h01538] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a9d] =  I0310077d53ae4ed9904df42e3f81c634['h0153a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a9e] =  I0310077d53ae4ed9904df42e3f81c634['h0153c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00a9f] =  I0310077d53ae4ed9904df42e3f81c634['h0153e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa0] =  I0310077d53ae4ed9904df42e3f81c634['h01540] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa1] =  I0310077d53ae4ed9904df42e3f81c634['h01542] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa2] =  I0310077d53ae4ed9904df42e3f81c634['h01544] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa3] =  I0310077d53ae4ed9904df42e3f81c634['h01546] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa4] =  I0310077d53ae4ed9904df42e3f81c634['h01548] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa5] =  I0310077d53ae4ed9904df42e3f81c634['h0154a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa6] =  I0310077d53ae4ed9904df42e3f81c634['h0154c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa7] =  I0310077d53ae4ed9904df42e3f81c634['h0154e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa8] =  I0310077d53ae4ed9904df42e3f81c634['h01550] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aa9] =  I0310077d53ae4ed9904df42e3f81c634['h01552] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aaa] =  I0310077d53ae4ed9904df42e3f81c634['h01554] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aab] =  I0310077d53ae4ed9904df42e3f81c634['h01556] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aac] =  I0310077d53ae4ed9904df42e3f81c634['h01558] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aad] =  I0310077d53ae4ed9904df42e3f81c634['h0155a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aae] =  I0310077d53ae4ed9904df42e3f81c634['h0155c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aaf] =  I0310077d53ae4ed9904df42e3f81c634['h0155e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab0] =  I0310077d53ae4ed9904df42e3f81c634['h01560] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab1] =  I0310077d53ae4ed9904df42e3f81c634['h01562] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab2] =  I0310077d53ae4ed9904df42e3f81c634['h01564] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab3] =  I0310077d53ae4ed9904df42e3f81c634['h01566] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab4] =  I0310077d53ae4ed9904df42e3f81c634['h01568] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab5] =  I0310077d53ae4ed9904df42e3f81c634['h0156a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab6] =  I0310077d53ae4ed9904df42e3f81c634['h0156c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab7] =  I0310077d53ae4ed9904df42e3f81c634['h0156e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab8] =  I0310077d53ae4ed9904df42e3f81c634['h01570] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ab9] =  I0310077d53ae4ed9904df42e3f81c634['h01572] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aba] =  I0310077d53ae4ed9904df42e3f81c634['h01574] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00abb] =  I0310077d53ae4ed9904df42e3f81c634['h01576] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00abc] =  I0310077d53ae4ed9904df42e3f81c634['h01578] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00abd] =  I0310077d53ae4ed9904df42e3f81c634['h0157a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00abe] =  I0310077d53ae4ed9904df42e3f81c634['h0157c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00abf] =  I0310077d53ae4ed9904df42e3f81c634['h0157e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac0] =  I0310077d53ae4ed9904df42e3f81c634['h01580] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac1] =  I0310077d53ae4ed9904df42e3f81c634['h01582] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac2] =  I0310077d53ae4ed9904df42e3f81c634['h01584] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac3] =  I0310077d53ae4ed9904df42e3f81c634['h01586] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac4] =  I0310077d53ae4ed9904df42e3f81c634['h01588] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac5] =  I0310077d53ae4ed9904df42e3f81c634['h0158a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac6] =  I0310077d53ae4ed9904df42e3f81c634['h0158c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac7] =  I0310077d53ae4ed9904df42e3f81c634['h0158e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac8] =  I0310077d53ae4ed9904df42e3f81c634['h01590] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ac9] =  I0310077d53ae4ed9904df42e3f81c634['h01592] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aca] =  I0310077d53ae4ed9904df42e3f81c634['h01594] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00acb] =  I0310077d53ae4ed9904df42e3f81c634['h01596] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00acc] =  I0310077d53ae4ed9904df42e3f81c634['h01598] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00acd] =  I0310077d53ae4ed9904df42e3f81c634['h0159a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ace] =  I0310077d53ae4ed9904df42e3f81c634['h0159c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00acf] =  I0310077d53ae4ed9904df42e3f81c634['h0159e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad0] =  I0310077d53ae4ed9904df42e3f81c634['h015a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad1] =  I0310077d53ae4ed9904df42e3f81c634['h015a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad2] =  I0310077d53ae4ed9904df42e3f81c634['h015a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad3] =  I0310077d53ae4ed9904df42e3f81c634['h015a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad4] =  I0310077d53ae4ed9904df42e3f81c634['h015a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad5] =  I0310077d53ae4ed9904df42e3f81c634['h015aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad6] =  I0310077d53ae4ed9904df42e3f81c634['h015ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad7] =  I0310077d53ae4ed9904df42e3f81c634['h015ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad8] =  I0310077d53ae4ed9904df42e3f81c634['h015b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ad9] =  I0310077d53ae4ed9904df42e3f81c634['h015b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ada] =  I0310077d53ae4ed9904df42e3f81c634['h015b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00adb] =  I0310077d53ae4ed9904df42e3f81c634['h015b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00adc] =  I0310077d53ae4ed9904df42e3f81c634['h015b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00add] =  I0310077d53ae4ed9904df42e3f81c634['h015ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ade] =  I0310077d53ae4ed9904df42e3f81c634['h015bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00adf] =  I0310077d53ae4ed9904df42e3f81c634['h015be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae0] =  I0310077d53ae4ed9904df42e3f81c634['h015c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae1] =  I0310077d53ae4ed9904df42e3f81c634['h015c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae2] =  I0310077d53ae4ed9904df42e3f81c634['h015c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae3] =  I0310077d53ae4ed9904df42e3f81c634['h015c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae4] =  I0310077d53ae4ed9904df42e3f81c634['h015c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae5] =  I0310077d53ae4ed9904df42e3f81c634['h015ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae6] =  I0310077d53ae4ed9904df42e3f81c634['h015cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae7] =  I0310077d53ae4ed9904df42e3f81c634['h015ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae8] =  I0310077d53ae4ed9904df42e3f81c634['h015d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ae9] =  I0310077d53ae4ed9904df42e3f81c634['h015d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aea] =  I0310077d53ae4ed9904df42e3f81c634['h015d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aeb] =  I0310077d53ae4ed9904df42e3f81c634['h015d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aec] =  I0310077d53ae4ed9904df42e3f81c634['h015d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aed] =  I0310077d53ae4ed9904df42e3f81c634['h015da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aee] =  I0310077d53ae4ed9904df42e3f81c634['h015dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aef] =  I0310077d53ae4ed9904df42e3f81c634['h015de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af0] =  I0310077d53ae4ed9904df42e3f81c634['h015e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af1] =  I0310077d53ae4ed9904df42e3f81c634['h015e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af2] =  I0310077d53ae4ed9904df42e3f81c634['h015e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af3] =  I0310077d53ae4ed9904df42e3f81c634['h015e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af4] =  I0310077d53ae4ed9904df42e3f81c634['h015e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af5] =  I0310077d53ae4ed9904df42e3f81c634['h015ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af6] =  I0310077d53ae4ed9904df42e3f81c634['h015ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af7] =  I0310077d53ae4ed9904df42e3f81c634['h015ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af8] =  I0310077d53ae4ed9904df42e3f81c634['h015f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00af9] =  I0310077d53ae4ed9904df42e3f81c634['h015f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00afa] =  I0310077d53ae4ed9904df42e3f81c634['h015f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00afb] =  I0310077d53ae4ed9904df42e3f81c634['h015f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00afc] =  I0310077d53ae4ed9904df42e3f81c634['h015f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00afd] =  I0310077d53ae4ed9904df42e3f81c634['h015fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00afe] =  I0310077d53ae4ed9904df42e3f81c634['h015fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00aff] =  I0310077d53ae4ed9904df42e3f81c634['h015fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b00] =  I0310077d53ae4ed9904df42e3f81c634['h01600] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b01] =  I0310077d53ae4ed9904df42e3f81c634['h01602] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b02] =  I0310077d53ae4ed9904df42e3f81c634['h01604] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b03] =  I0310077d53ae4ed9904df42e3f81c634['h01606] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b04] =  I0310077d53ae4ed9904df42e3f81c634['h01608] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b05] =  I0310077d53ae4ed9904df42e3f81c634['h0160a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b06] =  I0310077d53ae4ed9904df42e3f81c634['h0160c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b07] =  I0310077d53ae4ed9904df42e3f81c634['h0160e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b08] =  I0310077d53ae4ed9904df42e3f81c634['h01610] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b09] =  I0310077d53ae4ed9904df42e3f81c634['h01612] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b0a] =  I0310077d53ae4ed9904df42e3f81c634['h01614] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b0b] =  I0310077d53ae4ed9904df42e3f81c634['h01616] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b0c] =  I0310077d53ae4ed9904df42e3f81c634['h01618] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b0d] =  I0310077d53ae4ed9904df42e3f81c634['h0161a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b0e] =  I0310077d53ae4ed9904df42e3f81c634['h0161c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b0f] =  I0310077d53ae4ed9904df42e3f81c634['h0161e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b10] =  I0310077d53ae4ed9904df42e3f81c634['h01620] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b11] =  I0310077d53ae4ed9904df42e3f81c634['h01622] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b12] =  I0310077d53ae4ed9904df42e3f81c634['h01624] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b13] =  I0310077d53ae4ed9904df42e3f81c634['h01626] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b14] =  I0310077d53ae4ed9904df42e3f81c634['h01628] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b15] =  I0310077d53ae4ed9904df42e3f81c634['h0162a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b16] =  I0310077d53ae4ed9904df42e3f81c634['h0162c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b17] =  I0310077d53ae4ed9904df42e3f81c634['h0162e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b18] =  I0310077d53ae4ed9904df42e3f81c634['h01630] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b19] =  I0310077d53ae4ed9904df42e3f81c634['h01632] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b1a] =  I0310077d53ae4ed9904df42e3f81c634['h01634] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b1b] =  I0310077d53ae4ed9904df42e3f81c634['h01636] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b1c] =  I0310077d53ae4ed9904df42e3f81c634['h01638] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b1d] =  I0310077d53ae4ed9904df42e3f81c634['h0163a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b1e] =  I0310077d53ae4ed9904df42e3f81c634['h0163c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b1f] =  I0310077d53ae4ed9904df42e3f81c634['h0163e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b20] =  I0310077d53ae4ed9904df42e3f81c634['h01640] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b21] =  I0310077d53ae4ed9904df42e3f81c634['h01642] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b22] =  I0310077d53ae4ed9904df42e3f81c634['h01644] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b23] =  I0310077d53ae4ed9904df42e3f81c634['h01646] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b24] =  I0310077d53ae4ed9904df42e3f81c634['h01648] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b25] =  I0310077d53ae4ed9904df42e3f81c634['h0164a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b26] =  I0310077d53ae4ed9904df42e3f81c634['h0164c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b27] =  I0310077d53ae4ed9904df42e3f81c634['h0164e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b28] =  I0310077d53ae4ed9904df42e3f81c634['h01650] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b29] =  I0310077d53ae4ed9904df42e3f81c634['h01652] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b2a] =  I0310077d53ae4ed9904df42e3f81c634['h01654] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b2b] =  I0310077d53ae4ed9904df42e3f81c634['h01656] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b2c] =  I0310077d53ae4ed9904df42e3f81c634['h01658] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b2d] =  I0310077d53ae4ed9904df42e3f81c634['h0165a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b2e] =  I0310077d53ae4ed9904df42e3f81c634['h0165c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b2f] =  I0310077d53ae4ed9904df42e3f81c634['h0165e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b30] =  I0310077d53ae4ed9904df42e3f81c634['h01660] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b31] =  I0310077d53ae4ed9904df42e3f81c634['h01662] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b32] =  I0310077d53ae4ed9904df42e3f81c634['h01664] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b33] =  I0310077d53ae4ed9904df42e3f81c634['h01666] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b34] =  I0310077d53ae4ed9904df42e3f81c634['h01668] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b35] =  I0310077d53ae4ed9904df42e3f81c634['h0166a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b36] =  I0310077d53ae4ed9904df42e3f81c634['h0166c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b37] =  I0310077d53ae4ed9904df42e3f81c634['h0166e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b38] =  I0310077d53ae4ed9904df42e3f81c634['h01670] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b39] =  I0310077d53ae4ed9904df42e3f81c634['h01672] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b3a] =  I0310077d53ae4ed9904df42e3f81c634['h01674] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b3b] =  I0310077d53ae4ed9904df42e3f81c634['h01676] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b3c] =  I0310077d53ae4ed9904df42e3f81c634['h01678] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b3d] =  I0310077d53ae4ed9904df42e3f81c634['h0167a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b3e] =  I0310077d53ae4ed9904df42e3f81c634['h0167c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b3f] =  I0310077d53ae4ed9904df42e3f81c634['h0167e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b40] =  I0310077d53ae4ed9904df42e3f81c634['h01680] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b41] =  I0310077d53ae4ed9904df42e3f81c634['h01682] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b42] =  I0310077d53ae4ed9904df42e3f81c634['h01684] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b43] =  I0310077d53ae4ed9904df42e3f81c634['h01686] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b44] =  I0310077d53ae4ed9904df42e3f81c634['h01688] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b45] =  I0310077d53ae4ed9904df42e3f81c634['h0168a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b46] =  I0310077d53ae4ed9904df42e3f81c634['h0168c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b47] =  I0310077d53ae4ed9904df42e3f81c634['h0168e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b48] =  I0310077d53ae4ed9904df42e3f81c634['h01690] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b49] =  I0310077d53ae4ed9904df42e3f81c634['h01692] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b4a] =  I0310077d53ae4ed9904df42e3f81c634['h01694] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b4b] =  I0310077d53ae4ed9904df42e3f81c634['h01696] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b4c] =  I0310077d53ae4ed9904df42e3f81c634['h01698] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b4d] =  I0310077d53ae4ed9904df42e3f81c634['h0169a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b4e] =  I0310077d53ae4ed9904df42e3f81c634['h0169c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b4f] =  I0310077d53ae4ed9904df42e3f81c634['h0169e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b50] =  I0310077d53ae4ed9904df42e3f81c634['h016a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b51] =  I0310077d53ae4ed9904df42e3f81c634['h016a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b52] =  I0310077d53ae4ed9904df42e3f81c634['h016a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b53] =  I0310077d53ae4ed9904df42e3f81c634['h016a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b54] =  I0310077d53ae4ed9904df42e3f81c634['h016a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b55] =  I0310077d53ae4ed9904df42e3f81c634['h016aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b56] =  I0310077d53ae4ed9904df42e3f81c634['h016ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b57] =  I0310077d53ae4ed9904df42e3f81c634['h016ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b58] =  I0310077d53ae4ed9904df42e3f81c634['h016b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b59] =  I0310077d53ae4ed9904df42e3f81c634['h016b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b5a] =  I0310077d53ae4ed9904df42e3f81c634['h016b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b5b] =  I0310077d53ae4ed9904df42e3f81c634['h016b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b5c] =  I0310077d53ae4ed9904df42e3f81c634['h016b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b5d] =  I0310077d53ae4ed9904df42e3f81c634['h016ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b5e] =  I0310077d53ae4ed9904df42e3f81c634['h016bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b5f] =  I0310077d53ae4ed9904df42e3f81c634['h016be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b60] =  I0310077d53ae4ed9904df42e3f81c634['h016c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b61] =  I0310077d53ae4ed9904df42e3f81c634['h016c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b62] =  I0310077d53ae4ed9904df42e3f81c634['h016c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b63] =  I0310077d53ae4ed9904df42e3f81c634['h016c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b64] =  I0310077d53ae4ed9904df42e3f81c634['h016c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b65] =  I0310077d53ae4ed9904df42e3f81c634['h016ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b66] =  I0310077d53ae4ed9904df42e3f81c634['h016cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b67] =  I0310077d53ae4ed9904df42e3f81c634['h016ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b68] =  I0310077d53ae4ed9904df42e3f81c634['h016d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b69] =  I0310077d53ae4ed9904df42e3f81c634['h016d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b6a] =  I0310077d53ae4ed9904df42e3f81c634['h016d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b6b] =  I0310077d53ae4ed9904df42e3f81c634['h016d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b6c] =  I0310077d53ae4ed9904df42e3f81c634['h016d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b6d] =  I0310077d53ae4ed9904df42e3f81c634['h016da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b6e] =  I0310077d53ae4ed9904df42e3f81c634['h016dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b6f] =  I0310077d53ae4ed9904df42e3f81c634['h016de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b70] =  I0310077d53ae4ed9904df42e3f81c634['h016e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b71] =  I0310077d53ae4ed9904df42e3f81c634['h016e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b72] =  I0310077d53ae4ed9904df42e3f81c634['h016e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b73] =  I0310077d53ae4ed9904df42e3f81c634['h016e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b74] =  I0310077d53ae4ed9904df42e3f81c634['h016e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b75] =  I0310077d53ae4ed9904df42e3f81c634['h016ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b76] =  I0310077d53ae4ed9904df42e3f81c634['h016ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b77] =  I0310077d53ae4ed9904df42e3f81c634['h016ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b78] =  I0310077d53ae4ed9904df42e3f81c634['h016f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b79] =  I0310077d53ae4ed9904df42e3f81c634['h016f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b7a] =  I0310077d53ae4ed9904df42e3f81c634['h016f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b7b] =  I0310077d53ae4ed9904df42e3f81c634['h016f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b7c] =  I0310077d53ae4ed9904df42e3f81c634['h016f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b7d] =  I0310077d53ae4ed9904df42e3f81c634['h016fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b7e] =  I0310077d53ae4ed9904df42e3f81c634['h016fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b7f] =  I0310077d53ae4ed9904df42e3f81c634['h016fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b80] =  I0310077d53ae4ed9904df42e3f81c634['h01700] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b81] =  I0310077d53ae4ed9904df42e3f81c634['h01702] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b82] =  I0310077d53ae4ed9904df42e3f81c634['h01704] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b83] =  I0310077d53ae4ed9904df42e3f81c634['h01706] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b84] =  I0310077d53ae4ed9904df42e3f81c634['h01708] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b85] =  I0310077d53ae4ed9904df42e3f81c634['h0170a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b86] =  I0310077d53ae4ed9904df42e3f81c634['h0170c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b87] =  I0310077d53ae4ed9904df42e3f81c634['h0170e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b88] =  I0310077d53ae4ed9904df42e3f81c634['h01710] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b89] =  I0310077d53ae4ed9904df42e3f81c634['h01712] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b8a] =  I0310077d53ae4ed9904df42e3f81c634['h01714] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b8b] =  I0310077d53ae4ed9904df42e3f81c634['h01716] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b8c] =  I0310077d53ae4ed9904df42e3f81c634['h01718] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b8d] =  I0310077d53ae4ed9904df42e3f81c634['h0171a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b8e] =  I0310077d53ae4ed9904df42e3f81c634['h0171c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b8f] =  I0310077d53ae4ed9904df42e3f81c634['h0171e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b90] =  I0310077d53ae4ed9904df42e3f81c634['h01720] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b91] =  I0310077d53ae4ed9904df42e3f81c634['h01722] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b92] =  I0310077d53ae4ed9904df42e3f81c634['h01724] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b93] =  I0310077d53ae4ed9904df42e3f81c634['h01726] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b94] =  I0310077d53ae4ed9904df42e3f81c634['h01728] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b95] =  I0310077d53ae4ed9904df42e3f81c634['h0172a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b96] =  I0310077d53ae4ed9904df42e3f81c634['h0172c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b97] =  I0310077d53ae4ed9904df42e3f81c634['h0172e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b98] =  I0310077d53ae4ed9904df42e3f81c634['h01730] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b99] =  I0310077d53ae4ed9904df42e3f81c634['h01732] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b9a] =  I0310077d53ae4ed9904df42e3f81c634['h01734] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b9b] =  I0310077d53ae4ed9904df42e3f81c634['h01736] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b9c] =  I0310077d53ae4ed9904df42e3f81c634['h01738] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b9d] =  I0310077d53ae4ed9904df42e3f81c634['h0173a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b9e] =  I0310077d53ae4ed9904df42e3f81c634['h0173c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00b9f] =  I0310077d53ae4ed9904df42e3f81c634['h0173e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba0] =  I0310077d53ae4ed9904df42e3f81c634['h01740] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba1] =  I0310077d53ae4ed9904df42e3f81c634['h01742] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba2] =  I0310077d53ae4ed9904df42e3f81c634['h01744] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba3] =  I0310077d53ae4ed9904df42e3f81c634['h01746] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba4] =  I0310077d53ae4ed9904df42e3f81c634['h01748] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba5] =  I0310077d53ae4ed9904df42e3f81c634['h0174a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba6] =  I0310077d53ae4ed9904df42e3f81c634['h0174c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba7] =  I0310077d53ae4ed9904df42e3f81c634['h0174e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba8] =  I0310077d53ae4ed9904df42e3f81c634['h01750] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ba9] =  I0310077d53ae4ed9904df42e3f81c634['h01752] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00baa] =  I0310077d53ae4ed9904df42e3f81c634['h01754] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bab] =  I0310077d53ae4ed9904df42e3f81c634['h01756] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bac] =  I0310077d53ae4ed9904df42e3f81c634['h01758] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bad] =  I0310077d53ae4ed9904df42e3f81c634['h0175a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bae] =  I0310077d53ae4ed9904df42e3f81c634['h0175c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00baf] =  I0310077d53ae4ed9904df42e3f81c634['h0175e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb0] =  I0310077d53ae4ed9904df42e3f81c634['h01760] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb1] =  I0310077d53ae4ed9904df42e3f81c634['h01762] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb2] =  I0310077d53ae4ed9904df42e3f81c634['h01764] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb3] =  I0310077d53ae4ed9904df42e3f81c634['h01766] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb4] =  I0310077d53ae4ed9904df42e3f81c634['h01768] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb5] =  I0310077d53ae4ed9904df42e3f81c634['h0176a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb6] =  I0310077d53ae4ed9904df42e3f81c634['h0176c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb7] =  I0310077d53ae4ed9904df42e3f81c634['h0176e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb8] =  I0310077d53ae4ed9904df42e3f81c634['h01770] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bb9] =  I0310077d53ae4ed9904df42e3f81c634['h01772] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bba] =  I0310077d53ae4ed9904df42e3f81c634['h01774] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bbb] =  I0310077d53ae4ed9904df42e3f81c634['h01776] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bbc] =  I0310077d53ae4ed9904df42e3f81c634['h01778] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bbd] =  I0310077d53ae4ed9904df42e3f81c634['h0177a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bbe] =  I0310077d53ae4ed9904df42e3f81c634['h0177c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bbf] =  I0310077d53ae4ed9904df42e3f81c634['h0177e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc0] =  I0310077d53ae4ed9904df42e3f81c634['h01780] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc1] =  I0310077d53ae4ed9904df42e3f81c634['h01782] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc2] =  I0310077d53ae4ed9904df42e3f81c634['h01784] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc3] =  I0310077d53ae4ed9904df42e3f81c634['h01786] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc4] =  I0310077d53ae4ed9904df42e3f81c634['h01788] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc5] =  I0310077d53ae4ed9904df42e3f81c634['h0178a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc6] =  I0310077d53ae4ed9904df42e3f81c634['h0178c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc7] =  I0310077d53ae4ed9904df42e3f81c634['h0178e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc8] =  I0310077d53ae4ed9904df42e3f81c634['h01790] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bc9] =  I0310077d53ae4ed9904df42e3f81c634['h01792] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bca] =  I0310077d53ae4ed9904df42e3f81c634['h01794] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bcb] =  I0310077d53ae4ed9904df42e3f81c634['h01796] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bcc] =  I0310077d53ae4ed9904df42e3f81c634['h01798] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bcd] =  I0310077d53ae4ed9904df42e3f81c634['h0179a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bce] =  I0310077d53ae4ed9904df42e3f81c634['h0179c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bcf] =  I0310077d53ae4ed9904df42e3f81c634['h0179e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd0] =  I0310077d53ae4ed9904df42e3f81c634['h017a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd1] =  I0310077d53ae4ed9904df42e3f81c634['h017a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd2] =  I0310077d53ae4ed9904df42e3f81c634['h017a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd3] =  I0310077d53ae4ed9904df42e3f81c634['h017a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd4] =  I0310077d53ae4ed9904df42e3f81c634['h017a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd5] =  I0310077d53ae4ed9904df42e3f81c634['h017aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd6] =  I0310077d53ae4ed9904df42e3f81c634['h017ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd7] =  I0310077d53ae4ed9904df42e3f81c634['h017ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd8] =  I0310077d53ae4ed9904df42e3f81c634['h017b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bd9] =  I0310077d53ae4ed9904df42e3f81c634['h017b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bda] =  I0310077d53ae4ed9904df42e3f81c634['h017b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bdb] =  I0310077d53ae4ed9904df42e3f81c634['h017b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bdc] =  I0310077d53ae4ed9904df42e3f81c634['h017b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bdd] =  I0310077d53ae4ed9904df42e3f81c634['h017ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bde] =  I0310077d53ae4ed9904df42e3f81c634['h017bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bdf] =  I0310077d53ae4ed9904df42e3f81c634['h017be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be0] =  I0310077d53ae4ed9904df42e3f81c634['h017c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be1] =  I0310077d53ae4ed9904df42e3f81c634['h017c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be2] =  I0310077d53ae4ed9904df42e3f81c634['h017c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be3] =  I0310077d53ae4ed9904df42e3f81c634['h017c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be4] =  I0310077d53ae4ed9904df42e3f81c634['h017c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be5] =  I0310077d53ae4ed9904df42e3f81c634['h017ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be6] =  I0310077d53ae4ed9904df42e3f81c634['h017cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be7] =  I0310077d53ae4ed9904df42e3f81c634['h017ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be8] =  I0310077d53ae4ed9904df42e3f81c634['h017d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00be9] =  I0310077d53ae4ed9904df42e3f81c634['h017d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bea] =  I0310077d53ae4ed9904df42e3f81c634['h017d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00beb] =  I0310077d53ae4ed9904df42e3f81c634['h017d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bec] =  I0310077d53ae4ed9904df42e3f81c634['h017d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bed] =  I0310077d53ae4ed9904df42e3f81c634['h017da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bee] =  I0310077d53ae4ed9904df42e3f81c634['h017dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bef] =  I0310077d53ae4ed9904df42e3f81c634['h017de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf0] =  I0310077d53ae4ed9904df42e3f81c634['h017e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf1] =  I0310077d53ae4ed9904df42e3f81c634['h017e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf2] =  I0310077d53ae4ed9904df42e3f81c634['h017e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf3] =  I0310077d53ae4ed9904df42e3f81c634['h017e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf4] =  I0310077d53ae4ed9904df42e3f81c634['h017e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf5] =  I0310077d53ae4ed9904df42e3f81c634['h017ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf6] =  I0310077d53ae4ed9904df42e3f81c634['h017ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf7] =  I0310077d53ae4ed9904df42e3f81c634['h017ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf8] =  I0310077d53ae4ed9904df42e3f81c634['h017f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bf9] =  I0310077d53ae4ed9904df42e3f81c634['h017f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bfa] =  I0310077d53ae4ed9904df42e3f81c634['h017f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bfb] =  I0310077d53ae4ed9904df42e3f81c634['h017f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bfc] =  I0310077d53ae4ed9904df42e3f81c634['h017f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bfd] =  I0310077d53ae4ed9904df42e3f81c634['h017fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bfe] =  I0310077d53ae4ed9904df42e3f81c634['h017fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00bff] =  I0310077d53ae4ed9904df42e3f81c634['h017fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c00] =  I0310077d53ae4ed9904df42e3f81c634['h01800] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c01] =  I0310077d53ae4ed9904df42e3f81c634['h01802] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c02] =  I0310077d53ae4ed9904df42e3f81c634['h01804] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c03] =  I0310077d53ae4ed9904df42e3f81c634['h01806] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c04] =  I0310077d53ae4ed9904df42e3f81c634['h01808] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c05] =  I0310077d53ae4ed9904df42e3f81c634['h0180a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c06] =  I0310077d53ae4ed9904df42e3f81c634['h0180c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c07] =  I0310077d53ae4ed9904df42e3f81c634['h0180e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c08] =  I0310077d53ae4ed9904df42e3f81c634['h01810] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c09] =  I0310077d53ae4ed9904df42e3f81c634['h01812] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c0a] =  I0310077d53ae4ed9904df42e3f81c634['h01814] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c0b] =  I0310077d53ae4ed9904df42e3f81c634['h01816] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c0c] =  I0310077d53ae4ed9904df42e3f81c634['h01818] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c0d] =  I0310077d53ae4ed9904df42e3f81c634['h0181a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c0e] =  I0310077d53ae4ed9904df42e3f81c634['h0181c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c0f] =  I0310077d53ae4ed9904df42e3f81c634['h0181e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c10] =  I0310077d53ae4ed9904df42e3f81c634['h01820] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c11] =  I0310077d53ae4ed9904df42e3f81c634['h01822] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c12] =  I0310077d53ae4ed9904df42e3f81c634['h01824] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c13] =  I0310077d53ae4ed9904df42e3f81c634['h01826] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c14] =  I0310077d53ae4ed9904df42e3f81c634['h01828] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c15] =  I0310077d53ae4ed9904df42e3f81c634['h0182a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c16] =  I0310077d53ae4ed9904df42e3f81c634['h0182c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c17] =  I0310077d53ae4ed9904df42e3f81c634['h0182e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c18] =  I0310077d53ae4ed9904df42e3f81c634['h01830] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c19] =  I0310077d53ae4ed9904df42e3f81c634['h01832] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c1a] =  I0310077d53ae4ed9904df42e3f81c634['h01834] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c1b] =  I0310077d53ae4ed9904df42e3f81c634['h01836] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c1c] =  I0310077d53ae4ed9904df42e3f81c634['h01838] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c1d] =  I0310077d53ae4ed9904df42e3f81c634['h0183a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c1e] =  I0310077d53ae4ed9904df42e3f81c634['h0183c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c1f] =  I0310077d53ae4ed9904df42e3f81c634['h0183e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c20] =  I0310077d53ae4ed9904df42e3f81c634['h01840] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c21] =  I0310077d53ae4ed9904df42e3f81c634['h01842] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c22] =  I0310077d53ae4ed9904df42e3f81c634['h01844] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c23] =  I0310077d53ae4ed9904df42e3f81c634['h01846] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c24] =  I0310077d53ae4ed9904df42e3f81c634['h01848] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c25] =  I0310077d53ae4ed9904df42e3f81c634['h0184a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c26] =  I0310077d53ae4ed9904df42e3f81c634['h0184c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c27] =  I0310077d53ae4ed9904df42e3f81c634['h0184e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c28] =  I0310077d53ae4ed9904df42e3f81c634['h01850] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c29] =  I0310077d53ae4ed9904df42e3f81c634['h01852] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c2a] =  I0310077d53ae4ed9904df42e3f81c634['h01854] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c2b] =  I0310077d53ae4ed9904df42e3f81c634['h01856] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c2c] =  I0310077d53ae4ed9904df42e3f81c634['h01858] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c2d] =  I0310077d53ae4ed9904df42e3f81c634['h0185a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c2e] =  I0310077d53ae4ed9904df42e3f81c634['h0185c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c2f] =  I0310077d53ae4ed9904df42e3f81c634['h0185e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c30] =  I0310077d53ae4ed9904df42e3f81c634['h01860] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c31] =  I0310077d53ae4ed9904df42e3f81c634['h01862] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c32] =  I0310077d53ae4ed9904df42e3f81c634['h01864] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c33] =  I0310077d53ae4ed9904df42e3f81c634['h01866] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c34] =  I0310077d53ae4ed9904df42e3f81c634['h01868] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c35] =  I0310077d53ae4ed9904df42e3f81c634['h0186a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c36] =  I0310077d53ae4ed9904df42e3f81c634['h0186c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c37] =  I0310077d53ae4ed9904df42e3f81c634['h0186e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c38] =  I0310077d53ae4ed9904df42e3f81c634['h01870] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c39] =  I0310077d53ae4ed9904df42e3f81c634['h01872] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c3a] =  I0310077d53ae4ed9904df42e3f81c634['h01874] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c3b] =  I0310077d53ae4ed9904df42e3f81c634['h01876] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c3c] =  I0310077d53ae4ed9904df42e3f81c634['h01878] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c3d] =  I0310077d53ae4ed9904df42e3f81c634['h0187a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c3e] =  I0310077d53ae4ed9904df42e3f81c634['h0187c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c3f] =  I0310077d53ae4ed9904df42e3f81c634['h0187e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c40] =  I0310077d53ae4ed9904df42e3f81c634['h01880] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c41] =  I0310077d53ae4ed9904df42e3f81c634['h01882] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c42] =  I0310077d53ae4ed9904df42e3f81c634['h01884] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c43] =  I0310077d53ae4ed9904df42e3f81c634['h01886] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c44] =  I0310077d53ae4ed9904df42e3f81c634['h01888] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c45] =  I0310077d53ae4ed9904df42e3f81c634['h0188a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c46] =  I0310077d53ae4ed9904df42e3f81c634['h0188c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c47] =  I0310077d53ae4ed9904df42e3f81c634['h0188e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c48] =  I0310077d53ae4ed9904df42e3f81c634['h01890] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c49] =  I0310077d53ae4ed9904df42e3f81c634['h01892] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c4a] =  I0310077d53ae4ed9904df42e3f81c634['h01894] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c4b] =  I0310077d53ae4ed9904df42e3f81c634['h01896] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c4c] =  I0310077d53ae4ed9904df42e3f81c634['h01898] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c4d] =  I0310077d53ae4ed9904df42e3f81c634['h0189a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c4e] =  I0310077d53ae4ed9904df42e3f81c634['h0189c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c4f] =  I0310077d53ae4ed9904df42e3f81c634['h0189e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c50] =  I0310077d53ae4ed9904df42e3f81c634['h018a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c51] =  I0310077d53ae4ed9904df42e3f81c634['h018a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c52] =  I0310077d53ae4ed9904df42e3f81c634['h018a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c53] =  I0310077d53ae4ed9904df42e3f81c634['h018a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c54] =  I0310077d53ae4ed9904df42e3f81c634['h018a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c55] =  I0310077d53ae4ed9904df42e3f81c634['h018aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c56] =  I0310077d53ae4ed9904df42e3f81c634['h018ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c57] =  I0310077d53ae4ed9904df42e3f81c634['h018ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c58] =  I0310077d53ae4ed9904df42e3f81c634['h018b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c59] =  I0310077d53ae4ed9904df42e3f81c634['h018b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c5a] =  I0310077d53ae4ed9904df42e3f81c634['h018b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c5b] =  I0310077d53ae4ed9904df42e3f81c634['h018b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c5c] =  I0310077d53ae4ed9904df42e3f81c634['h018b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c5d] =  I0310077d53ae4ed9904df42e3f81c634['h018ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c5e] =  I0310077d53ae4ed9904df42e3f81c634['h018bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c5f] =  I0310077d53ae4ed9904df42e3f81c634['h018be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c60] =  I0310077d53ae4ed9904df42e3f81c634['h018c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c61] =  I0310077d53ae4ed9904df42e3f81c634['h018c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c62] =  I0310077d53ae4ed9904df42e3f81c634['h018c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c63] =  I0310077d53ae4ed9904df42e3f81c634['h018c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c64] =  I0310077d53ae4ed9904df42e3f81c634['h018c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c65] =  I0310077d53ae4ed9904df42e3f81c634['h018ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c66] =  I0310077d53ae4ed9904df42e3f81c634['h018cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c67] =  I0310077d53ae4ed9904df42e3f81c634['h018ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c68] =  I0310077d53ae4ed9904df42e3f81c634['h018d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c69] =  I0310077d53ae4ed9904df42e3f81c634['h018d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c6a] =  I0310077d53ae4ed9904df42e3f81c634['h018d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c6b] =  I0310077d53ae4ed9904df42e3f81c634['h018d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c6c] =  I0310077d53ae4ed9904df42e3f81c634['h018d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c6d] =  I0310077d53ae4ed9904df42e3f81c634['h018da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c6e] =  I0310077d53ae4ed9904df42e3f81c634['h018dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c6f] =  I0310077d53ae4ed9904df42e3f81c634['h018de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c70] =  I0310077d53ae4ed9904df42e3f81c634['h018e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c71] =  I0310077d53ae4ed9904df42e3f81c634['h018e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c72] =  I0310077d53ae4ed9904df42e3f81c634['h018e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c73] =  I0310077d53ae4ed9904df42e3f81c634['h018e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c74] =  I0310077d53ae4ed9904df42e3f81c634['h018e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c75] =  I0310077d53ae4ed9904df42e3f81c634['h018ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c76] =  I0310077d53ae4ed9904df42e3f81c634['h018ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c77] =  I0310077d53ae4ed9904df42e3f81c634['h018ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c78] =  I0310077d53ae4ed9904df42e3f81c634['h018f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c79] =  I0310077d53ae4ed9904df42e3f81c634['h018f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c7a] =  I0310077d53ae4ed9904df42e3f81c634['h018f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c7b] =  I0310077d53ae4ed9904df42e3f81c634['h018f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c7c] =  I0310077d53ae4ed9904df42e3f81c634['h018f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c7d] =  I0310077d53ae4ed9904df42e3f81c634['h018fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c7e] =  I0310077d53ae4ed9904df42e3f81c634['h018fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c7f] =  I0310077d53ae4ed9904df42e3f81c634['h018fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c80] =  I0310077d53ae4ed9904df42e3f81c634['h01900] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c81] =  I0310077d53ae4ed9904df42e3f81c634['h01902] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c82] =  I0310077d53ae4ed9904df42e3f81c634['h01904] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c83] =  I0310077d53ae4ed9904df42e3f81c634['h01906] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c84] =  I0310077d53ae4ed9904df42e3f81c634['h01908] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c85] =  I0310077d53ae4ed9904df42e3f81c634['h0190a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c86] =  I0310077d53ae4ed9904df42e3f81c634['h0190c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c87] =  I0310077d53ae4ed9904df42e3f81c634['h0190e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c88] =  I0310077d53ae4ed9904df42e3f81c634['h01910] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c89] =  I0310077d53ae4ed9904df42e3f81c634['h01912] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c8a] =  I0310077d53ae4ed9904df42e3f81c634['h01914] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c8b] =  I0310077d53ae4ed9904df42e3f81c634['h01916] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c8c] =  I0310077d53ae4ed9904df42e3f81c634['h01918] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c8d] =  I0310077d53ae4ed9904df42e3f81c634['h0191a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c8e] =  I0310077d53ae4ed9904df42e3f81c634['h0191c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c8f] =  I0310077d53ae4ed9904df42e3f81c634['h0191e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c90] =  I0310077d53ae4ed9904df42e3f81c634['h01920] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c91] =  I0310077d53ae4ed9904df42e3f81c634['h01922] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c92] =  I0310077d53ae4ed9904df42e3f81c634['h01924] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c93] =  I0310077d53ae4ed9904df42e3f81c634['h01926] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c94] =  I0310077d53ae4ed9904df42e3f81c634['h01928] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c95] =  I0310077d53ae4ed9904df42e3f81c634['h0192a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c96] =  I0310077d53ae4ed9904df42e3f81c634['h0192c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c97] =  I0310077d53ae4ed9904df42e3f81c634['h0192e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c98] =  I0310077d53ae4ed9904df42e3f81c634['h01930] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c99] =  I0310077d53ae4ed9904df42e3f81c634['h01932] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c9a] =  I0310077d53ae4ed9904df42e3f81c634['h01934] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c9b] =  I0310077d53ae4ed9904df42e3f81c634['h01936] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c9c] =  I0310077d53ae4ed9904df42e3f81c634['h01938] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c9d] =  I0310077d53ae4ed9904df42e3f81c634['h0193a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c9e] =  I0310077d53ae4ed9904df42e3f81c634['h0193c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00c9f] =  I0310077d53ae4ed9904df42e3f81c634['h0193e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca0] =  I0310077d53ae4ed9904df42e3f81c634['h01940] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca1] =  I0310077d53ae4ed9904df42e3f81c634['h01942] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca2] =  I0310077d53ae4ed9904df42e3f81c634['h01944] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca3] =  I0310077d53ae4ed9904df42e3f81c634['h01946] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca4] =  I0310077d53ae4ed9904df42e3f81c634['h01948] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca5] =  I0310077d53ae4ed9904df42e3f81c634['h0194a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca6] =  I0310077d53ae4ed9904df42e3f81c634['h0194c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca7] =  I0310077d53ae4ed9904df42e3f81c634['h0194e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca8] =  I0310077d53ae4ed9904df42e3f81c634['h01950] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ca9] =  I0310077d53ae4ed9904df42e3f81c634['h01952] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00caa] =  I0310077d53ae4ed9904df42e3f81c634['h01954] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cab] =  I0310077d53ae4ed9904df42e3f81c634['h01956] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cac] =  I0310077d53ae4ed9904df42e3f81c634['h01958] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cad] =  I0310077d53ae4ed9904df42e3f81c634['h0195a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cae] =  I0310077d53ae4ed9904df42e3f81c634['h0195c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00caf] =  I0310077d53ae4ed9904df42e3f81c634['h0195e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb0] =  I0310077d53ae4ed9904df42e3f81c634['h01960] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb1] =  I0310077d53ae4ed9904df42e3f81c634['h01962] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb2] =  I0310077d53ae4ed9904df42e3f81c634['h01964] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb3] =  I0310077d53ae4ed9904df42e3f81c634['h01966] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb4] =  I0310077d53ae4ed9904df42e3f81c634['h01968] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb5] =  I0310077d53ae4ed9904df42e3f81c634['h0196a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb6] =  I0310077d53ae4ed9904df42e3f81c634['h0196c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb7] =  I0310077d53ae4ed9904df42e3f81c634['h0196e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb8] =  I0310077d53ae4ed9904df42e3f81c634['h01970] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cb9] =  I0310077d53ae4ed9904df42e3f81c634['h01972] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cba] =  I0310077d53ae4ed9904df42e3f81c634['h01974] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cbb] =  I0310077d53ae4ed9904df42e3f81c634['h01976] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cbc] =  I0310077d53ae4ed9904df42e3f81c634['h01978] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cbd] =  I0310077d53ae4ed9904df42e3f81c634['h0197a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cbe] =  I0310077d53ae4ed9904df42e3f81c634['h0197c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cbf] =  I0310077d53ae4ed9904df42e3f81c634['h0197e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc0] =  I0310077d53ae4ed9904df42e3f81c634['h01980] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc1] =  I0310077d53ae4ed9904df42e3f81c634['h01982] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc2] =  I0310077d53ae4ed9904df42e3f81c634['h01984] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc3] =  I0310077d53ae4ed9904df42e3f81c634['h01986] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc4] =  I0310077d53ae4ed9904df42e3f81c634['h01988] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc5] =  I0310077d53ae4ed9904df42e3f81c634['h0198a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc6] =  I0310077d53ae4ed9904df42e3f81c634['h0198c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc7] =  I0310077d53ae4ed9904df42e3f81c634['h0198e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc8] =  I0310077d53ae4ed9904df42e3f81c634['h01990] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cc9] =  I0310077d53ae4ed9904df42e3f81c634['h01992] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cca] =  I0310077d53ae4ed9904df42e3f81c634['h01994] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ccb] =  I0310077d53ae4ed9904df42e3f81c634['h01996] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ccc] =  I0310077d53ae4ed9904df42e3f81c634['h01998] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ccd] =  I0310077d53ae4ed9904df42e3f81c634['h0199a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cce] =  I0310077d53ae4ed9904df42e3f81c634['h0199c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ccf] =  I0310077d53ae4ed9904df42e3f81c634['h0199e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd0] =  I0310077d53ae4ed9904df42e3f81c634['h019a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd1] =  I0310077d53ae4ed9904df42e3f81c634['h019a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd2] =  I0310077d53ae4ed9904df42e3f81c634['h019a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd3] =  I0310077d53ae4ed9904df42e3f81c634['h019a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd4] =  I0310077d53ae4ed9904df42e3f81c634['h019a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd5] =  I0310077d53ae4ed9904df42e3f81c634['h019aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd6] =  I0310077d53ae4ed9904df42e3f81c634['h019ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd7] =  I0310077d53ae4ed9904df42e3f81c634['h019ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd8] =  I0310077d53ae4ed9904df42e3f81c634['h019b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cd9] =  I0310077d53ae4ed9904df42e3f81c634['h019b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cda] =  I0310077d53ae4ed9904df42e3f81c634['h019b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cdb] =  I0310077d53ae4ed9904df42e3f81c634['h019b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cdc] =  I0310077d53ae4ed9904df42e3f81c634['h019b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cdd] =  I0310077d53ae4ed9904df42e3f81c634['h019ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cde] =  I0310077d53ae4ed9904df42e3f81c634['h019bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cdf] =  I0310077d53ae4ed9904df42e3f81c634['h019be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce0] =  I0310077d53ae4ed9904df42e3f81c634['h019c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce1] =  I0310077d53ae4ed9904df42e3f81c634['h019c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce2] =  I0310077d53ae4ed9904df42e3f81c634['h019c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce3] =  I0310077d53ae4ed9904df42e3f81c634['h019c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce4] =  I0310077d53ae4ed9904df42e3f81c634['h019c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce5] =  I0310077d53ae4ed9904df42e3f81c634['h019ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce6] =  I0310077d53ae4ed9904df42e3f81c634['h019cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce7] =  I0310077d53ae4ed9904df42e3f81c634['h019ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce8] =  I0310077d53ae4ed9904df42e3f81c634['h019d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ce9] =  I0310077d53ae4ed9904df42e3f81c634['h019d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cea] =  I0310077d53ae4ed9904df42e3f81c634['h019d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ceb] =  I0310077d53ae4ed9904df42e3f81c634['h019d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cec] =  I0310077d53ae4ed9904df42e3f81c634['h019d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ced] =  I0310077d53ae4ed9904df42e3f81c634['h019da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cee] =  I0310077d53ae4ed9904df42e3f81c634['h019dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cef] =  I0310077d53ae4ed9904df42e3f81c634['h019de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf0] =  I0310077d53ae4ed9904df42e3f81c634['h019e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf1] =  I0310077d53ae4ed9904df42e3f81c634['h019e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf2] =  I0310077d53ae4ed9904df42e3f81c634['h019e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf3] =  I0310077d53ae4ed9904df42e3f81c634['h019e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf4] =  I0310077d53ae4ed9904df42e3f81c634['h019e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf5] =  I0310077d53ae4ed9904df42e3f81c634['h019ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf6] =  I0310077d53ae4ed9904df42e3f81c634['h019ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf7] =  I0310077d53ae4ed9904df42e3f81c634['h019ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf8] =  I0310077d53ae4ed9904df42e3f81c634['h019f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cf9] =  I0310077d53ae4ed9904df42e3f81c634['h019f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cfa] =  I0310077d53ae4ed9904df42e3f81c634['h019f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cfb] =  I0310077d53ae4ed9904df42e3f81c634['h019f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cfc] =  I0310077d53ae4ed9904df42e3f81c634['h019f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cfd] =  I0310077d53ae4ed9904df42e3f81c634['h019fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cfe] =  I0310077d53ae4ed9904df42e3f81c634['h019fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00cff] =  I0310077d53ae4ed9904df42e3f81c634['h019fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d00] =  I0310077d53ae4ed9904df42e3f81c634['h01a00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d01] =  I0310077d53ae4ed9904df42e3f81c634['h01a02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d02] =  I0310077d53ae4ed9904df42e3f81c634['h01a04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d03] =  I0310077d53ae4ed9904df42e3f81c634['h01a06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d04] =  I0310077d53ae4ed9904df42e3f81c634['h01a08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d05] =  I0310077d53ae4ed9904df42e3f81c634['h01a0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d06] =  I0310077d53ae4ed9904df42e3f81c634['h01a0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d07] =  I0310077d53ae4ed9904df42e3f81c634['h01a0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d08] =  I0310077d53ae4ed9904df42e3f81c634['h01a10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d09] =  I0310077d53ae4ed9904df42e3f81c634['h01a12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d0a] =  I0310077d53ae4ed9904df42e3f81c634['h01a14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d0b] =  I0310077d53ae4ed9904df42e3f81c634['h01a16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d0c] =  I0310077d53ae4ed9904df42e3f81c634['h01a18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d0d] =  I0310077d53ae4ed9904df42e3f81c634['h01a1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d0e] =  I0310077d53ae4ed9904df42e3f81c634['h01a1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d0f] =  I0310077d53ae4ed9904df42e3f81c634['h01a1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d10] =  I0310077d53ae4ed9904df42e3f81c634['h01a20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d11] =  I0310077d53ae4ed9904df42e3f81c634['h01a22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d12] =  I0310077d53ae4ed9904df42e3f81c634['h01a24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d13] =  I0310077d53ae4ed9904df42e3f81c634['h01a26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d14] =  I0310077d53ae4ed9904df42e3f81c634['h01a28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d15] =  I0310077d53ae4ed9904df42e3f81c634['h01a2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d16] =  I0310077d53ae4ed9904df42e3f81c634['h01a2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d17] =  I0310077d53ae4ed9904df42e3f81c634['h01a2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d18] =  I0310077d53ae4ed9904df42e3f81c634['h01a30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d19] =  I0310077d53ae4ed9904df42e3f81c634['h01a32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d1a] =  I0310077d53ae4ed9904df42e3f81c634['h01a34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d1b] =  I0310077d53ae4ed9904df42e3f81c634['h01a36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d1c] =  I0310077d53ae4ed9904df42e3f81c634['h01a38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d1d] =  I0310077d53ae4ed9904df42e3f81c634['h01a3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d1e] =  I0310077d53ae4ed9904df42e3f81c634['h01a3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d1f] =  I0310077d53ae4ed9904df42e3f81c634['h01a3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d20] =  I0310077d53ae4ed9904df42e3f81c634['h01a40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d21] =  I0310077d53ae4ed9904df42e3f81c634['h01a42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d22] =  I0310077d53ae4ed9904df42e3f81c634['h01a44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d23] =  I0310077d53ae4ed9904df42e3f81c634['h01a46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d24] =  I0310077d53ae4ed9904df42e3f81c634['h01a48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d25] =  I0310077d53ae4ed9904df42e3f81c634['h01a4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d26] =  I0310077d53ae4ed9904df42e3f81c634['h01a4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d27] =  I0310077d53ae4ed9904df42e3f81c634['h01a4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d28] =  I0310077d53ae4ed9904df42e3f81c634['h01a50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d29] =  I0310077d53ae4ed9904df42e3f81c634['h01a52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d2a] =  I0310077d53ae4ed9904df42e3f81c634['h01a54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d2b] =  I0310077d53ae4ed9904df42e3f81c634['h01a56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d2c] =  I0310077d53ae4ed9904df42e3f81c634['h01a58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d2d] =  I0310077d53ae4ed9904df42e3f81c634['h01a5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d2e] =  I0310077d53ae4ed9904df42e3f81c634['h01a5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d2f] =  I0310077d53ae4ed9904df42e3f81c634['h01a5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d30] =  I0310077d53ae4ed9904df42e3f81c634['h01a60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d31] =  I0310077d53ae4ed9904df42e3f81c634['h01a62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d32] =  I0310077d53ae4ed9904df42e3f81c634['h01a64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d33] =  I0310077d53ae4ed9904df42e3f81c634['h01a66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d34] =  I0310077d53ae4ed9904df42e3f81c634['h01a68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d35] =  I0310077d53ae4ed9904df42e3f81c634['h01a6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d36] =  I0310077d53ae4ed9904df42e3f81c634['h01a6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d37] =  I0310077d53ae4ed9904df42e3f81c634['h01a6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d38] =  I0310077d53ae4ed9904df42e3f81c634['h01a70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d39] =  I0310077d53ae4ed9904df42e3f81c634['h01a72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d3a] =  I0310077d53ae4ed9904df42e3f81c634['h01a74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d3b] =  I0310077d53ae4ed9904df42e3f81c634['h01a76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d3c] =  I0310077d53ae4ed9904df42e3f81c634['h01a78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d3d] =  I0310077d53ae4ed9904df42e3f81c634['h01a7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d3e] =  I0310077d53ae4ed9904df42e3f81c634['h01a7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d3f] =  I0310077d53ae4ed9904df42e3f81c634['h01a7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d40] =  I0310077d53ae4ed9904df42e3f81c634['h01a80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d41] =  I0310077d53ae4ed9904df42e3f81c634['h01a82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d42] =  I0310077d53ae4ed9904df42e3f81c634['h01a84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d43] =  I0310077d53ae4ed9904df42e3f81c634['h01a86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d44] =  I0310077d53ae4ed9904df42e3f81c634['h01a88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d45] =  I0310077d53ae4ed9904df42e3f81c634['h01a8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d46] =  I0310077d53ae4ed9904df42e3f81c634['h01a8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d47] =  I0310077d53ae4ed9904df42e3f81c634['h01a8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d48] =  I0310077d53ae4ed9904df42e3f81c634['h01a90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d49] =  I0310077d53ae4ed9904df42e3f81c634['h01a92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d4a] =  I0310077d53ae4ed9904df42e3f81c634['h01a94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d4b] =  I0310077d53ae4ed9904df42e3f81c634['h01a96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d4c] =  I0310077d53ae4ed9904df42e3f81c634['h01a98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d4d] =  I0310077d53ae4ed9904df42e3f81c634['h01a9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d4e] =  I0310077d53ae4ed9904df42e3f81c634['h01a9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d4f] =  I0310077d53ae4ed9904df42e3f81c634['h01a9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d50] =  I0310077d53ae4ed9904df42e3f81c634['h01aa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d51] =  I0310077d53ae4ed9904df42e3f81c634['h01aa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d52] =  I0310077d53ae4ed9904df42e3f81c634['h01aa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d53] =  I0310077d53ae4ed9904df42e3f81c634['h01aa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d54] =  I0310077d53ae4ed9904df42e3f81c634['h01aa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d55] =  I0310077d53ae4ed9904df42e3f81c634['h01aaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d56] =  I0310077d53ae4ed9904df42e3f81c634['h01aac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d57] =  I0310077d53ae4ed9904df42e3f81c634['h01aae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d58] =  I0310077d53ae4ed9904df42e3f81c634['h01ab0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d59] =  I0310077d53ae4ed9904df42e3f81c634['h01ab2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d5a] =  I0310077d53ae4ed9904df42e3f81c634['h01ab4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d5b] =  I0310077d53ae4ed9904df42e3f81c634['h01ab6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d5c] =  I0310077d53ae4ed9904df42e3f81c634['h01ab8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d5d] =  I0310077d53ae4ed9904df42e3f81c634['h01aba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d5e] =  I0310077d53ae4ed9904df42e3f81c634['h01abc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d5f] =  I0310077d53ae4ed9904df42e3f81c634['h01abe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d60] =  I0310077d53ae4ed9904df42e3f81c634['h01ac0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d61] =  I0310077d53ae4ed9904df42e3f81c634['h01ac2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d62] =  I0310077d53ae4ed9904df42e3f81c634['h01ac4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d63] =  I0310077d53ae4ed9904df42e3f81c634['h01ac6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d64] =  I0310077d53ae4ed9904df42e3f81c634['h01ac8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d65] =  I0310077d53ae4ed9904df42e3f81c634['h01aca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d66] =  I0310077d53ae4ed9904df42e3f81c634['h01acc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d67] =  I0310077d53ae4ed9904df42e3f81c634['h01ace] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d68] =  I0310077d53ae4ed9904df42e3f81c634['h01ad0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d69] =  I0310077d53ae4ed9904df42e3f81c634['h01ad2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d6a] =  I0310077d53ae4ed9904df42e3f81c634['h01ad4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d6b] =  I0310077d53ae4ed9904df42e3f81c634['h01ad6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d6c] =  I0310077d53ae4ed9904df42e3f81c634['h01ad8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d6d] =  I0310077d53ae4ed9904df42e3f81c634['h01ada] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d6e] =  I0310077d53ae4ed9904df42e3f81c634['h01adc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d6f] =  I0310077d53ae4ed9904df42e3f81c634['h01ade] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d70] =  I0310077d53ae4ed9904df42e3f81c634['h01ae0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d71] =  I0310077d53ae4ed9904df42e3f81c634['h01ae2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d72] =  I0310077d53ae4ed9904df42e3f81c634['h01ae4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d73] =  I0310077d53ae4ed9904df42e3f81c634['h01ae6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d74] =  I0310077d53ae4ed9904df42e3f81c634['h01ae8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d75] =  I0310077d53ae4ed9904df42e3f81c634['h01aea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d76] =  I0310077d53ae4ed9904df42e3f81c634['h01aec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d77] =  I0310077d53ae4ed9904df42e3f81c634['h01aee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d78] =  I0310077d53ae4ed9904df42e3f81c634['h01af0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d79] =  I0310077d53ae4ed9904df42e3f81c634['h01af2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d7a] =  I0310077d53ae4ed9904df42e3f81c634['h01af4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d7b] =  I0310077d53ae4ed9904df42e3f81c634['h01af6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d7c] =  I0310077d53ae4ed9904df42e3f81c634['h01af8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d7d] =  I0310077d53ae4ed9904df42e3f81c634['h01afa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d7e] =  I0310077d53ae4ed9904df42e3f81c634['h01afc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d7f] =  I0310077d53ae4ed9904df42e3f81c634['h01afe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d80] =  I0310077d53ae4ed9904df42e3f81c634['h01b00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d81] =  I0310077d53ae4ed9904df42e3f81c634['h01b02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d82] =  I0310077d53ae4ed9904df42e3f81c634['h01b04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d83] =  I0310077d53ae4ed9904df42e3f81c634['h01b06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d84] =  I0310077d53ae4ed9904df42e3f81c634['h01b08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d85] =  I0310077d53ae4ed9904df42e3f81c634['h01b0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d86] =  I0310077d53ae4ed9904df42e3f81c634['h01b0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d87] =  I0310077d53ae4ed9904df42e3f81c634['h01b0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d88] =  I0310077d53ae4ed9904df42e3f81c634['h01b10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d89] =  I0310077d53ae4ed9904df42e3f81c634['h01b12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d8a] =  I0310077d53ae4ed9904df42e3f81c634['h01b14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d8b] =  I0310077d53ae4ed9904df42e3f81c634['h01b16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d8c] =  I0310077d53ae4ed9904df42e3f81c634['h01b18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d8d] =  I0310077d53ae4ed9904df42e3f81c634['h01b1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d8e] =  I0310077d53ae4ed9904df42e3f81c634['h01b1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d8f] =  I0310077d53ae4ed9904df42e3f81c634['h01b1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d90] =  I0310077d53ae4ed9904df42e3f81c634['h01b20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d91] =  I0310077d53ae4ed9904df42e3f81c634['h01b22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d92] =  I0310077d53ae4ed9904df42e3f81c634['h01b24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d93] =  I0310077d53ae4ed9904df42e3f81c634['h01b26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d94] =  I0310077d53ae4ed9904df42e3f81c634['h01b28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d95] =  I0310077d53ae4ed9904df42e3f81c634['h01b2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d96] =  I0310077d53ae4ed9904df42e3f81c634['h01b2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d97] =  I0310077d53ae4ed9904df42e3f81c634['h01b2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d98] =  I0310077d53ae4ed9904df42e3f81c634['h01b30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d99] =  I0310077d53ae4ed9904df42e3f81c634['h01b32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d9a] =  I0310077d53ae4ed9904df42e3f81c634['h01b34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d9b] =  I0310077d53ae4ed9904df42e3f81c634['h01b36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d9c] =  I0310077d53ae4ed9904df42e3f81c634['h01b38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d9d] =  I0310077d53ae4ed9904df42e3f81c634['h01b3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d9e] =  I0310077d53ae4ed9904df42e3f81c634['h01b3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00d9f] =  I0310077d53ae4ed9904df42e3f81c634['h01b3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da0] =  I0310077d53ae4ed9904df42e3f81c634['h01b40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da1] =  I0310077d53ae4ed9904df42e3f81c634['h01b42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da2] =  I0310077d53ae4ed9904df42e3f81c634['h01b44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da3] =  I0310077d53ae4ed9904df42e3f81c634['h01b46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da4] =  I0310077d53ae4ed9904df42e3f81c634['h01b48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da5] =  I0310077d53ae4ed9904df42e3f81c634['h01b4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da6] =  I0310077d53ae4ed9904df42e3f81c634['h01b4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da7] =  I0310077d53ae4ed9904df42e3f81c634['h01b4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da8] =  I0310077d53ae4ed9904df42e3f81c634['h01b50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00da9] =  I0310077d53ae4ed9904df42e3f81c634['h01b52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00daa] =  I0310077d53ae4ed9904df42e3f81c634['h01b54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dab] =  I0310077d53ae4ed9904df42e3f81c634['h01b56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dac] =  I0310077d53ae4ed9904df42e3f81c634['h01b58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dad] =  I0310077d53ae4ed9904df42e3f81c634['h01b5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dae] =  I0310077d53ae4ed9904df42e3f81c634['h01b5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00daf] =  I0310077d53ae4ed9904df42e3f81c634['h01b5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db0] =  I0310077d53ae4ed9904df42e3f81c634['h01b60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db1] =  I0310077d53ae4ed9904df42e3f81c634['h01b62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db2] =  I0310077d53ae4ed9904df42e3f81c634['h01b64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db3] =  I0310077d53ae4ed9904df42e3f81c634['h01b66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db4] =  I0310077d53ae4ed9904df42e3f81c634['h01b68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db5] =  I0310077d53ae4ed9904df42e3f81c634['h01b6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db6] =  I0310077d53ae4ed9904df42e3f81c634['h01b6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db7] =  I0310077d53ae4ed9904df42e3f81c634['h01b6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db8] =  I0310077d53ae4ed9904df42e3f81c634['h01b70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00db9] =  I0310077d53ae4ed9904df42e3f81c634['h01b72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dba] =  I0310077d53ae4ed9904df42e3f81c634['h01b74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dbb] =  I0310077d53ae4ed9904df42e3f81c634['h01b76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dbc] =  I0310077d53ae4ed9904df42e3f81c634['h01b78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dbd] =  I0310077d53ae4ed9904df42e3f81c634['h01b7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dbe] =  I0310077d53ae4ed9904df42e3f81c634['h01b7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dbf] =  I0310077d53ae4ed9904df42e3f81c634['h01b7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc0] =  I0310077d53ae4ed9904df42e3f81c634['h01b80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc1] =  I0310077d53ae4ed9904df42e3f81c634['h01b82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc2] =  I0310077d53ae4ed9904df42e3f81c634['h01b84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc3] =  I0310077d53ae4ed9904df42e3f81c634['h01b86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc4] =  I0310077d53ae4ed9904df42e3f81c634['h01b88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc5] =  I0310077d53ae4ed9904df42e3f81c634['h01b8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc6] =  I0310077d53ae4ed9904df42e3f81c634['h01b8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc7] =  I0310077d53ae4ed9904df42e3f81c634['h01b8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc8] =  I0310077d53ae4ed9904df42e3f81c634['h01b90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dc9] =  I0310077d53ae4ed9904df42e3f81c634['h01b92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dca] =  I0310077d53ae4ed9904df42e3f81c634['h01b94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dcb] =  I0310077d53ae4ed9904df42e3f81c634['h01b96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dcc] =  I0310077d53ae4ed9904df42e3f81c634['h01b98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dcd] =  I0310077d53ae4ed9904df42e3f81c634['h01b9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dce] =  I0310077d53ae4ed9904df42e3f81c634['h01b9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dcf] =  I0310077d53ae4ed9904df42e3f81c634['h01b9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd0] =  I0310077d53ae4ed9904df42e3f81c634['h01ba0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd1] =  I0310077d53ae4ed9904df42e3f81c634['h01ba2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd2] =  I0310077d53ae4ed9904df42e3f81c634['h01ba4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd3] =  I0310077d53ae4ed9904df42e3f81c634['h01ba6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd4] =  I0310077d53ae4ed9904df42e3f81c634['h01ba8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd5] =  I0310077d53ae4ed9904df42e3f81c634['h01baa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd6] =  I0310077d53ae4ed9904df42e3f81c634['h01bac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd7] =  I0310077d53ae4ed9904df42e3f81c634['h01bae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd8] =  I0310077d53ae4ed9904df42e3f81c634['h01bb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dd9] =  I0310077d53ae4ed9904df42e3f81c634['h01bb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dda] =  I0310077d53ae4ed9904df42e3f81c634['h01bb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ddb] =  I0310077d53ae4ed9904df42e3f81c634['h01bb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ddc] =  I0310077d53ae4ed9904df42e3f81c634['h01bb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ddd] =  I0310077d53ae4ed9904df42e3f81c634['h01bba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dde] =  I0310077d53ae4ed9904df42e3f81c634['h01bbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ddf] =  I0310077d53ae4ed9904df42e3f81c634['h01bbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de0] =  I0310077d53ae4ed9904df42e3f81c634['h01bc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de1] =  I0310077d53ae4ed9904df42e3f81c634['h01bc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de2] =  I0310077d53ae4ed9904df42e3f81c634['h01bc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de3] =  I0310077d53ae4ed9904df42e3f81c634['h01bc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de4] =  I0310077d53ae4ed9904df42e3f81c634['h01bc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de5] =  I0310077d53ae4ed9904df42e3f81c634['h01bca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de6] =  I0310077d53ae4ed9904df42e3f81c634['h01bcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de7] =  I0310077d53ae4ed9904df42e3f81c634['h01bce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de8] =  I0310077d53ae4ed9904df42e3f81c634['h01bd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00de9] =  I0310077d53ae4ed9904df42e3f81c634['h01bd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dea] =  I0310077d53ae4ed9904df42e3f81c634['h01bd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00deb] =  I0310077d53ae4ed9904df42e3f81c634['h01bd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dec] =  I0310077d53ae4ed9904df42e3f81c634['h01bd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ded] =  I0310077d53ae4ed9904df42e3f81c634['h01bda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dee] =  I0310077d53ae4ed9904df42e3f81c634['h01bdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00def] =  I0310077d53ae4ed9904df42e3f81c634['h01bde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df0] =  I0310077d53ae4ed9904df42e3f81c634['h01be0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df1] =  I0310077d53ae4ed9904df42e3f81c634['h01be2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df2] =  I0310077d53ae4ed9904df42e3f81c634['h01be4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df3] =  I0310077d53ae4ed9904df42e3f81c634['h01be6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df4] =  I0310077d53ae4ed9904df42e3f81c634['h01be8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df5] =  I0310077d53ae4ed9904df42e3f81c634['h01bea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df6] =  I0310077d53ae4ed9904df42e3f81c634['h01bec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df7] =  I0310077d53ae4ed9904df42e3f81c634['h01bee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df8] =  I0310077d53ae4ed9904df42e3f81c634['h01bf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00df9] =  I0310077d53ae4ed9904df42e3f81c634['h01bf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dfa] =  I0310077d53ae4ed9904df42e3f81c634['h01bf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dfb] =  I0310077d53ae4ed9904df42e3f81c634['h01bf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dfc] =  I0310077d53ae4ed9904df42e3f81c634['h01bf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dfd] =  I0310077d53ae4ed9904df42e3f81c634['h01bfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dfe] =  I0310077d53ae4ed9904df42e3f81c634['h01bfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00dff] =  I0310077d53ae4ed9904df42e3f81c634['h01bfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e00] =  I0310077d53ae4ed9904df42e3f81c634['h01c00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e01] =  I0310077d53ae4ed9904df42e3f81c634['h01c02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e02] =  I0310077d53ae4ed9904df42e3f81c634['h01c04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e03] =  I0310077d53ae4ed9904df42e3f81c634['h01c06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e04] =  I0310077d53ae4ed9904df42e3f81c634['h01c08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e05] =  I0310077d53ae4ed9904df42e3f81c634['h01c0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e06] =  I0310077d53ae4ed9904df42e3f81c634['h01c0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e07] =  I0310077d53ae4ed9904df42e3f81c634['h01c0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e08] =  I0310077d53ae4ed9904df42e3f81c634['h01c10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e09] =  I0310077d53ae4ed9904df42e3f81c634['h01c12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e0a] =  I0310077d53ae4ed9904df42e3f81c634['h01c14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e0b] =  I0310077d53ae4ed9904df42e3f81c634['h01c16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e0c] =  I0310077d53ae4ed9904df42e3f81c634['h01c18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e0d] =  I0310077d53ae4ed9904df42e3f81c634['h01c1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e0e] =  I0310077d53ae4ed9904df42e3f81c634['h01c1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e0f] =  I0310077d53ae4ed9904df42e3f81c634['h01c1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e10] =  I0310077d53ae4ed9904df42e3f81c634['h01c20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e11] =  I0310077d53ae4ed9904df42e3f81c634['h01c22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e12] =  I0310077d53ae4ed9904df42e3f81c634['h01c24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e13] =  I0310077d53ae4ed9904df42e3f81c634['h01c26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e14] =  I0310077d53ae4ed9904df42e3f81c634['h01c28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e15] =  I0310077d53ae4ed9904df42e3f81c634['h01c2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e16] =  I0310077d53ae4ed9904df42e3f81c634['h01c2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e17] =  I0310077d53ae4ed9904df42e3f81c634['h01c2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e18] =  I0310077d53ae4ed9904df42e3f81c634['h01c30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e19] =  I0310077d53ae4ed9904df42e3f81c634['h01c32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e1a] =  I0310077d53ae4ed9904df42e3f81c634['h01c34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e1b] =  I0310077d53ae4ed9904df42e3f81c634['h01c36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e1c] =  I0310077d53ae4ed9904df42e3f81c634['h01c38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e1d] =  I0310077d53ae4ed9904df42e3f81c634['h01c3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e1e] =  I0310077d53ae4ed9904df42e3f81c634['h01c3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e1f] =  I0310077d53ae4ed9904df42e3f81c634['h01c3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e20] =  I0310077d53ae4ed9904df42e3f81c634['h01c40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e21] =  I0310077d53ae4ed9904df42e3f81c634['h01c42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e22] =  I0310077d53ae4ed9904df42e3f81c634['h01c44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e23] =  I0310077d53ae4ed9904df42e3f81c634['h01c46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e24] =  I0310077d53ae4ed9904df42e3f81c634['h01c48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e25] =  I0310077d53ae4ed9904df42e3f81c634['h01c4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e26] =  I0310077d53ae4ed9904df42e3f81c634['h01c4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e27] =  I0310077d53ae4ed9904df42e3f81c634['h01c4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e28] =  I0310077d53ae4ed9904df42e3f81c634['h01c50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e29] =  I0310077d53ae4ed9904df42e3f81c634['h01c52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e2a] =  I0310077d53ae4ed9904df42e3f81c634['h01c54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e2b] =  I0310077d53ae4ed9904df42e3f81c634['h01c56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e2c] =  I0310077d53ae4ed9904df42e3f81c634['h01c58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e2d] =  I0310077d53ae4ed9904df42e3f81c634['h01c5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e2e] =  I0310077d53ae4ed9904df42e3f81c634['h01c5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e2f] =  I0310077d53ae4ed9904df42e3f81c634['h01c5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e30] =  I0310077d53ae4ed9904df42e3f81c634['h01c60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e31] =  I0310077d53ae4ed9904df42e3f81c634['h01c62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e32] =  I0310077d53ae4ed9904df42e3f81c634['h01c64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e33] =  I0310077d53ae4ed9904df42e3f81c634['h01c66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e34] =  I0310077d53ae4ed9904df42e3f81c634['h01c68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e35] =  I0310077d53ae4ed9904df42e3f81c634['h01c6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e36] =  I0310077d53ae4ed9904df42e3f81c634['h01c6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e37] =  I0310077d53ae4ed9904df42e3f81c634['h01c6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e38] =  I0310077d53ae4ed9904df42e3f81c634['h01c70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e39] =  I0310077d53ae4ed9904df42e3f81c634['h01c72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e3a] =  I0310077d53ae4ed9904df42e3f81c634['h01c74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e3b] =  I0310077d53ae4ed9904df42e3f81c634['h01c76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e3c] =  I0310077d53ae4ed9904df42e3f81c634['h01c78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e3d] =  I0310077d53ae4ed9904df42e3f81c634['h01c7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e3e] =  I0310077d53ae4ed9904df42e3f81c634['h01c7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e3f] =  I0310077d53ae4ed9904df42e3f81c634['h01c7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e40] =  I0310077d53ae4ed9904df42e3f81c634['h01c80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e41] =  I0310077d53ae4ed9904df42e3f81c634['h01c82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e42] =  I0310077d53ae4ed9904df42e3f81c634['h01c84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e43] =  I0310077d53ae4ed9904df42e3f81c634['h01c86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e44] =  I0310077d53ae4ed9904df42e3f81c634['h01c88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e45] =  I0310077d53ae4ed9904df42e3f81c634['h01c8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e46] =  I0310077d53ae4ed9904df42e3f81c634['h01c8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e47] =  I0310077d53ae4ed9904df42e3f81c634['h01c8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e48] =  I0310077d53ae4ed9904df42e3f81c634['h01c90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e49] =  I0310077d53ae4ed9904df42e3f81c634['h01c92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e4a] =  I0310077d53ae4ed9904df42e3f81c634['h01c94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e4b] =  I0310077d53ae4ed9904df42e3f81c634['h01c96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e4c] =  I0310077d53ae4ed9904df42e3f81c634['h01c98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e4d] =  I0310077d53ae4ed9904df42e3f81c634['h01c9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e4e] =  I0310077d53ae4ed9904df42e3f81c634['h01c9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e4f] =  I0310077d53ae4ed9904df42e3f81c634['h01c9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e50] =  I0310077d53ae4ed9904df42e3f81c634['h01ca0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e51] =  I0310077d53ae4ed9904df42e3f81c634['h01ca2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e52] =  I0310077d53ae4ed9904df42e3f81c634['h01ca4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e53] =  I0310077d53ae4ed9904df42e3f81c634['h01ca6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e54] =  I0310077d53ae4ed9904df42e3f81c634['h01ca8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e55] =  I0310077d53ae4ed9904df42e3f81c634['h01caa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e56] =  I0310077d53ae4ed9904df42e3f81c634['h01cac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e57] =  I0310077d53ae4ed9904df42e3f81c634['h01cae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e58] =  I0310077d53ae4ed9904df42e3f81c634['h01cb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e59] =  I0310077d53ae4ed9904df42e3f81c634['h01cb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e5a] =  I0310077d53ae4ed9904df42e3f81c634['h01cb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e5b] =  I0310077d53ae4ed9904df42e3f81c634['h01cb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e5c] =  I0310077d53ae4ed9904df42e3f81c634['h01cb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e5d] =  I0310077d53ae4ed9904df42e3f81c634['h01cba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e5e] =  I0310077d53ae4ed9904df42e3f81c634['h01cbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e5f] =  I0310077d53ae4ed9904df42e3f81c634['h01cbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e60] =  I0310077d53ae4ed9904df42e3f81c634['h01cc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e61] =  I0310077d53ae4ed9904df42e3f81c634['h01cc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e62] =  I0310077d53ae4ed9904df42e3f81c634['h01cc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e63] =  I0310077d53ae4ed9904df42e3f81c634['h01cc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e64] =  I0310077d53ae4ed9904df42e3f81c634['h01cc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e65] =  I0310077d53ae4ed9904df42e3f81c634['h01cca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e66] =  I0310077d53ae4ed9904df42e3f81c634['h01ccc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e67] =  I0310077d53ae4ed9904df42e3f81c634['h01cce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e68] =  I0310077d53ae4ed9904df42e3f81c634['h01cd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e69] =  I0310077d53ae4ed9904df42e3f81c634['h01cd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e6a] =  I0310077d53ae4ed9904df42e3f81c634['h01cd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e6b] =  I0310077d53ae4ed9904df42e3f81c634['h01cd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e6c] =  I0310077d53ae4ed9904df42e3f81c634['h01cd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e6d] =  I0310077d53ae4ed9904df42e3f81c634['h01cda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e6e] =  I0310077d53ae4ed9904df42e3f81c634['h01cdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e6f] =  I0310077d53ae4ed9904df42e3f81c634['h01cde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e70] =  I0310077d53ae4ed9904df42e3f81c634['h01ce0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e71] =  I0310077d53ae4ed9904df42e3f81c634['h01ce2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e72] =  I0310077d53ae4ed9904df42e3f81c634['h01ce4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e73] =  I0310077d53ae4ed9904df42e3f81c634['h01ce6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e74] =  I0310077d53ae4ed9904df42e3f81c634['h01ce8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e75] =  I0310077d53ae4ed9904df42e3f81c634['h01cea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e76] =  I0310077d53ae4ed9904df42e3f81c634['h01cec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e77] =  I0310077d53ae4ed9904df42e3f81c634['h01cee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e78] =  I0310077d53ae4ed9904df42e3f81c634['h01cf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e79] =  I0310077d53ae4ed9904df42e3f81c634['h01cf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e7a] =  I0310077d53ae4ed9904df42e3f81c634['h01cf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e7b] =  I0310077d53ae4ed9904df42e3f81c634['h01cf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e7c] =  I0310077d53ae4ed9904df42e3f81c634['h01cf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e7d] =  I0310077d53ae4ed9904df42e3f81c634['h01cfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e7e] =  I0310077d53ae4ed9904df42e3f81c634['h01cfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e7f] =  I0310077d53ae4ed9904df42e3f81c634['h01cfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e80] =  I0310077d53ae4ed9904df42e3f81c634['h01d00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e81] =  I0310077d53ae4ed9904df42e3f81c634['h01d02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e82] =  I0310077d53ae4ed9904df42e3f81c634['h01d04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e83] =  I0310077d53ae4ed9904df42e3f81c634['h01d06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e84] =  I0310077d53ae4ed9904df42e3f81c634['h01d08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e85] =  I0310077d53ae4ed9904df42e3f81c634['h01d0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e86] =  I0310077d53ae4ed9904df42e3f81c634['h01d0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e87] =  I0310077d53ae4ed9904df42e3f81c634['h01d0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e88] =  I0310077d53ae4ed9904df42e3f81c634['h01d10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e89] =  I0310077d53ae4ed9904df42e3f81c634['h01d12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e8a] =  I0310077d53ae4ed9904df42e3f81c634['h01d14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e8b] =  I0310077d53ae4ed9904df42e3f81c634['h01d16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e8c] =  I0310077d53ae4ed9904df42e3f81c634['h01d18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e8d] =  I0310077d53ae4ed9904df42e3f81c634['h01d1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e8e] =  I0310077d53ae4ed9904df42e3f81c634['h01d1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e8f] =  I0310077d53ae4ed9904df42e3f81c634['h01d1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e90] =  I0310077d53ae4ed9904df42e3f81c634['h01d20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e91] =  I0310077d53ae4ed9904df42e3f81c634['h01d22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e92] =  I0310077d53ae4ed9904df42e3f81c634['h01d24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e93] =  I0310077d53ae4ed9904df42e3f81c634['h01d26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e94] =  I0310077d53ae4ed9904df42e3f81c634['h01d28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e95] =  I0310077d53ae4ed9904df42e3f81c634['h01d2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e96] =  I0310077d53ae4ed9904df42e3f81c634['h01d2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e97] =  I0310077d53ae4ed9904df42e3f81c634['h01d2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e98] =  I0310077d53ae4ed9904df42e3f81c634['h01d30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e99] =  I0310077d53ae4ed9904df42e3f81c634['h01d32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e9a] =  I0310077d53ae4ed9904df42e3f81c634['h01d34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e9b] =  I0310077d53ae4ed9904df42e3f81c634['h01d36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e9c] =  I0310077d53ae4ed9904df42e3f81c634['h01d38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e9d] =  I0310077d53ae4ed9904df42e3f81c634['h01d3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e9e] =  I0310077d53ae4ed9904df42e3f81c634['h01d3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00e9f] =  I0310077d53ae4ed9904df42e3f81c634['h01d3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea0] =  I0310077d53ae4ed9904df42e3f81c634['h01d40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea1] =  I0310077d53ae4ed9904df42e3f81c634['h01d42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea2] =  I0310077d53ae4ed9904df42e3f81c634['h01d44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea3] =  I0310077d53ae4ed9904df42e3f81c634['h01d46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea4] =  I0310077d53ae4ed9904df42e3f81c634['h01d48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea5] =  I0310077d53ae4ed9904df42e3f81c634['h01d4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea6] =  I0310077d53ae4ed9904df42e3f81c634['h01d4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea7] =  I0310077d53ae4ed9904df42e3f81c634['h01d4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea8] =  I0310077d53ae4ed9904df42e3f81c634['h01d50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ea9] =  I0310077d53ae4ed9904df42e3f81c634['h01d52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eaa] =  I0310077d53ae4ed9904df42e3f81c634['h01d54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eab] =  I0310077d53ae4ed9904df42e3f81c634['h01d56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eac] =  I0310077d53ae4ed9904df42e3f81c634['h01d58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ead] =  I0310077d53ae4ed9904df42e3f81c634['h01d5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eae] =  I0310077d53ae4ed9904df42e3f81c634['h01d5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eaf] =  I0310077d53ae4ed9904df42e3f81c634['h01d5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb0] =  I0310077d53ae4ed9904df42e3f81c634['h01d60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb1] =  I0310077d53ae4ed9904df42e3f81c634['h01d62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb2] =  I0310077d53ae4ed9904df42e3f81c634['h01d64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb3] =  I0310077d53ae4ed9904df42e3f81c634['h01d66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb4] =  I0310077d53ae4ed9904df42e3f81c634['h01d68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb5] =  I0310077d53ae4ed9904df42e3f81c634['h01d6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb6] =  I0310077d53ae4ed9904df42e3f81c634['h01d6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb7] =  I0310077d53ae4ed9904df42e3f81c634['h01d6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb8] =  I0310077d53ae4ed9904df42e3f81c634['h01d70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eb9] =  I0310077d53ae4ed9904df42e3f81c634['h01d72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eba] =  I0310077d53ae4ed9904df42e3f81c634['h01d74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ebb] =  I0310077d53ae4ed9904df42e3f81c634['h01d76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ebc] =  I0310077d53ae4ed9904df42e3f81c634['h01d78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ebd] =  I0310077d53ae4ed9904df42e3f81c634['h01d7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ebe] =  I0310077d53ae4ed9904df42e3f81c634['h01d7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ebf] =  I0310077d53ae4ed9904df42e3f81c634['h01d7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec0] =  I0310077d53ae4ed9904df42e3f81c634['h01d80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec1] =  I0310077d53ae4ed9904df42e3f81c634['h01d82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec2] =  I0310077d53ae4ed9904df42e3f81c634['h01d84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec3] =  I0310077d53ae4ed9904df42e3f81c634['h01d86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec4] =  I0310077d53ae4ed9904df42e3f81c634['h01d88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec5] =  I0310077d53ae4ed9904df42e3f81c634['h01d8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec6] =  I0310077d53ae4ed9904df42e3f81c634['h01d8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec7] =  I0310077d53ae4ed9904df42e3f81c634['h01d8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec8] =  I0310077d53ae4ed9904df42e3f81c634['h01d90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ec9] =  I0310077d53ae4ed9904df42e3f81c634['h01d92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eca] =  I0310077d53ae4ed9904df42e3f81c634['h01d94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ecb] =  I0310077d53ae4ed9904df42e3f81c634['h01d96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ecc] =  I0310077d53ae4ed9904df42e3f81c634['h01d98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ecd] =  I0310077d53ae4ed9904df42e3f81c634['h01d9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ece] =  I0310077d53ae4ed9904df42e3f81c634['h01d9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ecf] =  I0310077d53ae4ed9904df42e3f81c634['h01d9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed0] =  I0310077d53ae4ed9904df42e3f81c634['h01da0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed1] =  I0310077d53ae4ed9904df42e3f81c634['h01da2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed2] =  I0310077d53ae4ed9904df42e3f81c634['h01da4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed3] =  I0310077d53ae4ed9904df42e3f81c634['h01da6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed4] =  I0310077d53ae4ed9904df42e3f81c634['h01da8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed5] =  I0310077d53ae4ed9904df42e3f81c634['h01daa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed6] =  I0310077d53ae4ed9904df42e3f81c634['h01dac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed7] =  I0310077d53ae4ed9904df42e3f81c634['h01dae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed8] =  I0310077d53ae4ed9904df42e3f81c634['h01db0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ed9] =  I0310077d53ae4ed9904df42e3f81c634['h01db2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eda] =  I0310077d53ae4ed9904df42e3f81c634['h01db4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00edb] =  I0310077d53ae4ed9904df42e3f81c634['h01db6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00edc] =  I0310077d53ae4ed9904df42e3f81c634['h01db8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00edd] =  I0310077d53ae4ed9904df42e3f81c634['h01dba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ede] =  I0310077d53ae4ed9904df42e3f81c634['h01dbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00edf] =  I0310077d53ae4ed9904df42e3f81c634['h01dbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee0] =  I0310077d53ae4ed9904df42e3f81c634['h01dc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee1] =  I0310077d53ae4ed9904df42e3f81c634['h01dc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee2] =  I0310077d53ae4ed9904df42e3f81c634['h01dc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee3] =  I0310077d53ae4ed9904df42e3f81c634['h01dc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee4] =  I0310077d53ae4ed9904df42e3f81c634['h01dc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee5] =  I0310077d53ae4ed9904df42e3f81c634['h01dca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee6] =  I0310077d53ae4ed9904df42e3f81c634['h01dcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee7] =  I0310077d53ae4ed9904df42e3f81c634['h01dce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee8] =  I0310077d53ae4ed9904df42e3f81c634['h01dd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ee9] =  I0310077d53ae4ed9904df42e3f81c634['h01dd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eea] =  I0310077d53ae4ed9904df42e3f81c634['h01dd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eeb] =  I0310077d53ae4ed9904df42e3f81c634['h01dd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eec] =  I0310077d53ae4ed9904df42e3f81c634['h01dd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eed] =  I0310077d53ae4ed9904df42e3f81c634['h01dda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eee] =  I0310077d53ae4ed9904df42e3f81c634['h01ddc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eef] =  I0310077d53ae4ed9904df42e3f81c634['h01dde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef0] =  I0310077d53ae4ed9904df42e3f81c634['h01de0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef1] =  I0310077d53ae4ed9904df42e3f81c634['h01de2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef2] =  I0310077d53ae4ed9904df42e3f81c634['h01de4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef3] =  I0310077d53ae4ed9904df42e3f81c634['h01de6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef4] =  I0310077d53ae4ed9904df42e3f81c634['h01de8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef5] =  I0310077d53ae4ed9904df42e3f81c634['h01dea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef6] =  I0310077d53ae4ed9904df42e3f81c634['h01dec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef7] =  I0310077d53ae4ed9904df42e3f81c634['h01dee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef8] =  I0310077d53ae4ed9904df42e3f81c634['h01df0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ef9] =  I0310077d53ae4ed9904df42e3f81c634['h01df2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00efa] =  I0310077d53ae4ed9904df42e3f81c634['h01df4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00efb] =  I0310077d53ae4ed9904df42e3f81c634['h01df6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00efc] =  I0310077d53ae4ed9904df42e3f81c634['h01df8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00efd] =  I0310077d53ae4ed9904df42e3f81c634['h01dfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00efe] =  I0310077d53ae4ed9904df42e3f81c634['h01dfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00eff] =  I0310077d53ae4ed9904df42e3f81c634['h01dfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f00] =  I0310077d53ae4ed9904df42e3f81c634['h01e00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f01] =  I0310077d53ae4ed9904df42e3f81c634['h01e02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f02] =  I0310077d53ae4ed9904df42e3f81c634['h01e04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f03] =  I0310077d53ae4ed9904df42e3f81c634['h01e06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f04] =  I0310077d53ae4ed9904df42e3f81c634['h01e08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f05] =  I0310077d53ae4ed9904df42e3f81c634['h01e0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f06] =  I0310077d53ae4ed9904df42e3f81c634['h01e0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f07] =  I0310077d53ae4ed9904df42e3f81c634['h01e0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f08] =  I0310077d53ae4ed9904df42e3f81c634['h01e10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f09] =  I0310077d53ae4ed9904df42e3f81c634['h01e12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f0a] =  I0310077d53ae4ed9904df42e3f81c634['h01e14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f0b] =  I0310077d53ae4ed9904df42e3f81c634['h01e16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f0c] =  I0310077d53ae4ed9904df42e3f81c634['h01e18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f0d] =  I0310077d53ae4ed9904df42e3f81c634['h01e1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f0e] =  I0310077d53ae4ed9904df42e3f81c634['h01e1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f0f] =  I0310077d53ae4ed9904df42e3f81c634['h01e1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f10] =  I0310077d53ae4ed9904df42e3f81c634['h01e20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f11] =  I0310077d53ae4ed9904df42e3f81c634['h01e22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f12] =  I0310077d53ae4ed9904df42e3f81c634['h01e24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f13] =  I0310077d53ae4ed9904df42e3f81c634['h01e26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f14] =  I0310077d53ae4ed9904df42e3f81c634['h01e28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f15] =  I0310077d53ae4ed9904df42e3f81c634['h01e2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f16] =  I0310077d53ae4ed9904df42e3f81c634['h01e2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f17] =  I0310077d53ae4ed9904df42e3f81c634['h01e2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f18] =  I0310077d53ae4ed9904df42e3f81c634['h01e30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f19] =  I0310077d53ae4ed9904df42e3f81c634['h01e32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f1a] =  I0310077d53ae4ed9904df42e3f81c634['h01e34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f1b] =  I0310077d53ae4ed9904df42e3f81c634['h01e36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f1c] =  I0310077d53ae4ed9904df42e3f81c634['h01e38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f1d] =  I0310077d53ae4ed9904df42e3f81c634['h01e3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f1e] =  I0310077d53ae4ed9904df42e3f81c634['h01e3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f1f] =  I0310077d53ae4ed9904df42e3f81c634['h01e3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f20] =  I0310077d53ae4ed9904df42e3f81c634['h01e40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f21] =  I0310077d53ae4ed9904df42e3f81c634['h01e42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f22] =  I0310077d53ae4ed9904df42e3f81c634['h01e44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f23] =  I0310077d53ae4ed9904df42e3f81c634['h01e46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f24] =  I0310077d53ae4ed9904df42e3f81c634['h01e48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f25] =  I0310077d53ae4ed9904df42e3f81c634['h01e4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f26] =  I0310077d53ae4ed9904df42e3f81c634['h01e4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f27] =  I0310077d53ae4ed9904df42e3f81c634['h01e4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f28] =  I0310077d53ae4ed9904df42e3f81c634['h01e50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f29] =  I0310077d53ae4ed9904df42e3f81c634['h01e52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f2a] =  I0310077d53ae4ed9904df42e3f81c634['h01e54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f2b] =  I0310077d53ae4ed9904df42e3f81c634['h01e56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f2c] =  I0310077d53ae4ed9904df42e3f81c634['h01e58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f2d] =  I0310077d53ae4ed9904df42e3f81c634['h01e5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f2e] =  I0310077d53ae4ed9904df42e3f81c634['h01e5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f2f] =  I0310077d53ae4ed9904df42e3f81c634['h01e5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f30] =  I0310077d53ae4ed9904df42e3f81c634['h01e60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f31] =  I0310077d53ae4ed9904df42e3f81c634['h01e62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f32] =  I0310077d53ae4ed9904df42e3f81c634['h01e64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f33] =  I0310077d53ae4ed9904df42e3f81c634['h01e66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f34] =  I0310077d53ae4ed9904df42e3f81c634['h01e68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f35] =  I0310077d53ae4ed9904df42e3f81c634['h01e6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f36] =  I0310077d53ae4ed9904df42e3f81c634['h01e6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f37] =  I0310077d53ae4ed9904df42e3f81c634['h01e6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f38] =  I0310077d53ae4ed9904df42e3f81c634['h01e70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f39] =  I0310077d53ae4ed9904df42e3f81c634['h01e72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f3a] =  I0310077d53ae4ed9904df42e3f81c634['h01e74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f3b] =  I0310077d53ae4ed9904df42e3f81c634['h01e76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f3c] =  I0310077d53ae4ed9904df42e3f81c634['h01e78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f3d] =  I0310077d53ae4ed9904df42e3f81c634['h01e7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f3e] =  I0310077d53ae4ed9904df42e3f81c634['h01e7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f3f] =  I0310077d53ae4ed9904df42e3f81c634['h01e7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f40] =  I0310077d53ae4ed9904df42e3f81c634['h01e80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f41] =  I0310077d53ae4ed9904df42e3f81c634['h01e82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f42] =  I0310077d53ae4ed9904df42e3f81c634['h01e84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f43] =  I0310077d53ae4ed9904df42e3f81c634['h01e86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f44] =  I0310077d53ae4ed9904df42e3f81c634['h01e88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f45] =  I0310077d53ae4ed9904df42e3f81c634['h01e8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f46] =  I0310077d53ae4ed9904df42e3f81c634['h01e8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f47] =  I0310077d53ae4ed9904df42e3f81c634['h01e8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f48] =  I0310077d53ae4ed9904df42e3f81c634['h01e90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f49] =  I0310077d53ae4ed9904df42e3f81c634['h01e92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f4a] =  I0310077d53ae4ed9904df42e3f81c634['h01e94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f4b] =  I0310077d53ae4ed9904df42e3f81c634['h01e96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f4c] =  I0310077d53ae4ed9904df42e3f81c634['h01e98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f4d] =  I0310077d53ae4ed9904df42e3f81c634['h01e9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f4e] =  I0310077d53ae4ed9904df42e3f81c634['h01e9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f4f] =  I0310077d53ae4ed9904df42e3f81c634['h01e9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f50] =  I0310077d53ae4ed9904df42e3f81c634['h01ea0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f51] =  I0310077d53ae4ed9904df42e3f81c634['h01ea2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f52] =  I0310077d53ae4ed9904df42e3f81c634['h01ea4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f53] =  I0310077d53ae4ed9904df42e3f81c634['h01ea6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f54] =  I0310077d53ae4ed9904df42e3f81c634['h01ea8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f55] =  I0310077d53ae4ed9904df42e3f81c634['h01eaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f56] =  I0310077d53ae4ed9904df42e3f81c634['h01eac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f57] =  I0310077d53ae4ed9904df42e3f81c634['h01eae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f58] =  I0310077d53ae4ed9904df42e3f81c634['h01eb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f59] =  I0310077d53ae4ed9904df42e3f81c634['h01eb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f5a] =  I0310077d53ae4ed9904df42e3f81c634['h01eb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f5b] =  I0310077d53ae4ed9904df42e3f81c634['h01eb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f5c] =  I0310077d53ae4ed9904df42e3f81c634['h01eb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f5d] =  I0310077d53ae4ed9904df42e3f81c634['h01eba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f5e] =  I0310077d53ae4ed9904df42e3f81c634['h01ebc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f5f] =  I0310077d53ae4ed9904df42e3f81c634['h01ebe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f60] =  I0310077d53ae4ed9904df42e3f81c634['h01ec0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f61] =  I0310077d53ae4ed9904df42e3f81c634['h01ec2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f62] =  I0310077d53ae4ed9904df42e3f81c634['h01ec4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f63] =  I0310077d53ae4ed9904df42e3f81c634['h01ec6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f64] =  I0310077d53ae4ed9904df42e3f81c634['h01ec8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f65] =  I0310077d53ae4ed9904df42e3f81c634['h01eca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f66] =  I0310077d53ae4ed9904df42e3f81c634['h01ecc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f67] =  I0310077d53ae4ed9904df42e3f81c634['h01ece] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f68] =  I0310077d53ae4ed9904df42e3f81c634['h01ed0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f69] =  I0310077d53ae4ed9904df42e3f81c634['h01ed2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f6a] =  I0310077d53ae4ed9904df42e3f81c634['h01ed4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f6b] =  I0310077d53ae4ed9904df42e3f81c634['h01ed6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f6c] =  I0310077d53ae4ed9904df42e3f81c634['h01ed8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f6d] =  I0310077d53ae4ed9904df42e3f81c634['h01eda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f6e] =  I0310077d53ae4ed9904df42e3f81c634['h01edc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f6f] =  I0310077d53ae4ed9904df42e3f81c634['h01ede] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f70] =  I0310077d53ae4ed9904df42e3f81c634['h01ee0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f71] =  I0310077d53ae4ed9904df42e3f81c634['h01ee2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f72] =  I0310077d53ae4ed9904df42e3f81c634['h01ee4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f73] =  I0310077d53ae4ed9904df42e3f81c634['h01ee6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f74] =  I0310077d53ae4ed9904df42e3f81c634['h01ee8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f75] =  I0310077d53ae4ed9904df42e3f81c634['h01eea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f76] =  I0310077d53ae4ed9904df42e3f81c634['h01eec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f77] =  I0310077d53ae4ed9904df42e3f81c634['h01eee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f78] =  I0310077d53ae4ed9904df42e3f81c634['h01ef0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f79] =  I0310077d53ae4ed9904df42e3f81c634['h01ef2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f7a] =  I0310077d53ae4ed9904df42e3f81c634['h01ef4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f7b] =  I0310077d53ae4ed9904df42e3f81c634['h01ef6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f7c] =  I0310077d53ae4ed9904df42e3f81c634['h01ef8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f7d] =  I0310077d53ae4ed9904df42e3f81c634['h01efa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f7e] =  I0310077d53ae4ed9904df42e3f81c634['h01efc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f7f] =  I0310077d53ae4ed9904df42e3f81c634['h01efe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f80] =  I0310077d53ae4ed9904df42e3f81c634['h01f00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f81] =  I0310077d53ae4ed9904df42e3f81c634['h01f02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f82] =  I0310077d53ae4ed9904df42e3f81c634['h01f04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f83] =  I0310077d53ae4ed9904df42e3f81c634['h01f06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f84] =  I0310077d53ae4ed9904df42e3f81c634['h01f08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f85] =  I0310077d53ae4ed9904df42e3f81c634['h01f0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f86] =  I0310077d53ae4ed9904df42e3f81c634['h01f0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f87] =  I0310077d53ae4ed9904df42e3f81c634['h01f0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f88] =  I0310077d53ae4ed9904df42e3f81c634['h01f10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f89] =  I0310077d53ae4ed9904df42e3f81c634['h01f12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f8a] =  I0310077d53ae4ed9904df42e3f81c634['h01f14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f8b] =  I0310077d53ae4ed9904df42e3f81c634['h01f16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f8c] =  I0310077d53ae4ed9904df42e3f81c634['h01f18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f8d] =  I0310077d53ae4ed9904df42e3f81c634['h01f1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f8e] =  I0310077d53ae4ed9904df42e3f81c634['h01f1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f8f] =  I0310077d53ae4ed9904df42e3f81c634['h01f1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f90] =  I0310077d53ae4ed9904df42e3f81c634['h01f20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f91] =  I0310077d53ae4ed9904df42e3f81c634['h01f22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f92] =  I0310077d53ae4ed9904df42e3f81c634['h01f24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f93] =  I0310077d53ae4ed9904df42e3f81c634['h01f26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f94] =  I0310077d53ae4ed9904df42e3f81c634['h01f28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f95] =  I0310077d53ae4ed9904df42e3f81c634['h01f2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f96] =  I0310077d53ae4ed9904df42e3f81c634['h01f2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f97] =  I0310077d53ae4ed9904df42e3f81c634['h01f2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f98] =  I0310077d53ae4ed9904df42e3f81c634['h01f30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f99] =  I0310077d53ae4ed9904df42e3f81c634['h01f32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f9a] =  I0310077d53ae4ed9904df42e3f81c634['h01f34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f9b] =  I0310077d53ae4ed9904df42e3f81c634['h01f36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f9c] =  I0310077d53ae4ed9904df42e3f81c634['h01f38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f9d] =  I0310077d53ae4ed9904df42e3f81c634['h01f3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f9e] =  I0310077d53ae4ed9904df42e3f81c634['h01f3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00f9f] =  I0310077d53ae4ed9904df42e3f81c634['h01f3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa0] =  I0310077d53ae4ed9904df42e3f81c634['h01f40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa1] =  I0310077d53ae4ed9904df42e3f81c634['h01f42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa2] =  I0310077d53ae4ed9904df42e3f81c634['h01f44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa3] =  I0310077d53ae4ed9904df42e3f81c634['h01f46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa4] =  I0310077d53ae4ed9904df42e3f81c634['h01f48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa5] =  I0310077d53ae4ed9904df42e3f81c634['h01f4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa6] =  I0310077d53ae4ed9904df42e3f81c634['h01f4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa7] =  I0310077d53ae4ed9904df42e3f81c634['h01f4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa8] =  I0310077d53ae4ed9904df42e3f81c634['h01f50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fa9] =  I0310077d53ae4ed9904df42e3f81c634['h01f52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00faa] =  I0310077d53ae4ed9904df42e3f81c634['h01f54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fab] =  I0310077d53ae4ed9904df42e3f81c634['h01f56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fac] =  I0310077d53ae4ed9904df42e3f81c634['h01f58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fad] =  I0310077d53ae4ed9904df42e3f81c634['h01f5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fae] =  I0310077d53ae4ed9904df42e3f81c634['h01f5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00faf] =  I0310077d53ae4ed9904df42e3f81c634['h01f5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb0] =  I0310077d53ae4ed9904df42e3f81c634['h01f60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb1] =  I0310077d53ae4ed9904df42e3f81c634['h01f62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb2] =  I0310077d53ae4ed9904df42e3f81c634['h01f64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb3] =  I0310077d53ae4ed9904df42e3f81c634['h01f66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb4] =  I0310077d53ae4ed9904df42e3f81c634['h01f68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb5] =  I0310077d53ae4ed9904df42e3f81c634['h01f6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb6] =  I0310077d53ae4ed9904df42e3f81c634['h01f6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb7] =  I0310077d53ae4ed9904df42e3f81c634['h01f6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb8] =  I0310077d53ae4ed9904df42e3f81c634['h01f70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fb9] =  I0310077d53ae4ed9904df42e3f81c634['h01f72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fba] =  I0310077d53ae4ed9904df42e3f81c634['h01f74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fbb] =  I0310077d53ae4ed9904df42e3f81c634['h01f76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fbc] =  I0310077d53ae4ed9904df42e3f81c634['h01f78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fbd] =  I0310077d53ae4ed9904df42e3f81c634['h01f7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fbe] =  I0310077d53ae4ed9904df42e3f81c634['h01f7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fbf] =  I0310077d53ae4ed9904df42e3f81c634['h01f7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc0] =  I0310077d53ae4ed9904df42e3f81c634['h01f80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc1] =  I0310077d53ae4ed9904df42e3f81c634['h01f82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc2] =  I0310077d53ae4ed9904df42e3f81c634['h01f84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc3] =  I0310077d53ae4ed9904df42e3f81c634['h01f86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc4] =  I0310077d53ae4ed9904df42e3f81c634['h01f88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc5] =  I0310077d53ae4ed9904df42e3f81c634['h01f8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc6] =  I0310077d53ae4ed9904df42e3f81c634['h01f8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc7] =  I0310077d53ae4ed9904df42e3f81c634['h01f8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc8] =  I0310077d53ae4ed9904df42e3f81c634['h01f90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fc9] =  I0310077d53ae4ed9904df42e3f81c634['h01f92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fca] =  I0310077d53ae4ed9904df42e3f81c634['h01f94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fcb] =  I0310077d53ae4ed9904df42e3f81c634['h01f96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fcc] =  I0310077d53ae4ed9904df42e3f81c634['h01f98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fcd] =  I0310077d53ae4ed9904df42e3f81c634['h01f9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fce] =  I0310077d53ae4ed9904df42e3f81c634['h01f9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fcf] =  I0310077d53ae4ed9904df42e3f81c634['h01f9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd0] =  I0310077d53ae4ed9904df42e3f81c634['h01fa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd1] =  I0310077d53ae4ed9904df42e3f81c634['h01fa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd2] =  I0310077d53ae4ed9904df42e3f81c634['h01fa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd3] =  I0310077d53ae4ed9904df42e3f81c634['h01fa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd4] =  I0310077d53ae4ed9904df42e3f81c634['h01fa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd5] =  I0310077d53ae4ed9904df42e3f81c634['h01faa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd6] =  I0310077d53ae4ed9904df42e3f81c634['h01fac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd7] =  I0310077d53ae4ed9904df42e3f81c634['h01fae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd8] =  I0310077d53ae4ed9904df42e3f81c634['h01fb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fd9] =  I0310077d53ae4ed9904df42e3f81c634['h01fb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fda] =  I0310077d53ae4ed9904df42e3f81c634['h01fb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fdb] =  I0310077d53ae4ed9904df42e3f81c634['h01fb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fdc] =  I0310077d53ae4ed9904df42e3f81c634['h01fb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fdd] =  I0310077d53ae4ed9904df42e3f81c634['h01fba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fde] =  I0310077d53ae4ed9904df42e3f81c634['h01fbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fdf] =  I0310077d53ae4ed9904df42e3f81c634['h01fbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe0] =  I0310077d53ae4ed9904df42e3f81c634['h01fc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe1] =  I0310077d53ae4ed9904df42e3f81c634['h01fc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe2] =  I0310077d53ae4ed9904df42e3f81c634['h01fc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe3] =  I0310077d53ae4ed9904df42e3f81c634['h01fc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe4] =  I0310077d53ae4ed9904df42e3f81c634['h01fc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe5] =  I0310077d53ae4ed9904df42e3f81c634['h01fca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe6] =  I0310077d53ae4ed9904df42e3f81c634['h01fcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe7] =  I0310077d53ae4ed9904df42e3f81c634['h01fce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe8] =  I0310077d53ae4ed9904df42e3f81c634['h01fd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fe9] =  I0310077d53ae4ed9904df42e3f81c634['h01fd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fea] =  I0310077d53ae4ed9904df42e3f81c634['h01fd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00feb] =  I0310077d53ae4ed9904df42e3f81c634['h01fd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fec] =  I0310077d53ae4ed9904df42e3f81c634['h01fd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fed] =  I0310077d53ae4ed9904df42e3f81c634['h01fda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fee] =  I0310077d53ae4ed9904df42e3f81c634['h01fdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fef] =  I0310077d53ae4ed9904df42e3f81c634['h01fde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff0] =  I0310077d53ae4ed9904df42e3f81c634['h01fe0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff1] =  I0310077d53ae4ed9904df42e3f81c634['h01fe2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff2] =  I0310077d53ae4ed9904df42e3f81c634['h01fe4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff3] =  I0310077d53ae4ed9904df42e3f81c634['h01fe6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff4] =  I0310077d53ae4ed9904df42e3f81c634['h01fe8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff5] =  I0310077d53ae4ed9904df42e3f81c634['h01fea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff6] =  I0310077d53ae4ed9904df42e3f81c634['h01fec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff7] =  I0310077d53ae4ed9904df42e3f81c634['h01fee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff8] =  I0310077d53ae4ed9904df42e3f81c634['h01ff0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ff9] =  I0310077d53ae4ed9904df42e3f81c634['h01ff2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ffa] =  I0310077d53ae4ed9904df42e3f81c634['h01ff4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ffb] =  I0310077d53ae4ed9904df42e3f81c634['h01ff6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ffc] =  I0310077d53ae4ed9904df42e3f81c634['h01ff8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ffd] =  I0310077d53ae4ed9904df42e3f81c634['h01ffa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00ffe] =  I0310077d53ae4ed9904df42e3f81c634['h01ffc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h00fff] =  I0310077d53ae4ed9904df42e3f81c634['h01ffe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01000] =  I0310077d53ae4ed9904df42e3f81c634['h02000] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01001] =  I0310077d53ae4ed9904df42e3f81c634['h02002] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01002] =  I0310077d53ae4ed9904df42e3f81c634['h02004] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01003] =  I0310077d53ae4ed9904df42e3f81c634['h02006] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01004] =  I0310077d53ae4ed9904df42e3f81c634['h02008] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01005] =  I0310077d53ae4ed9904df42e3f81c634['h0200a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01006] =  I0310077d53ae4ed9904df42e3f81c634['h0200c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01007] =  I0310077d53ae4ed9904df42e3f81c634['h0200e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01008] =  I0310077d53ae4ed9904df42e3f81c634['h02010] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01009] =  I0310077d53ae4ed9904df42e3f81c634['h02012] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0100a] =  I0310077d53ae4ed9904df42e3f81c634['h02014] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0100b] =  I0310077d53ae4ed9904df42e3f81c634['h02016] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0100c] =  I0310077d53ae4ed9904df42e3f81c634['h02018] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0100d] =  I0310077d53ae4ed9904df42e3f81c634['h0201a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0100e] =  I0310077d53ae4ed9904df42e3f81c634['h0201c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0100f] =  I0310077d53ae4ed9904df42e3f81c634['h0201e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01010] =  I0310077d53ae4ed9904df42e3f81c634['h02020] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01011] =  I0310077d53ae4ed9904df42e3f81c634['h02022] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01012] =  I0310077d53ae4ed9904df42e3f81c634['h02024] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01013] =  I0310077d53ae4ed9904df42e3f81c634['h02026] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01014] =  I0310077d53ae4ed9904df42e3f81c634['h02028] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01015] =  I0310077d53ae4ed9904df42e3f81c634['h0202a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01016] =  I0310077d53ae4ed9904df42e3f81c634['h0202c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01017] =  I0310077d53ae4ed9904df42e3f81c634['h0202e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01018] =  I0310077d53ae4ed9904df42e3f81c634['h02030] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01019] =  I0310077d53ae4ed9904df42e3f81c634['h02032] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0101a] =  I0310077d53ae4ed9904df42e3f81c634['h02034] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0101b] =  I0310077d53ae4ed9904df42e3f81c634['h02036] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0101c] =  I0310077d53ae4ed9904df42e3f81c634['h02038] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0101d] =  I0310077d53ae4ed9904df42e3f81c634['h0203a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0101e] =  I0310077d53ae4ed9904df42e3f81c634['h0203c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0101f] =  I0310077d53ae4ed9904df42e3f81c634['h0203e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01020] =  I0310077d53ae4ed9904df42e3f81c634['h02040] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01021] =  I0310077d53ae4ed9904df42e3f81c634['h02042] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01022] =  I0310077d53ae4ed9904df42e3f81c634['h02044] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01023] =  I0310077d53ae4ed9904df42e3f81c634['h02046] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01024] =  I0310077d53ae4ed9904df42e3f81c634['h02048] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01025] =  I0310077d53ae4ed9904df42e3f81c634['h0204a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01026] =  I0310077d53ae4ed9904df42e3f81c634['h0204c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01027] =  I0310077d53ae4ed9904df42e3f81c634['h0204e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01028] =  I0310077d53ae4ed9904df42e3f81c634['h02050] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01029] =  I0310077d53ae4ed9904df42e3f81c634['h02052] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0102a] =  I0310077d53ae4ed9904df42e3f81c634['h02054] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0102b] =  I0310077d53ae4ed9904df42e3f81c634['h02056] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0102c] =  I0310077d53ae4ed9904df42e3f81c634['h02058] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0102d] =  I0310077d53ae4ed9904df42e3f81c634['h0205a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0102e] =  I0310077d53ae4ed9904df42e3f81c634['h0205c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0102f] =  I0310077d53ae4ed9904df42e3f81c634['h0205e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01030] =  I0310077d53ae4ed9904df42e3f81c634['h02060] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01031] =  I0310077d53ae4ed9904df42e3f81c634['h02062] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01032] =  I0310077d53ae4ed9904df42e3f81c634['h02064] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01033] =  I0310077d53ae4ed9904df42e3f81c634['h02066] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01034] =  I0310077d53ae4ed9904df42e3f81c634['h02068] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01035] =  I0310077d53ae4ed9904df42e3f81c634['h0206a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01036] =  I0310077d53ae4ed9904df42e3f81c634['h0206c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01037] =  I0310077d53ae4ed9904df42e3f81c634['h0206e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01038] =  I0310077d53ae4ed9904df42e3f81c634['h02070] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01039] =  I0310077d53ae4ed9904df42e3f81c634['h02072] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0103a] =  I0310077d53ae4ed9904df42e3f81c634['h02074] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0103b] =  I0310077d53ae4ed9904df42e3f81c634['h02076] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0103c] =  I0310077d53ae4ed9904df42e3f81c634['h02078] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0103d] =  I0310077d53ae4ed9904df42e3f81c634['h0207a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0103e] =  I0310077d53ae4ed9904df42e3f81c634['h0207c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0103f] =  I0310077d53ae4ed9904df42e3f81c634['h0207e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01040] =  I0310077d53ae4ed9904df42e3f81c634['h02080] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01041] =  I0310077d53ae4ed9904df42e3f81c634['h02082] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01042] =  I0310077d53ae4ed9904df42e3f81c634['h02084] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01043] =  I0310077d53ae4ed9904df42e3f81c634['h02086] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01044] =  I0310077d53ae4ed9904df42e3f81c634['h02088] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01045] =  I0310077d53ae4ed9904df42e3f81c634['h0208a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01046] =  I0310077d53ae4ed9904df42e3f81c634['h0208c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01047] =  I0310077d53ae4ed9904df42e3f81c634['h0208e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01048] =  I0310077d53ae4ed9904df42e3f81c634['h02090] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01049] =  I0310077d53ae4ed9904df42e3f81c634['h02092] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0104a] =  I0310077d53ae4ed9904df42e3f81c634['h02094] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0104b] =  I0310077d53ae4ed9904df42e3f81c634['h02096] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0104c] =  I0310077d53ae4ed9904df42e3f81c634['h02098] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0104d] =  I0310077d53ae4ed9904df42e3f81c634['h0209a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0104e] =  I0310077d53ae4ed9904df42e3f81c634['h0209c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0104f] =  I0310077d53ae4ed9904df42e3f81c634['h0209e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01050] =  I0310077d53ae4ed9904df42e3f81c634['h020a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01051] =  I0310077d53ae4ed9904df42e3f81c634['h020a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01052] =  I0310077d53ae4ed9904df42e3f81c634['h020a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01053] =  I0310077d53ae4ed9904df42e3f81c634['h020a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01054] =  I0310077d53ae4ed9904df42e3f81c634['h020a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01055] =  I0310077d53ae4ed9904df42e3f81c634['h020aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01056] =  I0310077d53ae4ed9904df42e3f81c634['h020ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01057] =  I0310077d53ae4ed9904df42e3f81c634['h020ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01058] =  I0310077d53ae4ed9904df42e3f81c634['h020b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01059] =  I0310077d53ae4ed9904df42e3f81c634['h020b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0105a] =  I0310077d53ae4ed9904df42e3f81c634['h020b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0105b] =  I0310077d53ae4ed9904df42e3f81c634['h020b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0105c] =  I0310077d53ae4ed9904df42e3f81c634['h020b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0105d] =  I0310077d53ae4ed9904df42e3f81c634['h020ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0105e] =  I0310077d53ae4ed9904df42e3f81c634['h020bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0105f] =  I0310077d53ae4ed9904df42e3f81c634['h020be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01060] =  I0310077d53ae4ed9904df42e3f81c634['h020c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01061] =  I0310077d53ae4ed9904df42e3f81c634['h020c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01062] =  I0310077d53ae4ed9904df42e3f81c634['h020c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01063] =  I0310077d53ae4ed9904df42e3f81c634['h020c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01064] =  I0310077d53ae4ed9904df42e3f81c634['h020c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01065] =  I0310077d53ae4ed9904df42e3f81c634['h020ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01066] =  I0310077d53ae4ed9904df42e3f81c634['h020cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01067] =  I0310077d53ae4ed9904df42e3f81c634['h020ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01068] =  I0310077d53ae4ed9904df42e3f81c634['h020d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01069] =  I0310077d53ae4ed9904df42e3f81c634['h020d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0106a] =  I0310077d53ae4ed9904df42e3f81c634['h020d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0106b] =  I0310077d53ae4ed9904df42e3f81c634['h020d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0106c] =  I0310077d53ae4ed9904df42e3f81c634['h020d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0106d] =  I0310077d53ae4ed9904df42e3f81c634['h020da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0106e] =  I0310077d53ae4ed9904df42e3f81c634['h020dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0106f] =  I0310077d53ae4ed9904df42e3f81c634['h020de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01070] =  I0310077d53ae4ed9904df42e3f81c634['h020e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01071] =  I0310077d53ae4ed9904df42e3f81c634['h020e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01072] =  I0310077d53ae4ed9904df42e3f81c634['h020e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01073] =  I0310077d53ae4ed9904df42e3f81c634['h020e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01074] =  I0310077d53ae4ed9904df42e3f81c634['h020e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01075] =  I0310077d53ae4ed9904df42e3f81c634['h020ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01076] =  I0310077d53ae4ed9904df42e3f81c634['h020ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01077] =  I0310077d53ae4ed9904df42e3f81c634['h020ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01078] =  I0310077d53ae4ed9904df42e3f81c634['h020f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01079] =  I0310077d53ae4ed9904df42e3f81c634['h020f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0107a] =  I0310077d53ae4ed9904df42e3f81c634['h020f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0107b] =  I0310077d53ae4ed9904df42e3f81c634['h020f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0107c] =  I0310077d53ae4ed9904df42e3f81c634['h020f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0107d] =  I0310077d53ae4ed9904df42e3f81c634['h020fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0107e] =  I0310077d53ae4ed9904df42e3f81c634['h020fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0107f] =  I0310077d53ae4ed9904df42e3f81c634['h020fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01080] =  I0310077d53ae4ed9904df42e3f81c634['h02100] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01081] =  I0310077d53ae4ed9904df42e3f81c634['h02102] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01082] =  I0310077d53ae4ed9904df42e3f81c634['h02104] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01083] =  I0310077d53ae4ed9904df42e3f81c634['h02106] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01084] =  I0310077d53ae4ed9904df42e3f81c634['h02108] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01085] =  I0310077d53ae4ed9904df42e3f81c634['h0210a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01086] =  I0310077d53ae4ed9904df42e3f81c634['h0210c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01087] =  I0310077d53ae4ed9904df42e3f81c634['h0210e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01088] =  I0310077d53ae4ed9904df42e3f81c634['h02110] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01089] =  I0310077d53ae4ed9904df42e3f81c634['h02112] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0108a] =  I0310077d53ae4ed9904df42e3f81c634['h02114] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0108b] =  I0310077d53ae4ed9904df42e3f81c634['h02116] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0108c] =  I0310077d53ae4ed9904df42e3f81c634['h02118] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0108d] =  I0310077d53ae4ed9904df42e3f81c634['h0211a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0108e] =  I0310077d53ae4ed9904df42e3f81c634['h0211c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0108f] =  I0310077d53ae4ed9904df42e3f81c634['h0211e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01090] =  I0310077d53ae4ed9904df42e3f81c634['h02120] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01091] =  I0310077d53ae4ed9904df42e3f81c634['h02122] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01092] =  I0310077d53ae4ed9904df42e3f81c634['h02124] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01093] =  I0310077d53ae4ed9904df42e3f81c634['h02126] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01094] =  I0310077d53ae4ed9904df42e3f81c634['h02128] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01095] =  I0310077d53ae4ed9904df42e3f81c634['h0212a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01096] =  I0310077d53ae4ed9904df42e3f81c634['h0212c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01097] =  I0310077d53ae4ed9904df42e3f81c634['h0212e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01098] =  I0310077d53ae4ed9904df42e3f81c634['h02130] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01099] =  I0310077d53ae4ed9904df42e3f81c634['h02132] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0109a] =  I0310077d53ae4ed9904df42e3f81c634['h02134] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0109b] =  I0310077d53ae4ed9904df42e3f81c634['h02136] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0109c] =  I0310077d53ae4ed9904df42e3f81c634['h02138] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0109d] =  I0310077d53ae4ed9904df42e3f81c634['h0213a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0109e] =  I0310077d53ae4ed9904df42e3f81c634['h0213c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0109f] =  I0310077d53ae4ed9904df42e3f81c634['h0213e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a0] =  I0310077d53ae4ed9904df42e3f81c634['h02140] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a1] =  I0310077d53ae4ed9904df42e3f81c634['h02142] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a2] =  I0310077d53ae4ed9904df42e3f81c634['h02144] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a3] =  I0310077d53ae4ed9904df42e3f81c634['h02146] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a4] =  I0310077d53ae4ed9904df42e3f81c634['h02148] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a5] =  I0310077d53ae4ed9904df42e3f81c634['h0214a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a6] =  I0310077d53ae4ed9904df42e3f81c634['h0214c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a7] =  I0310077d53ae4ed9904df42e3f81c634['h0214e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a8] =  I0310077d53ae4ed9904df42e3f81c634['h02150] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010a9] =  I0310077d53ae4ed9904df42e3f81c634['h02152] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010aa] =  I0310077d53ae4ed9904df42e3f81c634['h02154] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ab] =  I0310077d53ae4ed9904df42e3f81c634['h02156] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ac] =  I0310077d53ae4ed9904df42e3f81c634['h02158] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ad] =  I0310077d53ae4ed9904df42e3f81c634['h0215a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ae] =  I0310077d53ae4ed9904df42e3f81c634['h0215c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010af] =  I0310077d53ae4ed9904df42e3f81c634['h0215e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b0] =  I0310077d53ae4ed9904df42e3f81c634['h02160] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b1] =  I0310077d53ae4ed9904df42e3f81c634['h02162] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b2] =  I0310077d53ae4ed9904df42e3f81c634['h02164] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b3] =  I0310077d53ae4ed9904df42e3f81c634['h02166] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b4] =  I0310077d53ae4ed9904df42e3f81c634['h02168] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b5] =  I0310077d53ae4ed9904df42e3f81c634['h0216a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b6] =  I0310077d53ae4ed9904df42e3f81c634['h0216c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b7] =  I0310077d53ae4ed9904df42e3f81c634['h0216e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b8] =  I0310077d53ae4ed9904df42e3f81c634['h02170] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010b9] =  I0310077d53ae4ed9904df42e3f81c634['h02172] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ba] =  I0310077d53ae4ed9904df42e3f81c634['h02174] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010bb] =  I0310077d53ae4ed9904df42e3f81c634['h02176] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010bc] =  I0310077d53ae4ed9904df42e3f81c634['h02178] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010bd] =  I0310077d53ae4ed9904df42e3f81c634['h0217a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010be] =  I0310077d53ae4ed9904df42e3f81c634['h0217c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010bf] =  I0310077d53ae4ed9904df42e3f81c634['h0217e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c0] =  I0310077d53ae4ed9904df42e3f81c634['h02180] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c1] =  I0310077d53ae4ed9904df42e3f81c634['h02182] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c2] =  I0310077d53ae4ed9904df42e3f81c634['h02184] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c3] =  I0310077d53ae4ed9904df42e3f81c634['h02186] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c4] =  I0310077d53ae4ed9904df42e3f81c634['h02188] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c5] =  I0310077d53ae4ed9904df42e3f81c634['h0218a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c6] =  I0310077d53ae4ed9904df42e3f81c634['h0218c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c7] =  I0310077d53ae4ed9904df42e3f81c634['h0218e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c8] =  I0310077d53ae4ed9904df42e3f81c634['h02190] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010c9] =  I0310077d53ae4ed9904df42e3f81c634['h02192] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ca] =  I0310077d53ae4ed9904df42e3f81c634['h02194] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010cb] =  I0310077d53ae4ed9904df42e3f81c634['h02196] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010cc] =  I0310077d53ae4ed9904df42e3f81c634['h02198] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010cd] =  I0310077d53ae4ed9904df42e3f81c634['h0219a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ce] =  I0310077d53ae4ed9904df42e3f81c634['h0219c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010cf] =  I0310077d53ae4ed9904df42e3f81c634['h0219e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d0] =  I0310077d53ae4ed9904df42e3f81c634['h021a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d1] =  I0310077d53ae4ed9904df42e3f81c634['h021a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d2] =  I0310077d53ae4ed9904df42e3f81c634['h021a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d3] =  I0310077d53ae4ed9904df42e3f81c634['h021a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d4] =  I0310077d53ae4ed9904df42e3f81c634['h021a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d5] =  I0310077d53ae4ed9904df42e3f81c634['h021aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d6] =  I0310077d53ae4ed9904df42e3f81c634['h021ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d7] =  I0310077d53ae4ed9904df42e3f81c634['h021ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d8] =  I0310077d53ae4ed9904df42e3f81c634['h021b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010d9] =  I0310077d53ae4ed9904df42e3f81c634['h021b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010da] =  I0310077d53ae4ed9904df42e3f81c634['h021b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010db] =  I0310077d53ae4ed9904df42e3f81c634['h021b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010dc] =  I0310077d53ae4ed9904df42e3f81c634['h021b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010dd] =  I0310077d53ae4ed9904df42e3f81c634['h021ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010de] =  I0310077d53ae4ed9904df42e3f81c634['h021bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010df] =  I0310077d53ae4ed9904df42e3f81c634['h021be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e0] =  I0310077d53ae4ed9904df42e3f81c634['h021c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e1] =  I0310077d53ae4ed9904df42e3f81c634['h021c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e2] =  I0310077d53ae4ed9904df42e3f81c634['h021c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e3] =  I0310077d53ae4ed9904df42e3f81c634['h021c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e4] =  I0310077d53ae4ed9904df42e3f81c634['h021c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e5] =  I0310077d53ae4ed9904df42e3f81c634['h021ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e6] =  I0310077d53ae4ed9904df42e3f81c634['h021cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e7] =  I0310077d53ae4ed9904df42e3f81c634['h021ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e8] =  I0310077d53ae4ed9904df42e3f81c634['h021d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010e9] =  I0310077d53ae4ed9904df42e3f81c634['h021d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ea] =  I0310077d53ae4ed9904df42e3f81c634['h021d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010eb] =  I0310077d53ae4ed9904df42e3f81c634['h021d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ec] =  I0310077d53ae4ed9904df42e3f81c634['h021d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ed] =  I0310077d53ae4ed9904df42e3f81c634['h021da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ee] =  I0310077d53ae4ed9904df42e3f81c634['h021dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ef] =  I0310077d53ae4ed9904df42e3f81c634['h021de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f0] =  I0310077d53ae4ed9904df42e3f81c634['h021e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f1] =  I0310077d53ae4ed9904df42e3f81c634['h021e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f2] =  I0310077d53ae4ed9904df42e3f81c634['h021e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f3] =  I0310077d53ae4ed9904df42e3f81c634['h021e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f4] =  I0310077d53ae4ed9904df42e3f81c634['h021e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f5] =  I0310077d53ae4ed9904df42e3f81c634['h021ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f6] =  I0310077d53ae4ed9904df42e3f81c634['h021ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f7] =  I0310077d53ae4ed9904df42e3f81c634['h021ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f8] =  I0310077d53ae4ed9904df42e3f81c634['h021f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010f9] =  I0310077d53ae4ed9904df42e3f81c634['h021f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010fa] =  I0310077d53ae4ed9904df42e3f81c634['h021f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010fb] =  I0310077d53ae4ed9904df42e3f81c634['h021f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010fc] =  I0310077d53ae4ed9904df42e3f81c634['h021f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010fd] =  I0310077d53ae4ed9904df42e3f81c634['h021fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010fe] =  I0310077d53ae4ed9904df42e3f81c634['h021fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h010ff] =  I0310077d53ae4ed9904df42e3f81c634['h021fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01100] =  I0310077d53ae4ed9904df42e3f81c634['h02200] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01101] =  I0310077d53ae4ed9904df42e3f81c634['h02202] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01102] =  I0310077d53ae4ed9904df42e3f81c634['h02204] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01103] =  I0310077d53ae4ed9904df42e3f81c634['h02206] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01104] =  I0310077d53ae4ed9904df42e3f81c634['h02208] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01105] =  I0310077d53ae4ed9904df42e3f81c634['h0220a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01106] =  I0310077d53ae4ed9904df42e3f81c634['h0220c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01107] =  I0310077d53ae4ed9904df42e3f81c634['h0220e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01108] =  I0310077d53ae4ed9904df42e3f81c634['h02210] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01109] =  I0310077d53ae4ed9904df42e3f81c634['h02212] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0110a] =  I0310077d53ae4ed9904df42e3f81c634['h02214] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0110b] =  I0310077d53ae4ed9904df42e3f81c634['h02216] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0110c] =  I0310077d53ae4ed9904df42e3f81c634['h02218] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0110d] =  I0310077d53ae4ed9904df42e3f81c634['h0221a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0110e] =  I0310077d53ae4ed9904df42e3f81c634['h0221c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0110f] =  I0310077d53ae4ed9904df42e3f81c634['h0221e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01110] =  I0310077d53ae4ed9904df42e3f81c634['h02220] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01111] =  I0310077d53ae4ed9904df42e3f81c634['h02222] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01112] =  I0310077d53ae4ed9904df42e3f81c634['h02224] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01113] =  I0310077d53ae4ed9904df42e3f81c634['h02226] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01114] =  I0310077d53ae4ed9904df42e3f81c634['h02228] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01115] =  I0310077d53ae4ed9904df42e3f81c634['h0222a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01116] =  I0310077d53ae4ed9904df42e3f81c634['h0222c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01117] =  I0310077d53ae4ed9904df42e3f81c634['h0222e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01118] =  I0310077d53ae4ed9904df42e3f81c634['h02230] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01119] =  I0310077d53ae4ed9904df42e3f81c634['h02232] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0111a] =  I0310077d53ae4ed9904df42e3f81c634['h02234] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0111b] =  I0310077d53ae4ed9904df42e3f81c634['h02236] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0111c] =  I0310077d53ae4ed9904df42e3f81c634['h02238] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0111d] =  I0310077d53ae4ed9904df42e3f81c634['h0223a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0111e] =  I0310077d53ae4ed9904df42e3f81c634['h0223c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0111f] =  I0310077d53ae4ed9904df42e3f81c634['h0223e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01120] =  I0310077d53ae4ed9904df42e3f81c634['h02240] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01121] =  I0310077d53ae4ed9904df42e3f81c634['h02242] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01122] =  I0310077d53ae4ed9904df42e3f81c634['h02244] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01123] =  I0310077d53ae4ed9904df42e3f81c634['h02246] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01124] =  I0310077d53ae4ed9904df42e3f81c634['h02248] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01125] =  I0310077d53ae4ed9904df42e3f81c634['h0224a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01126] =  I0310077d53ae4ed9904df42e3f81c634['h0224c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01127] =  I0310077d53ae4ed9904df42e3f81c634['h0224e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01128] =  I0310077d53ae4ed9904df42e3f81c634['h02250] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01129] =  I0310077d53ae4ed9904df42e3f81c634['h02252] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0112a] =  I0310077d53ae4ed9904df42e3f81c634['h02254] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0112b] =  I0310077d53ae4ed9904df42e3f81c634['h02256] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0112c] =  I0310077d53ae4ed9904df42e3f81c634['h02258] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0112d] =  I0310077d53ae4ed9904df42e3f81c634['h0225a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0112e] =  I0310077d53ae4ed9904df42e3f81c634['h0225c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0112f] =  I0310077d53ae4ed9904df42e3f81c634['h0225e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01130] =  I0310077d53ae4ed9904df42e3f81c634['h02260] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01131] =  I0310077d53ae4ed9904df42e3f81c634['h02262] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01132] =  I0310077d53ae4ed9904df42e3f81c634['h02264] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01133] =  I0310077d53ae4ed9904df42e3f81c634['h02266] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01134] =  I0310077d53ae4ed9904df42e3f81c634['h02268] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01135] =  I0310077d53ae4ed9904df42e3f81c634['h0226a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01136] =  I0310077d53ae4ed9904df42e3f81c634['h0226c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01137] =  I0310077d53ae4ed9904df42e3f81c634['h0226e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01138] =  I0310077d53ae4ed9904df42e3f81c634['h02270] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01139] =  I0310077d53ae4ed9904df42e3f81c634['h02272] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0113a] =  I0310077d53ae4ed9904df42e3f81c634['h02274] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0113b] =  I0310077d53ae4ed9904df42e3f81c634['h02276] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0113c] =  I0310077d53ae4ed9904df42e3f81c634['h02278] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0113d] =  I0310077d53ae4ed9904df42e3f81c634['h0227a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0113e] =  I0310077d53ae4ed9904df42e3f81c634['h0227c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0113f] =  I0310077d53ae4ed9904df42e3f81c634['h0227e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01140] =  I0310077d53ae4ed9904df42e3f81c634['h02280] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01141] =  I0310077d53ae4ed9904df42e3f81c634['h02282] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01142] =  I0310077d53ae4ed9904df42e3f81c634['h02284] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01143] =  I0310077d53ae4ed9904df42e3f81c634['h02286] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01144] =  I0310077d53ae4ed9904df42e3f81c634['h02288] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01145] =  I0310077d53ae4ed9904df42e3f81c634['h0228a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01146] =  I0310077d53ae4ed9904df42e3f81c634['h0228c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01147] =  I0310077d53ae4ed9904df42e3f81c634['h0228e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01148] =  I0310077d53ae4ed9904df42e3f81c634['h02290] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01149] =  I0310077d53ae4ed9904df42e3f81c634['h02292] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0114a] =  I0310077d53ae4ed9904df42e3f81c634['h02294] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0114b] =  I0310077d53ae4ed9904df42e3f81c634['h02296] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0114c] =  I0310077d53ae4ed9904df42e3f81c634['h02298] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0114d] =  I0310077d53ae4ed9904df42e3f81c634['h0229a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0114e] =  I0310077d53ae4ed9904df42e3f81c634['h0229c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0114f] =  I0310077d53ae4ed9904df42e3f81c634['h0229e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01150] =  I0310077d53ae4ed9904df42e3f81c634['h022a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01151] =  I0310077d53ae4ed9904df42e3f81c634['h022a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01152] =  I0310077d53ae4ed9904df42e3f81c634['h022a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01153] =  I0310077d53ae4ed9904df42e3f81c634['h022a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01154] =  I0310077d53ae4ed9904df42e3f81c634['h022a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01155] =  I0310077d53ae4ed9904df42e3f81c634['h022aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01156] =  I0310077d53ae4ed9904df42e3f81c634['h022ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01157] =  I0310077d53ae4ed9904df42e3f81c634['h022ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01158] =  I0310077d53ae4ed9904df42e3f81c634['h022b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01159] =  I0310077d53ae4ed9904df42e3f81c634['h022b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0115a] =  I0310077d53ae4ed9904df42e3f81c634['h022b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0115b] =  I0310077d53ae4ed9904df42e3f81c634['h022b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0115c] =  I0310077d53ae4ed9904df42e3f81c634['h022b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0115d] =  I0310077d53ae4ed9904df42e3f81c634['h022ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0115e] =  I0310077d53ae4ed9904df42e3f81c634['h022bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0115f] =  I0310077d53ae4ed9904df42e3f81c634['h022be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01160] =  I0310077d53ae4ed9904df42e3f81c634['h022c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01161] =  I0310077d53ae4ed9904df42e3f81c634['h022c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01162] =  I0310077d53ae4ed9904df42e3f81c634['h022c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01163] =  I0310077d53ae4ed9904df42e3f81c634['h022c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01164] =  I0310077d53ae4ed9904df42e3f81c634['h022c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01165] =  I0310077d53ae4ed9904df42e3f81c634['h022ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01166] =  I0310077d53ae4ed9904df42e3f81c634['h022cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01167] =  I0310077d53ae4ed9904df42e3f81c634['h022ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01168] =  I0310077d53ae4ed9904df42e3f81c634['h022d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01169] =  I0310077d53ae4ed9904df42e3f81c634['h022d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0116a] =  I0310077d53ae4ed9904df42e3f81c634['h022d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0116b] =  I0310077d53ae4ed9904df42e3f81c634['h022d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0116c] =  I0310077d53ae4ed9904df42e3f81c634['h022d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0116d] =  I0310077d53ae4ed9904df42e3f81c634['h022da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0116e] =  I0310077d53ae4ed9904df42e3f81c634['h022dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0116f] =  I0310077d53ae4ed9904df42e3f81c634['h022de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01170] =  I0310077d53ae4ed9904df42e3f81c634['h022e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01171] =  I0310077d53ae4ed9904df42e3f81c634['h022e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01172] =  I0310077d53ae4ed9904df42e3f81c634['h022e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01173] =  I0310077d53ae4ed9904df42e3f81c634['h022e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01174] =  I0310077d53ae4ed9904df42e3f81c634['h022e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01175] =  I0310077d53ae4ed9904df42e3f81c634['h022ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01176] =  I0310077d53ae4ed9904df42e3f81c634['h022ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01177] =  I0310077d53ae4ed9904df42e3f81c634['h022ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01178] =  I0310077d53ae4ed9904df42e3f81c634['h022f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01179] =  I0310077d53ae4ed9904df42e3f81c634['h022f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0117a] =  I0310077d53ae4ed9904df42e3f81c634['h022f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0117b] =  I0310077d53ae4ed9904df42e3f81c634['h022f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0117c] =  I0310077d53ae4ed9904df42e3f81c634['h022f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0117d] =  I0310077d53ae4ed9904df42e3f81c634['h022fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0117e] =  I0310077d53ae4ed9904df42e3f81c634['h022fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0117f] =  I0310077d53ae4ed9904df42e3f81c634['h022fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01180] =  I0310077d53ae4ed9904df42e3f81c634['h02300] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01181] =  I0310077d53ae4ed9904df42e3f81c634['h02302] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01182] =  I0310077d53ae4ed9904df42e3f81c634['h02304] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01183] =  I0310077d53ae4ed9904df42e3f81c634['h02306] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01184] =  I0310077d53ae4ed9904df42e3f81c634['h02308] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01185] =  I0310077d53ae4ed9904df42e3f81c634['h0230a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01186] =  I0310077d53ae4ed9904df42e3f81c634['h0230c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01187] =  I0310077d53ae4ed9904df42e3f81c634['h0230e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01188] =  I0310077d53ae4ed9904df42e3f81c634['h02310] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01189] =  I0310077d53ae4ed9904df42e3f81c634['h02312] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0118a] =  I0310077d53ae4ed9904df42e3f81c634['h02314] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0118b] =  I0310077d53ae4ed9904df42e3f81c634['h02316] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0118c] =  I0310077d53ae4ed9904df42e3f81c634['h02318] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0118d] =  I0310077d53ae4ed9904df42e3f81c634['h0231a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0118e] =  I0310077d53ae4ed9904df42e3f81c634['h0231c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0118f] =  I0310077d53ae4ed9904df42e3f81c634['h0231e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01190] =  I0310077d53ae4ed9904df42e3f81c634['h02320] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01191] =  I0310077d53ae4ed9904df42e3f81c634['h02322] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01192] =  I0310077d53ae4ed9904df42e3f81c634['h02324] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01193] =  I0310077d53ae4ed9904df42e3f81c634['h02326] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01194] =  I0310077d53ae4ed9904df42e3f81c634['h02328] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01195] =  I0310077d53ae4ed9904df42e3f81c634['h0232a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01196] =  I0310077d53ae4ed9904df42e3f81c634['h0232c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01197] =  I0310077d53ae4ed9904df42e3f81c634['h0232e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01198] =  I0310077d53ae4ed9904df42e3f81c634['h02330] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01199] =  I0310077d53ae4ed9904df42e3f81c634['h02332] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0119a] =  I0310077d53ae4ed9904df42e3f81c634['h02334] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0119b] =  I0310077d53ae4ed9904df42e3f81c634['h02336] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0119c] =  I0310077d53ae4ed9904df42e3f81c634['h02338] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0119d] =  I0310077d53ae4ed9904df42e3f81c634['h0233a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0119e] =  I0310077d53ae4ed9904df42e3f81c634['h0233c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0119f] =  I0310077d53ae4ed9904df42e3f81c634['h0233e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a0] =  I0310077d53ae4ed9904df42e3f81c634['h02340] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a1] =  I0310077d53ae4ed9904df42e3f81c634['h02342] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a2] =  I0310077d53ae4ed9904df42e3f81c634['h02344] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a3] =  I0310077d53ae4ed9904df42e3f81c634['h02346] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a4] =  I0310077d53ae4ed9904df42e3f81c634['h02348] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a5] =  I0310077d53ae4ed9904df42e3f81c634['h0234a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a6] =  I0310077d53ae4ed9904df42e3f81c634['h0234c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a7] =  I0310077d53ae4ed9904df42e3f81c634['h0234e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a8] =  I0310077d53ae4ed9904df42e3f81c634['h02350] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011a9] =  I0310077d53ae4ed9904df42e3f81c634['h02352] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011aa] =  I0310077d53ae4ed9904df42e3f81c634['h02354] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ab] =  I0310077d53ae4ed9904df42e3f81c634['h02356] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ac] =  I0310077d53ae4ed9904df42e3f81c634['h02358] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ad] =  I0310077d53ae4ed9904df42e3f81c634['h0235a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ae] =  I0310077d53ae4ed9904df42e3f81c634['h0235c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011af] =  I0310077d53ae4ed9904df42e3f81c634['h0235e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b0] =  I0310077d53ae4ed9904df42e3f81c634['h02360] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b1] =  I0310077d53ae4ed9904df42e3f81c634['h02362] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b2] =  I0310077d53ae4ed9904df42e3f81c634['h02364] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b3] =  I0310077d53ae4ed9904df42e3f81c634['h02366] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b4] =  I0310077d53ae4ed9904df42e3f81c634['h02368] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b5] =  I0310077d53ae4ed9904df42e3f81c634['h0236a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b6] =  I0310077d53ae4ed9904df42e3f81c634['h0236c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b7] =  I0310077d53ae4ed9904df42e3f81c634['h0236e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b8] =  I0310077d53ae4ed9904df42e3f81c634['h02370] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011b9] =  I0310077d53ae4ed9904df42e3f81c634['h02372] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ba] =  I0310077d53ae4ed9904df42e3f81c634['h02374] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011bb] =  I0310077d53ae4ed9904df42e3f81c634['h02376] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011bc] =  I0310077d53ae4ed9904df42e3f81c634['h02378] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011bd] =  I0310077d53ae4ed9904df42e3f81c634['h0237a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011be] =  I0310077d53ae4ed9904df42e3f81c634['h0237c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011bf] =  I0310077d53ae4ed9904df42e3f81c634['h0237e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c0] =  I0310077d53ae4ed9904df42e3f81c634['h02380] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c1] =  I0310077d53ae4ed9904df42e3f81c634['h02382] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c2] =  I0310077d53ae4ed9904df42e3f81c634['h02384] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c3] =  I0310077d53ae4ed9904df42e3f81c634['h02386] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c4] =  I0310077d53ae4ed9904df42e3f81c634['h02388] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c5] =  I0310077d53ae4ed9904df42e3f81c634['h0238a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c6] =  I0310077d53ae4ed9904df42e3f81c634['h0238c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c7] =  I0310077d53ae4ed9904df42e3f81c634['h0238e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c8] =  I0310077d53ae4ed9904df42e3f81c634['h02390] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011c9] =  I0310077d53ae4ed9904df42e3f81c634['h02392] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ca] =  I0310077d53ae4ed9904df42e3f81c634['h02394] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011cb] =  I0310077d53ae4ed9904df42e3f81c634['h02396] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011cc] =  I0310077d53ae4ed9904df42e3f81c634['h02398] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011cd] =  I0310077d53ae4ed9904df42e3f81c634['h0239a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ce] =  I0310077d53ae4ed9904df42e3f81c634['h0239c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011cf] =  I0310077d53ae4ed9904df42e3f81c634['h0239e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d0] =  I0310077d53ae4ed9904df42e3f81c634['h023a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d1] =  I0310077d53ae4ed9904df42e3f81c634['h023a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d2] =  I0310077d53ae4ed9904df42e3f81c634['h023a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d3] =  I0310077d53ae4ed9904df42e3f81c634['h023a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d4] =  I0310077d53ae4ed9904df42e3f81c634['h023a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d5] =  I0310077d53ae4ed9904df42e3f81c634['h023aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d6] =  I0310077d53ae4ed9904df42e3f81c634['h023ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d7] =  I0310077d53ae4ed9904df42e3f81c634['h023ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d8] =  I0310077d53ae4ed9904df42e3f81c634['h023b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011d9] =  I0310077d53ae4ed9904df42e3f81c634['h023b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011da] =  I0310077d53ae4ed9904df42e3f81c634['h023b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011db] =  I0310077d53ae4ed9904df42e3f81c634['h023b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011dc] =  I0310077d53ae4ed9904df42e3f81c634['h023b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011dd] =  I0310077d53ae4ed9904df42e3f81c634['h023ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011de] =  I0310077d53ae4ed9904df42e3f81c634['h023bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011df] =  I0310077d53ae4ed9904df42e3f81c634['h023be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e0] =  I0310077d53ae4ed9904df42e3f81c634['h023c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e1] =  I0310077d53ae4ed9904df42e3f81c634['h023c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e2] =  I0310077d53ae4ed9904df42e3f81c634['h023c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e3] =  I0310077d53ae4ed9904df42e3f81c634['h023c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e4] =  I0310077d53ae4ed9904df42e3f81c634['h023c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e5] =  I0310077d53ae4ed9904df42e3f81c634['h023ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e6] =  I0310077d53ae4ed9904df42e3f81c634['h023cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e7] =  I0310077d53ae4ed9904df42e3f81c634['h023ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e8] =  I0310077d53ae4ed9904df42e3f81c634['h023d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011e9] =  I0310077d53ae4ed9904df42e3f81c634['h023d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ea] =  I0310077d53ae4ed9904df42e3f81c634['h023d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011eb] =  I0310077d53ae4ed9904df42e3f81c634['h023d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ec] =  I0310077d53ae4ed9904df42e3f81c634['h023d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ed] =  I0310077d53ae4ed9904df42e3f81c634['h023da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ee] =  I0310077d53ae4ed9904df42e3f81c634['h023dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ef] =  I0310077d53ae4ed9904df42e3f81c634['h023de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f0] =  I0310077d53ae4ed9904df42e3f81c634['h023e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f1] =  I0310077d53ae4ed9904df42e3f81c634['h023e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f2] =  I0310077d53ae4ed9904df42e3f81c634['h023e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f3] =  I0310077d53ae4ed9904df42e3f81c634['h023e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f4] =  I0310077d53ae4ed9904df42e3f81c634['h023e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f5] =  I0310077d53ae4ed9904df42e3f81c634['h023ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f6] =  I0310077d53ae4ed9904df42e3f81c634['h023ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f7] =  I0310077d53ae4ed9904df42e3f81c634['h023ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f8] =  I0310077d53ae4ed9904df42e3f81c634['h023f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011f9] =  I0310077d53ae4ed9904df42e3f81c634['h023f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011fa] =  I0310077d53ae4ed9904df42e3f81c634['h023f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011fb] =  I0310077d53ae4ed9904df42e3f81c634['h023f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011fc] =  I0310077d53ae4ed9904df42e3f81c634['h023f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011fd] =  I0310077d53ae4ed9904df42e3f81c634['h023fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011fe] =  I0310077d53ae4ed9904df42e3f81c634['h023fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h011ff] =  I0310077d53ae4ed9904df42e3f81c634['h023fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01200] =  I0310077d53ae4ed9904df42e3f81c634['h02400] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01201] =  I0310077d53ae4ed9904df42e3f81c634['h02402] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01202] =  I0310077d53ae4ed9904df42e3f81c634['h02404] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01203] =  I0310077d53ae4ed9904df42e3f81c634['h02406] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01204] =  I0310077d53ae4ed9904df42e3f81c634['h02408] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01205] =  I0310077d53ae4ed9904df42e3f81c634['h0240a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01206] =  I0310077d53ae4ed9904df42e3f81c634['h0240c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01207] =  I0310077d53ae4ed9904df42e3f81c634['h0240e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01208] =  I0310077d53ae4ed9904df42e3f81c634['h02410] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01209] =  I0310077d53ae4ed9904df42e3f81c634['h02412] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0120a] =  I0310077d53ae4ed9904df42e3f81c634['h02414] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0120b] =  I0310077d53ae4ed9904df42e3f81c634['h02416] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0120c] =  I0310077d53ae4ed9904df42e3f81c634['h02418] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0120d] =  I0310077d53ae4ed9904df42e3f81c634['h0241a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0120e] =  I0310077d53ae4ed9904df42e3f81c634['h0241c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0120f] =  I0310077d53ae4ed9904df42e3f81c634['h0241e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01210] =  I0310077d53ae4ed9904df42e3f81c634['h02420] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01211] =  I0310077d53ae4ed9904df42e3f81c634['h02422] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01212] =  I0310077d53ae4ed9904df42e3f81c634['h02424] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01213] =  I0310077d53ae4ed9904df42e3f81c634['h02426] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01214] =  I0310077d53ae4ed9904df42e3f81c634['h02428] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01215] =  I0310077d53ae4ed9904df42e3f81c634['h0242a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01216] =  I0310077d53ae4ed9904df42e3f81c634['h0242c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01217] =  I0310077d53ae4ed9904df42e3f81c634['h0242e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01218] =  I0310077d53ae4ed9904df42e3f81c634['h02430] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01219] =  I0310077d53ae4ed9904df42e3f81c634['h02432] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0121a] =  I0310077d53ae4ed9904df42e3f81c634['h02434] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0121b] =  I0310077d53ae4ed9904df42e3f81c634['h02436] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0121c] =  I0310077d53ae4ed9904df42e3f81c634['h02438] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0121d] =  I0310077d53ae4ed9904df42e3f81c634['h0243a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0121e] =  I0310077d53ae4ed9904df42e3f81c634['h0243c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0121f] =  I0310077d53ae4ed9904df42e3f81c634['h0243e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01220] =  I0310077d53ae4ed9904df42e3f81c634['h02440] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01221] =  I0310077d53ae4ed9904df42e3f81c634['h02442] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01222] =  I0310077d53ae4ed9904df42e3f81c634['h02444] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01223] =  I0310077d53ae4ed9904df42e3f81c634['h02446] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01224] =  I0310077d53ae4ed9904df42e3f81c634['h02448] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01225] =  I0310077d53ae4ed9904df42e3f81c634['h0244a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01226] =  I0310077d53ae4ed9904df42e3f81c634['h0244c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01227] =  I0310077d53ae4ed9904df42e3f81c634['h0244e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01228] =  I0310077d53ae4ed9904df42e3f81c634['h02450] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01229] =  I0310077d53ae4ed9904df42e3f81c634['h02452] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0122a] =  I0310077d53ae4ed9904df42e3f81c634['h02454] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0122b] =  I0310077d53ae4ed9904df42e3f81c634['h02456] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0122c] =  I0310077d53ae4ed9904df42e3f81c634['h02458] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0122d] =  I0310077d53ae4ed9904df42e3f81c634['h0245a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0122e] =  I0310077d53ae4ed9904df42e3f81c634['h0245c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0122f] =  I0310077d53ae4ed9904df42e3f81c634['h0245e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01230] =  I0310077d53ae4ed9904df42e3f81c634['h02460] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01231] =  I0310077d53ae4ed9904df42e3f81c634['h02462] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01232] =  I0310077d53ae4ed9904df42e3f81c634['h02464] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01233] =  I0310077d53ae4ed9904df42e3f81c634['h02466] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01234] =  I0310077d53ae4ed9904df42e3f81c634['h02468] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01235] =  I0310077d53ae4ed9904df42e3f81c634['h0246a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01236] =  I0310077d53ae4ed9904df42e3f81c634['h0246c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01237] =  I0310077d53ae4ed9904df42e3f81c634['h0246e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01238] =  I0310077d53ae4ed9904df42e3f81c634['h02470] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01239] =  I0310077d53ae4ed9904df42e3f81c634['h02472] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0123a] =  I0310077d53ae4ed9904df42e3f81c634['h02474] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0123b] =  I0310077d53ae4ed9904df42e3f81c634['h02476] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0123c] =  I0310077d53ae4ed9904df42e3f81c634['h02478] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0123d] =  I0310077d53ae4ed9904df42e3f81c634['h0247a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0123e] =  I0310077d53ae4ed9904df42e3f81c634['h0247c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0123f] =  I0310077d53ae4ed9904df42e3f81c634['h0247e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01240] =  I0310077d53ae4ed9904df42e3f81c634['h02480] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01241] =  I0310077d53ae4ed9904df42e3f81c634['h02482] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01242] =  I0310077d53ae4ed9904df42e3f81c634['h02484] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01243] =  I0310077d53ae4ed9904df42e3f81c634['h02486] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01244] =  I0310077d53ae4ed9904df42e3f81c634['h02488] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01245] =  I0310077d53ae4ed9904df42e3f81c634['h0248a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01246] =  I0310077d53ae4ed9904df42e3f81c634['h0248c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01247] =  I0310077d53ae4ed9904df42e3f81c634['h0248e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01248] =  I0310077d53ae4ed9904df42e3f81c634['h02490] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01249] =  I0310077d53ae4ed9904df42e3f81c634['h02492] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0124a] =  I0310077d53ae4ed9904df42e3f81c634['h02494] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0124b] =  I0310077d53ae4ed9904df42e3f81c634['h02496] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0124c] =  I0310077d53ae4ed9904df42e3f81c634['h02498] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0124d] =  I0310077d53ae4ed9904df42e3f81c634['h0249a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0124e] =  I0310077d53ae4ed9904df42e3f81c634['h0249c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0124f] =  I0310077d53ae4ed9904df42e3f81c634['h0249e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01250] =  I0310077d53ae4ed9904df42e3f81c634['h024a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01251] =  I0310077d53ae4ed9904df42e3f81c634['h024a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01252] =  I0310077d53ae4ed9904df42e3f81c634['h024a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01253] =  I0310077d53ae4ed9904df42e3f81c634['h024a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01254] =  I0310077d53ae4ed9904df42e3f81c634['h024a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01255] =  I0310077d53ae4ed9904df42e3f81c634['h024aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01256] =  I0310077d53ae4ed9904df42e3f81c634['h024ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01257] =  I0310077d53ae4ed9904df42e3f81c634['h024ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01258] =  I0310077d53ae4ed9904df42e3f81c634['h024b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01259] =  I0310077d53ae4ed9904df42e3f81c634['h024b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0125a] =  I0310077d53ae4ed9904df42e3f81c634['h024b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0125b] =  I0310077d53ae4ed9904df42e3f81c634['h024b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0125c] =  I0310077d53ae4ed9904df42e3f81c634['h024b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0125d] =  I0310077d53ae4ed9904df42e3f81c634['h024ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0125e] =  I0310077d53ae4ed9904df42e3f81c634['h024bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0125f] =  I0310077d53ae4ed9904df42e3f81c634['h024be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01260] =  I0310077d53ae4ed9904df42e3f81c634['h024c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01261] =  I0310077d53ae4ed9904df42e3f81c634['h024c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01262] =  I0310077d53ae4ed9904df42e3f81c634['h024c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01263] =  I0310077d53ae4ed9904df42e3f81c634['h024c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01264] =  I0310077d53ae4ed9904df42e3f81c634['h024c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01265] =  I0310077d53ae4ed9904df42e3f81c634['h024ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01266] =  I0310077d53ae4ed9904df42e3f81c634['h024cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01267] =  I0310077d53ae4ed9904df42e3f81c634['h024ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01268] =  I0310077d53ae4ed9904df42e3f81c634['h024d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01269] =  I0310077d53ae4ed9904df42e3f81c634['h024d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0126a] =  I0310077d53ae4ed9904df42e3f81c634['h024d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0126b] =  I0310077d53ae4ed9904df42e3f81c634['h024d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0126c] =  I0310077d53ae4ed9904df42e3f81c634['h024d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0126d] =  I0310077d53ae4ed9904df42e3f81c634['h024da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0126e] =  I0310077d53ae4ed9904df42e3f81c634['h024dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0126f] =  I0310077d53ae4ed9904df42e3f81c634['h024de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01270] =  I0310077d53ae4ed9904df42e3f81c634['h024e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01271] =  I0310077d53ae4ed9904df42e3f81c634['h024e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01272] =  I0310077d53ae4ed9904df42e3f81c634['h024e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01273] =  I0310077d53ae4ed9904df42e3f81c634['h024e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01274] =  I0310077d53ae4ed9904df42e3f81c634['h024e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01275] =  I0310077d53ae4ed9904df42e3f81c634['h024ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01276] =  I0310077d53ae4ed9904df42e3f81c634['h024ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01277] =  I0310077d53ae4ed9904df42e3f81c634['h024ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01278] =  I0310077d53ae4ed9904df42e3f81c634['h024f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01279] =  I0310077d53ae4ed9904df42e3f81c634['h024f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0127a] =  I0310077d53ae4ed9904df42e3f81c634['h024f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0127b] =  I0310077d53ae4ed9904df42e3f81c634['h024f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0127c] =  I0310077d53ae4ed9904df42e3f81c634['h024f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0127d] =  I0310077d53ae4ed9904df42e3f81c634['h024fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0127e] =  I0310077d53ae4ed9904df42e3f81c634['h024fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0127f] =  I0310077d53ae4ed9904df42e3f81c634['h024fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01280] =  I0310077d53ae4ed9904df42e3f81c634['h02500] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01281] =  I0310077d53ae4ed9904df42e3f81c634['h02502] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01282] =  I0310077d53ae4ed9904df42e3f81c634['h02504] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01283] =  I0310077d53ae4ed9904df42e3f81c634['h02506] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01284] =  I0310077d53ae4ed9904df42e3f81c634['h02508] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01285] =  I0310077d53ae4ed9904df42e3f81c634['h0250a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01286] =  I0310077d53ae4ed9904df42e3f81c634['h0250c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01287] =  I0310077d53ae4ed9904df42e3f81c634['h0250e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01288] =  I0310077d53ae4ed9904df42e3f81c634['h02510] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01289] =  I0310077d53ae4ed9904df42e3f81c634['h02512] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0128a] =  I0310077d53ae4ed9904df42e3f81c634['h02514] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0128b] =  I0310077d53ae4ed9904df42e3f81c634['h02516] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0128c] =  I0310077d53ae4ed9904df42e3f81c634['h02518] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0128d] =  I0310077d53ae4ed9904df42e3f81c634['h0251a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0128e] =  I0310077d53ae4ed9904df42e3f81c634['h0251c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0128f] =  I0310077d53ae4ed9904df42e3f81c634['h0251e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01290] =  I0310077d53ae4ed9904df42e3f81c634['h02520] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01291] =  I0310077d53ae4ed9904df42e3f81c634['h02522] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01292] =  I0310077d53ae4ed9904df42e3f81c634['h02524] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01293] =  I0310077d53ae4ed9904df42e3f81c634['h02526] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01294] =  I0310077d53ae4ed9904df42e3f81c634['h02528] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01295] =  I0310077d53ae4ed9904df42e3f81c634['h0252a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01296] =  I0310077d53ae4ed9904df42e3f81c634['h0252c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01297] =  I0310077d53ae4ed9904df42e3f81c634['h0252e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01298] =  I0310077d53ae4ed9904df42e3f81c634['h02530] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01299] =  I0310077d53ae4ed9904df42e3f81c634['h02532] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0129a] =  I0310077d53ae4ed9904df42e3f81c634['h02534] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0129b] =  I0310077d53ae4ed9904df42e3f81c634['h02536] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0129c] =  I0310077d53ae4ed9904df42e3f81c634['h02538] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0129d] =  I0310077d53ae4ed9904df42e3f81c634['h0253a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0129e] =  I0310077d53ae4ed9904df42e3f81c634['h0253c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0129f] =  I0310077d53ae4ed9904df42e3f81c634['h0253e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a0] =  I0310077d53ae4ed9904df42e3f81c634['h02540] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a1] =  I0310077d53ae4ed9904df42e3f81c634['h02542] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a2] =  I0310077d53ae4ed9904df42e3f81c634['h02544] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a3] =  I0310077d53ae4ed9904df42e3f81c634['h02546] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a4] =  I0310077d53ae4ed9904df42e3f81c634['h02548] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a5] =  I0310077d53ae4ed9904df42e3f81c634['h0254a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a6] =  I0310077d53ae4ed9904df42e3f81c634['h0254c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a7] =  I0310077d53ae4ed9904df42e3f81c634['h0254e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a8] =  I0310077d53ae4ed9904df42e3f81c634['h02550] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012a9] =  I0310077d53ae4ed9904df42e3f81c634['h02552] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012aa] =  I0310077d53ae4ed9904df42e3f81c634['h02554] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ab] =  I0310077d53ae4ed9904df42e3f81c634['h02556] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ac] =  I0310077d53ae4ed9904df42e3f81c634['h02558] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ad] =  I0310077d53ae4ed9904df42e3f81c634['h0255a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ae] =  I0310077d53ae4ed9904df42e3f81c634['h0255c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012af] =  I0310077d53ae4ed9904df42e3f81c634['h0255e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b0] =  I0310077d53ae4ed9904df42e3f81c634['h02560] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b1] =  I0310077d53ae4ed9904df42e3f81c634['h02562] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b2] =  I0310077d53ae4ed9904df42e3f81c634['h02564] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b3] =  I0310077d53ae4ed9904df42e3f81c634['h02566] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b4] =  I0310077d53ae4ed9904df42e3f81c634['h02568] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b5] =  I0310077d53ae4ed9904df42e3f81c634['h0256a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b6] =  I0310077d53ae4ed9904df42e3f81c634['h0256c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b7] =  I0310077d53ae4ed9904df42e3f81c634['h0256e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b8] =  I0310077d53ae4ed9904df42e3f81c634['h02570] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012b9] =  I0310077d53ae4ed9904df42e3f81c634['h02572] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ba] =  I0310077d53ae4ed9904df42e3f81c634['h02574] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012bb] =  I0310077d53ae4ed9904df42e3f81c634['h02576] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012bc] =  I0310077d53ae4ed9904df42e3f81c634['h02578] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012bd] =  I0310077d53ae4ed9904df42e3f81c634['h0257a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012be] =  I0310077d53ae4ed9904df42e3f81c634['h0257c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012bf] =  I0310077d53ae4ed9904df42e3f81c634['h0257e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c0] =  I0310077d53ae4ed9904df42e3f81c634['h02580] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c1] =  I0310077d53ae4ed9904df42e3f81c634['h02582] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c2] =  I0310077d53ae4ed9904df42e3f81c634['h02584] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c3] =  I0310077d53ae4ed9904df42e3f81c634['h02586] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c4] =  I0310077d53ae4ed9904df42e3f81c634['h02588] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c5] =  I0310077d53ae4ed9904df42e3f81c634['h0258a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c6] =  I0310077d53ae4ed9904df42e3f81c634['h0258c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c7] =  I0310077d53ae4ed9904df42e3f81c634['h0258e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c8] =  I0310077d53ae4ed9904df42e3f81c634['h02590] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012c9] =  I0310077d53ae4ed9904df42e3f81c634['h02592] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ca] =  I0310077d53ae4ed9904df42e3f81c634['h02594] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012cb] =  I0310077d53ae4ed9904df42e3f81c634['h02596] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012cc] =  I0310077d53ae4ed9904df42e3f81c634['h02598] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012cd] =  I0310077d53ae4ed9904df42e3f81c634['h0259a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ce] =  I0310077d53ae4ed9904df42e3f81c634['h0259c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012cf] =  I0310077d53ae4ed9904df42e3f81c634['h0259e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d0] =  I0310077d53ae4ed9904df42e3f81c634['h025a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d1] =  I0310077d53ae4ed9904df42e3f81c634['h025a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d2] =  I0310077d53ae4ed9904df42e3f81c634['h025a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d3] =  I0310077d53ae4ed9904df42e3f81c634['h025a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d4] =  I0310077d53ae4ed9904df42e3f81c634['h025a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d5] =  I0310077d53ae4ed9904df42e3f81c634['h025aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d6] =  I0310077d53ae4ed9904df42e3f81c634['h025ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d7] =  I0310077d53ae4ed9904df42e3f81c634['h025ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d8] =  I0310077d53ae4ed9904df42e3f81c634['h025b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012d9] =  I0310077d53ae4ed9904df42e3f81c634['h025b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012da] =  I0310077d53ae4ed9904df42e3f81c634['h025b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012db] =  I0310077d53ae4ed9904df42e3f81c634['h025b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012dc] =  I0310077d53ae4ed9904df42e3f81c634['h025b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012dd] =  I0310077d53ae4ed9904df42e3f81c634['h025ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012de] =  I0310077d53ae4ed9904df42e3f81c634['h025bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012df] =  I0310077d53ae4ed9904df42e3f81c634['h025be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e0] =  I0310077d53ae4ed9904df42e3f81c634['h025c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e1] =  I0310077d53ae4ed9904df42e3f81c634['h025c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e2] =  I0310077d53ae4ed9904df42e3f81c634['h025c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e3] =  I0310077d53ae4ed9904df42e3f81c634['h025c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e4] =  I0310077d53ae4ed9904df42e3f81c634['h025c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e5] =  I0310077d53ae4ed9904df42e3f81c634['h025ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e6] =  I0310077d53ae4ed9904df42e3f81c634['h025cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e7] =  I0310077d53ae4ed9904df42e3f81c634['h025ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e8] =  I0310077d53ae4ed9904df42e3f81c634['h025d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012e9] =  I0310077d53ae4ed9904df42e3f81c634['h025d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ea] =  I0310077d53ae4ed9904df42e3f81c634['h025d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012eb] =  I0310077d53ae4ed9904df42e3f81c634['h025d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ec] =  I0310077d53ae4ed9904df42e3f81c634['h025d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ed] =  I0310077d53ae4ed9904df42e3f81c634['h025da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ee] =  I0310077d53ae4ed9904df42e3f81c634['h025dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ef] =  I0310077d53ae4ed9904df42e3f81c634['h025de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f0] =  I0310077d53ae4ed9904df42e3f81c634['h025e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f1] =  I0310077d53ae4ed9904df42e3f81c634['h025e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f2] =  I0310077d53ae4ed9904df42e3f81c634['h025e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f3] =  I0310077d53ae4ed9904df42e3f81c634['h025e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f4] =  I0310077d53ae4ed9904df42e3f81c634['h025e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f5] =  I0310077d53ae4ed9904df42e3f81c634['h025ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f6] =  I0310077d53ae4ed9904df42e3f81c634['h025ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f7] =  I0310077d53ae4ed9904df42e3f81c634['h025ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f8] =  I0310077d53ae4ed9904df42e3f81c634['h025f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012f9] =  I0310077d53ae4ed9904df42e3f81c634['h025f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012fa] =  I0310077d53ae4ed9904df42e3f81c634['h025f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012fb] =  I0310077d53ae4ed9904df42e3f81c634['h025f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012fc] =  I0310077d53ae4ed9904df42e3f81c634['h025f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012fd] =  I0310077d53ae4ed9904df42e3f81c634['h025fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012fe] =  I0310077d53ae4ed9904df42e3f81c634['h025fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h012ff] =  I0310077d53ae4ed9904df42e3f81c634['h025fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01300] =  I0310077d53ae4ed9904df42e3f81c634['h02600] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01301] =  I0310077d53ae4ed9904df42e3f81c634['h02602] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01302] =  I0310077d53ae4ed9904df42e3f81c634['h02604] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01303] =  I0310077d53ae4ed9904df42e3f81c634['h02606] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01304] =  I0310077d53ae4ed9904df42e3f81c634['h02608] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01305] =  I0310077d53ae4ed9904df42e3f81c634['h0260a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01306] =  I0310077d53ae4ed9904df42e3f81c634['h0260c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01307] =  I0310077d53ae4ed9904df42e3f81c634['h0260e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01308] =  I0310077d53ae4ed9904df42e3f81c634['h02610] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01309] =  I0310077d53ae4ed9904df42e3f81c634['h02612] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0130a] =  I0310077d53ae4ed9904df42e3f81c634['h02614] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0130b] =  I0310077d53ae4ed9904df42e3f81c634['h02616] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0130c] =  I0310077d53ae4ed9904df42e3f81c634['h02618] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0130d] =  I0310077d53ae4ed9904df42e3f81c634['h0261a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0130e] =  I0310077d53ae4ed9904df42e3f81c634['h0261c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0130f] =  I0310077d53ae4ed9904df42e3f81c634['h0261e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01310] =  I0310077d53ae4ed9904df42e3f81c634['h02620] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01311] =  I0310077d53ae4ed9904df42e3f81c634['h02622] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01312] =  I0310077d53ae4ed9904df42e3f81c634['h02624] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01313] =  I0310077d53ae4ed9904df42e3f81c634['h02626] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01314] =  I0310077d53ae4ed9904df42e3f81c634['h02628] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01315] =  I0310077d53ae4ed9904df42e3f81c634['h0262a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01316] =  I0310077d53ae4ed9904df42e3f81c634['h0262c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01317] =  I0310077d53ae4ed9904df42e3f81c634['h0262e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01318] =  I0310077d53ae4ed9904df42e3f81c634['h02630] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01319] =  I0310077d53ae4ed9904df42e3f81c634['h02632] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0131a] =  I0310077d53ae4ed9904df42e3f81c634['h02634] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0131b] =  I0310077d53ae4ed9904df42e3f81c634['h02636] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0131c] =  I0310077d53ae4ed9904df42e3f81c634['h02638] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0131d] =  I0310077d53ae4ed9904df42e3f81c634['h0263a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0131e] =  I0310077d53ae4ed9904df42e3f81c634['h0263c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0131f] =  I0310077d53ae4ed9904df42e3f81c634['h0263e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01320] =  I0310077d53ae4ed9904df42e3f81c634['h02640] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01321] =  I0310077d53ae4ed9904df42e3f81c634['h02642] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01322] =  I0310077d53ae4ed9904df42e3f81c634['h02644] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01323] =  I0310077d53ae4ed9904df42e3f81c634['h02646] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01324] =  I0310077d53ae4ed9904df42e3f81c634['h02648] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01325] =  I0310077d53ae4ed9904df42e3f81c634['h0264a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01326] =  I0310077d53ae4ed9904df42e3f81c634['h0264c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01327] =  I0310077d53ae4ed9904df42e3f81c634['h0264e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01328] =  I0310077d53ae4ed9904df42e3f81c634['h02650] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01329] =  I0310077d53ae4ed9904df42e3f81c634['h02652] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0132a] =  I0310077d53ae4ed9904df42e3f81c634['h02654] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0132b] =  I0310077d53ae4ed9904df42e3f81c634['h02656] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0132c] =  I0310077d53ae4ed9904df42e3f81c634['h02658] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0132d] =  I0310077d53ae4ed9904df42e3f81c634['h0265a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0132e] =  I0310077d53ae4ed9904df42e3f81c634['h0265c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0132f] =  I0310077d53ae4ed9904df42e3f81c634['h0265e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01330] =  I0310077d53ae4ed9904df42e3f81c634['h02660] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01331] =  I0310077d53ae4ed9904df42e3f81c634['h02662] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01332] =  I0310077d53ae4ed9904df42e3f81c634['h02664] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01333] =  I0310077d53ae4ed9904df42e3f81c634['h02666] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01334] =  I0310077d53ae4ed9904df42e3f81c634['h02668] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01335] =  I0310077d53ae4ed9904df42e3f81c634['h0266a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01336] =  I0310077d53ae4ed9904df42e3f81c634['h0266c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01337] =  I0310077d53ae4ed9904df42e3f81c634['h0266e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01338] =  I0310077d53ae4ed9904df42e3f81c634['h02670] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01339] =  I0310077d53ae4ed9904df42e3f81c634['h02672] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0133a] =  I0310077d53ae4ed9904df42e3f81c634['h02674] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0133b] =  I0310077d53ae4ed9904df42e3f81c634['h02676] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0133c] =  I0310077d53ae4ed9904df42e3f81c634['h02678] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0133d] =  I0310077d53ae4ed9904df42e3f81c634['h0267a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0133e] =  I0310077d53ae4ed9904df42e3f81c634['h0267c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0133f] =  I0310077d53ae4ed9904df42e3f81c634['h0267e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01340] =  I0310077d53ae4ed9904df42e3f81c634['h02680] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01341] =  I0310077d53ae4ed9904df42e3f81c634['h02682] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01342] =  I0310077d53ae4ed9904df42e3f81c634['h02684] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01343] =  I0310077d53ae4ed9904df42e3f81c634['h02686] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01344] =  I0310077d53ae4ed9904df42e3f81c634['h02688] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01345] =  I0310077d53ae4ed9904df42e3f81c634['h0268a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01346] =  I0310077d53ae4ed9904df42e3f81c634['h0268c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01347] =  I0310077d53ae4ed9904df42e3f81c634['h0268e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01348] =  I0310077d53ae4ed9904df42e3f81c634['h02690] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01349] =  I0310077d53ae4ed9904df42e3f81c634['h02692] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0134a] =  I0310077d53ae4ed9904df42e3f81c634['h02694] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0134b] =  I0310077d53ae4ed9904df42e3f81c634['h02696] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0134c] =  I0310077d53ae4ed9904df42e3f81c634['h02698] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0134d] =  I0310077d53ae4ed9904df42e3f81c634['h0269a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0134e] =  I0310077d53ae4ed9904df42e3f81c634['h0269c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0134f] =  I0310077d53ae4ed9904df42e3f81c634['h0269e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01350] =  I0310077d53ae4ed9904df42e3f81c634['h026a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01351] =  I0310077d53ae4ed9904df42e3f81c634['h026a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01352] =  I0310077d53ae4ed9904df42e3f81c634['h026a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01353] =  I0310077d53ae4ed9904df42e3f81c634['h026a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01354] =  I0310077d53ae4ed9904df42e3f81c634['h026a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01355] =  I0310077d53ae4ed9904df42e3f81c634['h026aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01356] =  I0310077d53ae4ed9904df42e3f81c634['h026ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01357] =  I0310077d53ae4ed9904df42e3f81c634['h026ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01358] =  I0310077d53ae4ed9904df42e3f81c634['h026b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01359] =  I0310077d53ae4ed9904df42e3f81c634['h026b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0135a] =  I0310077d53ae4ed9904df42e3f81c634['h026b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0135b] =  I0310077d53ae4ed9904df42e3f81c634['h026b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0135c] =  I0310077d53ae4ed9904df42e3f81c634['h026b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0135d] =  I0310077d53ae4ed9904df42e3f81c634['h026ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0135e] =  I0310077d53ae4ed9904df42e3f81c634['h026bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0135f] =  I0310077d53ae4ed9904df42e3f81c634['h026be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01360] =  I0310077d53ae4ed9904df42e3f81c634['h026c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01361] =  I0310077d53ae4ed9904df42e3f81c634['h026c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01362] =  I0310077d53ae4ed9904df42e3f81c634['h026c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01363] =  I0310077d53ae4ed9904df42e3f81c634['h026c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01364] =  I0310077d53ae4ed9904df42e3f81c634['h026c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01365] =  I0310077d53ae4ed9904df42e3f81c634['h026ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01366] =  I0310077d53ae4ed9904df42e3f81c634['h026cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01367] =  I0310077d53ae4ed9904df42e3f81c634['h026ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01368] =  I0310077d53ae4ed9904df42e3f81c634['h026d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01369] =  I0310077d53ae4ed9904df42e3f81c634['h026d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0136a] =  I0310077d53ae4ed9904df42e3f81c634['h026d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0136b] =  I0310077d53ae4ed9904df42e3f81c634['h026d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0136c] =  I0310077d53ae4ed9904df42e3f81c634['h026d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0136d] =  I0310077d53ae4ed9904df42e3f81c634['h026da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0136e] =  I0310077d53ae4ed9904df42e3f81c634['h026dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0136f] =  I0310077d53ae4ed9904df42e3f81c634['h026de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01370] =  I0310077d53ae4ed9904df42e3f81c634['h026e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01371] =  I0310077d53ae4ed9904df42e3f81c634['h026e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01372] =  I0310077d53ae4ed9904df42e3f81c634['h026e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01373] =  I0310077d53ae4ed9904df42e3f81c634['h026e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01374] =  I0310077d53ae4ed9904df42e3f81c634['h026e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01375] =  I0310077d53ae4ed9904df42e3f81c634['h026ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01376] =  I0310077d53ae4ed9904df42e3f81c634['h026ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01377] =  I0310077d53ae4ed9904df42e3f81c634['h026ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01378] =  I0310077d53ae4ed9904df42e3f81c634['h026f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01379] =  I0310077d53ae4ed9904df42e3f81c634['h026f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0137a] =  I0310077d53ae4ed9904df42e3f81c634['h026f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0137b] =  I0310077d53ae4ed9904df42e3f81c634['h026f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0137c] =  I0310077d53ae4ed9904df42e3f81c634['h026f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0137d] =  I0310077d53ae4ed9904df42e3f81c634['h026fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0137e] =  I0310077d53ae4ed9904df42e3f81c634['h026fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0137f] =  I0310077d53ae4ed9904df42e3f81c634['h026fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01380] =  I0310077d53ae4ed9904df42e3f81c634['h02700] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01381] =  I0310077d53ae4ed9904df42e3f81c634['h02702] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01382] =  I0310077d53ae4ed9904df42e3f81c634['h02704] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01383] =  I0310077d53ae4ed9904df42e3f81c634['h02706] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01384] =  I0310077d53ae4ed9904df42e3f81c634['h02708] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01385] =  I0310077d53ae4ed9904df42e3f81c634['h0270a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01386] =  I0310077d53ae4ed9904df42e3f81c634['h0270c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01387] =  I0310077d53ae4ed9904df42e3f81c634['h0270e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01388] =  I0310077d53ae4ed9904df42e3f81c634['h02710] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01389] =  I0310077d53ae4ed9904df42e3f81c634['h02712] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0138a] =  I0310077d53ae4ed9904df42e3f81c634['h02714] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0138b] =  I0310077d53ae4ed9904df42e3f81c634['h02716] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0138c] =  I0310077d53ae4ed9904df42e3f81c634['h02718] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0138d] =  I0310077d53ae4ed9904df42e3f81c634['h0271a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0138e] =  I0310077d53ae4ed9904df42e3f81c634['h0271c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0138f] =  I0310077d53ae4ed9904df42e3f81c634['h0271e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01390] =  I0310077d53ae4ed9904df42e3f81c634['h02720] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01391] =  I0310077d53ae4ed9904df42e3f81c634['h02722] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01392] =  I0310077d53ae4ed9904df42e3f81c634['h02724] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01393] =  I0310077d53ae4ed9904df42e3f81c634['h02726] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01394] =  I0310077d53ae4ed9904df42e3f81c634['h02728] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01395] =  I0310077d53ae4ed9904df42e3f81c634['h0272a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01396] =  I0310077d53ae4ed9904df42e3f81c634['h0272c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01397] =  I0310077d53ae4ed9904df42e3f81c634['h0272e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01398] =  I0310077d53ae4ed9904df42e3f81c634['h02730] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01399] =  I0310077d53ae4ed9904df42e3f81c634['h02732] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0139a] =  I0310077d53ae4ed9904df42e3f81c634['h02734] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0139b] =  I0310077d53ae4ed9904df42e3f81c634['h02736] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0139c] =  I0310077d53ae4ed9904df42e3f81c634['h02738] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0139d] =  I0310077d53ae4ed9904df42e3f81c634['h0273a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0139e] =  I0310077d53ae4ed9904df42e3f81c634['h0273c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0139f] =  I0310077d53ae4ed9904df42e3f81c634['h0273e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a0] =  I0310077d53ae4ed9904df42e3f81c634['h02740] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a1] =  I0310077d53ae4ed9904df42e3f81c634['h02742] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a2] =  I0310077d53ae4ed9904df42e3f81c634['h02744] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a3] =  I0310077d53ae4ed9904df42e3f81c634['h02746] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a4] =  I0310077d53ae4ed9904df42e3f81c634['h02748] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a5] =  I0310077d53ae4ed9904df42e3f81c634['h0274a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a6] =  I0310077d53ae4ed9904df42e3f81c634['h0274c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a7] =  I0310077d53ae4ed9904df42e3f81c634['h0274e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a8] =  I0310077d53ae4ed9904df42e3f81c634['h02750] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013a9] =  I0310077d53ae4ed9904df42e3f81c634['h02752] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013aa] =  I0310077d53ae4ed9904df42e3f81c634['h02754] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ab] =  I0310077d53ae4ed9904df42e3f81c634['h02756] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ac] =  I0310077d53ae4ed9904df42e3f81c634['h02758] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ad] =  I0310077d53ae4ed9904df42e3f81c634['h0275a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ae] =  I0310077d53ae4ed9904df42e3f81c634['h0275c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013af] =  I0310077d53ae4ed9904df42e3f81c634['h0275e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b0] =  I0310077d53ae4ed9904df42e3f81c634['h02760] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b1] =  I0310077d53ae4ed9904df42e3f81c634['h02762] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b2] =  I0310077d53ae4ed9904df42e3f81c634['h02764] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b3] =  I0310077d53ae4ed9904df42e3f81c634['h02766] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b4] =  I0310077d53ae4ed9904df42e3f81c634['h02768] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b5] =  I0310077d53ae4ed9904df42e3f81c634['h0276a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b6] =  I0310077d53ae4ed9904df42e3f81c634['h0276c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b7] =  I0310077d53ae4ed9904df42e3f81c634['h0276e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b8] =  I0310077d53ae4ed9904df42e3f81c634['h02770] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013b9] =  I0310077d53ae4ed9904df42e3f81c634['h02772] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ba] =  I0310077d53ae4ed9904df42e3f81c634['h02774] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013bb] =  I0310077d53ae4ed9904df42e3f81c634['h02776] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013bc] =  I0310077d53ae4ed9904df42e3f81c634['h02778] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013bd] =  I0310077d53ae4ed9904df42e3f81c634['h0277a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013be] =  I0310077d53ae4ed9904df42e3f81c634['h0277c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013bf] =  I0310077d53ae4ed9904df42e3f81c634['h0277e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c0] =  I0310077d53ae4ed9904df42e3f81c634['h02780] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c1] =  I0310077d53ae4ed9904df42e3f81c634['h02782] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c2] =  I0310077d53ae4ed9904df42e3f81c634['h02784] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c3] =  I0310077d53ae4ed9904df42e3f81c634['h02786] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c4] =  I0310077d53ae4ed9904df42e3f81c634['h02788] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c5] =  I0310077d53ae4ed9904df42e3f81c634['h0278a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c6] =  I0310077d53ae4ed9904df42e3f81c634['h0278c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c7] =  I0310077d53ae4ed9904df42e3f81c634['h0278e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c8] =  I0310077d53ae4ed9904df42e3f81c634['h02790] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013c9] =  I0310077d53ae4ed9904df42e3f81c634['h02792] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ca] =  I0310077d53ae4ed9904df42e3f81c634['h02794] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013cb] =  I0310077d53ae4ed9904df42e3f81c634['h02796] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013cc] =  I0310077d53ae4ed9904df42e3f81c634['h02798] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013cd] =  I0310077d53ae4ed9904df42e3f81c634['h0279a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ce] =  I0310077d53ae4ed9904df42e3f81c634['h0279c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013cf] =  I0310077d53ae4ed9904df42e3f81c634['h0279e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d0] =  I0310077d53ae4ed9904df42e3f81c634['h027a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d1] =  I0310077d53ae4ed9904df42e3f81c634['h027a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d2] =  I0310077d53ae4ed9904df42e3f81c634['h027a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d3] =  I0310077d53ae4ed9904df42e3f81c634['h027a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d4] =  I0310077d53ae4ed9904df42e3f81c634['h027a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d5] =  I0310077d53ae4ed9904df42e3f81c634['h027aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d6] =  I0310077d53ae4ed9904df42e3f81c634['h027ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d7] =  I0310077d53ae4ed9904df42e3f81c634['h027ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d8] =  I0310077d53ae4ed9904df42e3f81c634['h027b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013d9] =  I0310077d53ae4ed9904df42e3f81c634['h027b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013da] =  I0310077d53ae4ed9904df42e3f81c634['h027b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013db] =  I0310077d53ae4ed9904df42e3f81c634['h027b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013dc] =  I0310077d53ae4ed9904df42e3f81c634['h027b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013dd] =  I0310077d53ae4ed9904df42e3f81c634['h027ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013de] =  I0310077d53ae4ed9904df42e3f81c634['h027bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013df] =  I0310077d53ae4ed9904df42e3f81c634['h027be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e0] =  I0310077d53ae4ed9904df42e3f81c634['h027c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e1] =  I0310077d53ae4ed9904df42e3f81c634['h027c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e2] =  I0310077d53ae4ed9904df42e3f81c634['h027c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e3] =  I0310077d53ae4ed9904df42e3f81c634['h027c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e4] =  I0310077d53ae4ed9904df42e3f81c634['h027c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e5] =  I0310077d53ae4ed9904df42e3f81c634['h027ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e6] =  I0310077d53ae4ed9904df42e3f81c634['h027cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e7] =  I0310077d53ae4ed9904df42e3f81c634['h027ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e8] =  I0310077d53ae4ed9904df42e3f81c634['h027d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013e9] =  I0310077d53ae4ed9904df42e3f81c634['h027d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ea] =  I0310077d53ae4ed9904df42e3f81c634['h027d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013eb] =  I0310077d53ae4ed9904df42e3f81c634['h027d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ec] =  I0310077d53ae4ed9904df42e3f81c634['h027d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ed] =  I0310077d53ae4ed9904df42e3f81c634['h027da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ee] =  I0310077d53ae4ed9904df42e3f81c634['h027dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ef] =  I0310077d53ae4ed9904df42e3f81c634['h027de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f0] =  I0310077d53ae4ed9904df42e3f81c634['h027e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f1] =  I0310077d53ae4ed9904df42e3f81c634['h027e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f2] =  I0310077d53ae4ed9904df42e3f81c634['h027e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f3] =  I0310077d53ae4ed9904df42e3f81c634['h027e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f4] =  I0310077d53ae4ed9904df42e3f81c634['h027e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f5] =  I0310077d53ae4ed9904df42e3f81c634['h027ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f6] =  I0310077d53ae4ed9904df42e3f81c634['h027ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f7] =  I0310077d53ae4ed9904df42e3f81c634['h027ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f8] =  I0310077d53ae4ed9904df42e3f81c634['h027f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013f9] =  I0310077d53ae4ed9904df42e3f81c634['h027f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013fa] =  I0310077d53ae4ed9904df42e3f81c634['h027f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013fb] =  I0310077d53ae4ed9904df42e3f81c634['h027f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013fc] =  I0310077d53ae4ed9904df42e3f81c634['h027f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013fd] =  I0310077d53ae4ed9904df42e3f81c634['h027fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013fe] =  I0310077d53ae4ed9904df42e3f81c634['h027fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h013ff] =  I0310077d53ae4ed9904df42e3f81c634['h027fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01400] =  I0310077d53ae4ed9904df42e3f81c634['h02800] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01401] =  I0310077d53ae4ed9904df42e3f81c634['h02802] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01402] =  I0310077d53ae4ed9904df42e3f81c634['h02804] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01403] =  I0310077d53ae4ed9904df42e3f81c634['h02806] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01404] =  I0310077d53ae4ed9904df42e3f81c634['h02808] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01405] =  I0310077d53ae4ed9904df42e3f81c634['h0280a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01406] =  I0310077d53ae4ed9904df42e3f81c634['h0280c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01407] =  I0310077d53ae4ed9904df42e3f81c634['h0280e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01408] =  I0310077d53ae4ed9904df42e3f81c634['h02810] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01409] =  I0310077d53ae4ed9904df42e3f81c634['h02812] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0140a] =  I0310077d53ae4ed9904df42e3f81c634['h02814] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0140b] =  I0310077d53ae4ed9904df42e3f81c634['h02816] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0140c] =  I0310077d53ae4ed9904df42e3f81c634['h02818] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0140d] =  I0310077d53ae4ed9904df42e3f81c634['h0281a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0140e] =  I0310077d53ae4ed9904df42e3f81c634['h0281c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0140f] =  I0310077d53ae4ed9904df42e3f81c634['h0281e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01410] =  I0310077d53ae4ed9904df42e3f81c634['h02820] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01411] =  I0310077d53ae4ed9904df42e3f81c634['h02822] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01412] =  I0310077d53ae4ed9904df42e3f81c634['h02824] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01413] =  I0310077d53ae4ed9904df42e3f81c634['h02826] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01414] =  I0310077d53ae4ed9904df42e3f81c634['h02828] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01415] =  I0310077d53ae4ed9904df42e3f81c634['h0282a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01416] =  I0310077d53ae4ed9904df42e3f81c634['h0282c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01417] =  I0310077d53ae4ed9904df42e3f81c634['h0282e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01418] =  I0310077d53ae4ed9904df42e3f81c634['h02830] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01419] =  I0310077d53ae4ed9904df42e3f81c634['h02832] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0141a] =  I0310077d53ae4ed9904df42e3f81c634['h02834] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0141b] =  I0310077d53ae4ed9904df42e3f81c634['h02836] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0141c] =  I0310077d53ae4ed9904df42e3f81c634['h02838] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0141d] =  I0310077d53ae4ed9904df42e3f81c634['h0283a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0141e] =  I0310077d53ae4ed9904df42e3f81c634['h0283c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0141f] =  I0310077d53ae4ed9904df42e3f81c634['h0283e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01420] =  I0310077d53ae4ed9904df42e3f81c634['h02840] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01421] =  I0310077d53ae4ed9904df42e3f81c634['h02842] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01422] =  I0310077d53ae4ed9904df42e3f81c634['h02844] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01423] =  I0310077d53ae4ed9904df42e3f81c634['h02846] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01424] =  I0310077d53ae4ed9904df42e3f81c634['h02848] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01425] =  I0310077d53ae4ed9904df42e3f81c634['h0284a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01426] =  I0310077d53ae4ed9904df42e3f81c634['h0284c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01427] =  I0310077d53ae4ed9904df42e3f81c634['h0284e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01428] =  I0310077d53ae4ed9904df42e3f81c634['h02850] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01429] =  I0310077d53ae4ed9904df42e3f81c634['h02852] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0142a] =  I0310077d53ae4ed9904df42e3f81c634['h02854] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0142b] =  I0310077d53ae4ed9904df42e3f81c634['h02856] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0142c] =  I0310077d53ae4ed9904df42e3f81c634['h02858] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0142d] =  I0310077d53ae4ed9904df42e3f81c634['h0285a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0142e] =  I0310077d53ae4ed9904df42e3f81c634['h0285c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0142f] =  I0310077d53ae4ed9904df42e3f81c634['h0285e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01430] =  I0310077d53ae4ed9904df42e3f81c634['h02860] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01431] =  I0310077d53ae4ed9904df42e3f81c634['h02862] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01432] =  I0310077d53ae4ed9904df42e3f81c634['h02864] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01433] =  I0310077d53ae4ed9904df42e3f81c634['h02866] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01434] =  I0310077d53ae4ed9904df42e3f81c634['h02868] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01435] =  I0310077d53ae4ed9904df42e3f81c634['h0286a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01436] =  I0310077d53ae4ed9904df42e3f81c634['h0286c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01437] =  I0310077d53ae4ed9904df42e3f81c634['h0286e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01438] =  I0310077d53ae4ed9904df42e3f81c634['h02870] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01439] =  I0310077d53ae4ed9904df42e3f81c634['h02872] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0143a] =  I0310077d53ae4ed9904df42e3f81c634['h02874] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0143b] =  I0310077d53ae4ed9904df42e3f81c634['h02876] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0143c] =  I0310077d53ae4ed9904df42e3f81c634['h02878] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0143d] =  I0310077d53ae4ed9904df42e3f81c634['h0287a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0143e] =  I0310077d53ae4ed9904df42e3f81c634['h0287c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0143f] =  I0310077d53ae4ed9904df42e3f81c634['h0287e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01440] =  I0310077d53ae4ed9904df42e3f81c634['h02880] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01441] =  I0310077d53ae4ed9904df42e3f81c634['h02882] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01442] =  I0310077d53ae4ed9904df42e3f81c634['h02884] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01443] =  I0310077d53ae4ed9904df42e3f81c634['h02886] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01444] =  I0310077d53ae4ed9904df42e3f81c634['h02888] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01445] =  I0310077d53ae4ed9904df42e3f81c634['h0288a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01446] =  I0310077d53ae4ed9904df42e3f81c634['h0288c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01447] =  I0310077d53ae4ed9904df42e3f81c634['h0288e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01448] =  I0310077d53ae4ed9904df42e3f81c634['h02890] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01449] =  I0310077d53ae4ed9904df42e3f81c634['h02892] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0144a] =  I0310077d53ae4ed9904df42e3f81c634['h02894] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0144b] =  I0310077d53ae4ed9904df42e3f81c634['h02896] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0144c] =  I0310077d53ae4ed9904df42e3f81c634['h02898] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0144d] =  I0310077d53ae4ed9904df42e3f81c634['h0289a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0144e] =  I0310077d53ae4ed9904df42e3f81c634['h0289c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0144f] =  I0310077d53ae4ed9904df42e3f81c634['h0289e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01450] =  I0310077d53ae4ed9904df42e3f81c634['h028a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01451] =  I0310077d53ae4ed9904df42e3f81c634['h028a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01452] =  I0310077d53ae4ed9904df42e3f81c634['h028a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01453] =  I0310077d53ae4ed9904df42e3f81c634['h028a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01454] =  I0310077d53ae4ed9904df42e3f81c634['h028a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01455] =  I0310077d53ae4ed9904df42e3f81c634['h028aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01456] =  I0310077d53ae4ed9904df42e3f81c634['h028ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01457] =  I0310077d53ae4ed9904df42e3f81c634['h028ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01458] =  I0310077d53ae4ed9904df42e3f81c634['h028b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01459] =  I0310077d53ae4ed9904df42e3f81c634['h028b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0145a] =  I0310077d53ae4ed9904df42e3f81c634['h028b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0145b] =  I0310077d53ae4ed9904df42e3f81c634['h028b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0145c] =  I0310077d53ae4ed9904df42e3f81c634['h028b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0145d] =  I0310077d53ae4ed9904df42e3f81c634['h028ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0145e] =  I0310077d53ae4ed9904df42e3f81c634['h028bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0145f] =  I0310077d53ae4ed9904df42e3f81c634['h028be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01460] =  I0310077d53ae4ed9904df42e3f81c634['h028c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01461] =  I0310077d53ae4ed9904df42e3f81c634['h028c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01462] =  I0310077d53ae4ed9904df42e3f81c634['h028c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01463] =  I0310077d53ae4ed9904df42e3f81c634['h028c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01464] =  I0310077d53ae4ed9904df42e3f81c634['h028c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01465] =  I0310077d53ae4ed9904df42e3f81c634['h028ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01466] =  I0310077d53ae4ed9904df42e3f81c634['h028cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01467] =  I0310077d53ae4ed9904df42e3f81c634['h028ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01468] =  I0310077d53ae4ed9904df42e3f81c634['h028d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01469] =  I0310077d53ae4ed9904df42e3f81c634['h028d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0146a] =  I0310077d53ae4ed9904df42e3f81c634['h028d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0146b] =  I0310077d53ae4ed9904df42e3f81c634['h028d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0146c] =  I0310077d53ae4ed9904df42e3f81c634['h028d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0146d] =  I0310077d53ae4ed9904df42e3f81c634['h028da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0146e] =  I0310077d53ae4ed9904df42e3f81c634['h028dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0146f] =  I0310077d53ae4ed9904df42e3f81c634['h028de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01470] =  I0310077d53ae4ed9904df42e3f81c634['h028e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01471] =  I0310077d53ae4ed9904df42e3f81c634['h028e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01472] =  I0310077d53ae4ed9904df42e3f81c634['h028e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01473] =  I0310077d53ae4ed9904df42e3f81c634['h028e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01474] =  I0310077d53ae4ed9904df42e3f81c634['h028e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01475] =  I0310077d53ae4ed9904df42e3f81c634['h028ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01476] =  I0310077d53ae4ed9904df42e3f81c634['h028ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01477] =  I0310077d53ae4ed9904df42e3f81c634['h028ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01478] =  I0310077d53ae4ed9904df42e3f81c634['h028f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01479] =  I0310077d53ae4ed9904df42e3f81c634['h028f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0147a] =  I0310077d53ae4ed9904df42e3f81c634['h028f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0147b] =  I0310077d53ae4ed9904df42e3f81c634['h028f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0147c] =  I0310077d53ae4ed9904df42e3f81c634['h028f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0147d] =  I0310077d53ae4ed9904df42e3f81c634['h028fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0147e] =  I0310077d53ae4ed9904df42e3f81c634['h028fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0147f] =  I0310077d53ae4ed9904df42e3f81c634['h028fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01480] =  I0310077d53ae4ed9904df42e3f81c634['h02900] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01481] =  I0310077d53ae4ed9904df42e3f81c634['h02902] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01482] =  I0310077d53ae4ed9904df42e3f81c634['h02904] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01483] =  I0310077d53ae4ed9904df42e3f81c634['h02906] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01484] =  I0310077d53ae4ed9904df42e3f81c634['h02908] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01485] =  I0310077d53ae4ed9904df42e3f81c634['h0290a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01486] =  I0310077d53ae4ed9904df42e3f81c634['h0290c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01487] =  I0310077d53ae4ed9904df42e3f81c634['h0290e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01488] =  I0310077d53ae4ed9904df42e3f81c634['h02910] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01489] =  I0310077d53ae4ed9904df42e3f81c634['h02912] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0148a] =  I0310077d53ae4ed9904df42e3f81c634['h02914] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0148b] =  I0310077d53ae4ed9904df42e3f81c634['h02916] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0148c] =  I0310077d53ae4ed9904df42e3f81c634['h02918] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0148d] =  I0310077d53ae4ed9904df42e3f81c634['h0291a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0148e] =  I0310077d53ae4ed9904df42e3f81c634['h0291c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0148f] =  I0310077d53ae4ed9904df42e3f81c634['h0291e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01490] =  I0310077d53ae4ed9904df42e3f81c634['h02920] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01491] =  I0310077d53ae4ed9904df42e3f81c634['h02922] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01492] =  I0310077d53ae4ed9904df42e3f81c634['h02924] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01493] =  I0310077d53ae4ed9904df42e3f81c634['h02926] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01494] =  I0310077d53ae4ed9904df42e3f81c634['h02928] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01495] =  I0310077d53ae4ed9904df42e3f81c634['h0292a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01496] =  I0310077d53ae4ed9904df42e3f81c634['h0292c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01497] =  I0310077d53ae4ed9904df42e3f81c634['h0292e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01498] =  I0310077d53ae4ed9904df42e3f81c634['h02930] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01499] =  I0310077d53ae4ed9904df42e3f81c634['h02932] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0149a] =  I0310077d53ae4ed9904df42e3f81c634['h02934] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0149b] =  I0310077d53ae4ed9904df42e3f81c634['h02936] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0149c] =  I0310077d53ae4ed9904df42e3f81c634['h02938] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0149d] =  I0310077d53ae4ed9904df42e3f81c634['h0293a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0149e] =  I0310077d53ae4ed9904df42e3f81c634['h0293c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0149f] =  I0310077d53ae4ed9904df42e3f81c634['h0293e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a0] =  I0310077d53ae4ed9904df42e3f81c634['h02940] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a1] =  I0310077d53ae4ed9904df42e3f81c634['h02942] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a2] =  I0310077d53ae4ed9904df42e3f81c634['h02944] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a3] =  I0310077d53ae4ed9904df42e3f81c634['h02946] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a4] =  I0310077d53ae4ed9904df42e3f81c634['h02948] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a5] =  I0310077d53ae4ed9904df42e3f81c634['h0294a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a6] =  I0310077d53ae4ed9904df42e3f81c634['h0294c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a7] =  I0310077d53ae4ed9904df42e3f81c634['h0294e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a8] =  I0310077d53ae4ed9904df42e3f81c634['h02950] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014a9] =  I0310077d53ae4ed9904df42e3f81c634['h02952] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014aa] =  I0310077d53ae4ed9904df42e3f81c634['h02954] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ab] =  I0310077d53ae4ed9904df42e3f81c634['h02956] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ac] =  I0310077d53ae4ed9904df42e3f81c634['h02958] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ad] =  I0310077d53ae4ed9904df42e3f81c634['h0295a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ae] =  I0310077d53ae4ed9904df42e3f81c634['h0295c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014af] =  I0310077d53ae4ed9904df42e3f81c634['h0295e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b0] =  I0310077d53ae4ed9904df42e3f81c634['h02960] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b1] =  I0310077d53ae4ed9904df42e3f81c634['h02962] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b2] =  I0310077d53ae4ed9904df42e3f81c634['h02964] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b3] =  I0310077d53ae4ed9904df42e3f81c634['h02966] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b4] =  I0310077d53ae4ed9904df42e3f81c634['h02968] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b5] =  I0310077d53ae4ed9904df42e3f81c634['h0296a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b6] =  I0310077d53ae4ed9904df42e3f81c634['h0296c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b7] =  I0310077d53ae4ed9904df42e3f81c634['h0296e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b8] =  I0310077d53ae4ed9904df42e3f81c634['h02970] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014b9] =  I0310077d53ae4ed9904df42e3f81c634['h02972] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ba] =  I0310077d53ae4ed9904df42e3f81c634['h02974] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014bb] =  I0310077d53ae4ed9904df42e3f81c634['h02976] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014bc] =  I0310077d53ae4ed9904df42e3f81c634['h02978] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014bd] =  I0310077d53ae4ed9904df42e3f81c634['h0297a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014be] =  I0310077d53ae4ed9904df42e3f81c634['h0297c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014bf] =  I0310077d53ae4ed9904df42e3f81c634['h0297e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c0] =  I0310077d53ae4ed9904df42e3f81c634['h02980] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c1] =  I0310077d53ae4ed9904df42e3f81c634['h02982] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c2] =  I0310077d53ae4ed9904df42e3f81c634['h02984] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c3] =  I0310077d53ae4ed9904df42e3f81c634['h02986] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c4] =  I0310077d53ae4ed9904df42e3f81c634['h02988] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c5] =  I0310077d53ae4ed9904df42e3f81c634['h0298a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c6] =  I0310077d53ae4ed9904df42e3f81c634['h0298c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c7] =  I0310077d53ae4ed9904df42e3f81c634['h0298e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c8] =  I0310077d53ae4ed9904df42e3f81c634['h02990] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014c9] =  I0310077d53ae4ed9904df42e3f81c634['h02992] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ca] =  I0310077d53ae4ed9904df42e3f81c634['h02994] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014cb] =  I0310077d53ae4ed9904df42e3f81c634['h02996] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014cc] =  I0310077d53ae4ed9904df42e3f81c634['h02998] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014cd] =  I0310077d53ae4ed9904df42e3f81c634['h0299a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ce] =  I0310077d53ae4ed9904df42e3f81c634['h0299c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014cf] =  I0310077d53ae4ed9904df42e3f81c634['h0299e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d0] =  I0310077d53ae4ed9904df42e3f81c634['h029a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d1] =  I0310077d53ae4ed9904df42e3f81c634['h029a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d2] =  I0310077d53ae4ed9904df42e3f81c634['h029a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d3] =  I0310077d53ae4ed9904df42e3f81c634['h029a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d4] =  I0310077d53ae4ed9904df42e3f81c634['h029a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d5] =  I0310077d53ae4ed9904df42e3f81c634['h029aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d6] =  I0310077d53ae4ed9904df42e3f81c634['h029ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d7] =  I0310077d53ae4ed9904df42e3f81c634['h029ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d8] =  I0310077d53ae4ed9904df42e3f81c634['h029b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014d9] =  I0310077d53ae4ed9904df42e3f81c634['h029b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014da] =  I0310077d53ae4ed9904df42e3f81c634['h029b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014db] =  I0310077d53ae4ed9904df42e3f81c634['h029b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014dc] =  I0310077d53ae4ed9904df42e3f81c634['h029b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014dd] =  I0310077d53ae4ed9904df42e3f81c634['h029ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014de] =  I0310077d53ae4ed9904df42e3f81c634['h029bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014df] =  I0310077d53ae4ed9904df42e3f81c634['h029be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e0] =  I0310077d53ae4ed9904df42e3f81c634['h029c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e1] =  I0310077d53ae4ed9904df42e3f81c634['h029c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e2] =  I0310077d53ae4ed9904df42e3f81c634['h029c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e3] =  I0310077d53ae4ed9904df42e3f81c634['h029c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e4] =  I0310077d53ae4ed9904df42e3f81c634['h029c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e5] =  I0310077d53ae4ed9904df42e3f81c634['h029ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e6] =  I0310077d53ae4ed9904df42e3f81c634['h029cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e7] =  I0310077d53ae4ed9904df42e3f81c634['h029ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e8] =  I0310077d53ae4ed9904df42e3f81c634['h029d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014e9] =  I0310077d53ae4ed9904df42e3f81c634['h029d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ea] =  I0310077d53ae4ed9904df42e3f81c634['h029d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014eb] =  I0310077d53ae4ed9904df42e3f81c634['h029d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ec] =  I0310077d53ae4ed9904df42e3f81c634['h029d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ed] =  I0310077d53ae4ed9904df42e3f81c634['h029da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ee] =  I0310077d53ae4ed9904df42e3f81c634['h029dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ef] =  I0310077d53ae4ed9904df42e3f81c634['h029de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f0] =  I0310077d53ae4ed9904df42e3f81c634['h029e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f1] =  I0310077d53ae4ed9904df42e3f81c634['h029e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f2] =  I0310077d53ae4ed9904df42e3f81c634['h029e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f3] =  I0310077d53ae4ed9904df42e3f81c634['h029e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f4] =  I0310077d53ae4ed9904df42e3f81c634['h029e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f5] =  I0310077d53ae4ed9904df42e3f81c634['h029ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f6] =  I0310077d53ae4ed9904df42e3f81c634['h029ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f7] =  I0310077d53ae4ed9904df42e3f81c634['h029ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f8] =  I0310077d53ae4ed9904df42e3f81c634['h029f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014f9] =  I0310077d53ae4ed9904df42e3f81c634['h029f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014fa] =  I0310077d53ae4ed9904df42e3f81c634['h029f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014fb] =  I0310077d53ae4ed9904df42e3f81c634['h029f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014fc] =  I0310077d53ae4ed9904df42e3f81c634['h029f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014fd] =  I0310077d53ae4ed9904df42e3f81c634['h029fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014fe] =  I0310077d53ae4ed9904df42e3f81c634['h029fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h014ff] =  I0310077d53ae4ed9904df42e3f81c634['h029fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01500] =  I0310077d53ae4ed9904df42e3f81c634['h02a00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01501] =  I0310077d53ae4ed9904df42e3f81c634['h02a02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01502] =  I0310077d53ae4ed9904df42e3f81c634['h02a04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01503] =  I0310077d53ae4ed9904df42e3f81c634['h02a06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01504] =  I0310077d53ae4ed9904df42e3f81c634['h02a08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01505] =  I0310077d53ae4ed9904df42e3f81c634['h02a0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01506] =  I0310077d53ae4ed9904df42e3f81c634['h02a0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01507] =  I0310077d53ae4ed9904df42e3f81c634['h02a0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01508] =  I0310077d53ae4ed9904df42e3f81c634['h02a10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01509] =  I0310077d53ae4ed9904df42e3f81c634['h02a12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0150a] =  I0310077d53ae4ed9904df42e3f81c634['h02a14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0150b] =  I0310077d53ae4ed9904df42e3f81c634['h02a16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0150c] =  I0310077d53ae4ed9904df42e3f81c634['h02a18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0150d] =  I0310077d53ae4ed9904df42e3f81c634['h02a1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0150e] =  I0310077d53ae4ed9904df42e3f81c634['h02a1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0150f] =  I0310077d53ae4ed9904df42e3f81c634['h02a1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01510] =  I0310077d53ae4ed9904df42e3f81c634['h02a20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01511] =  I0310077d53ae4ed9904df42e3f81c634['h02a22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01512] =  I0310077d53ae4ed9904df42e3f81c634['h02a24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01513] =  I0310077d53ae4ed9904df42e3f81c634['h02a26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01514] =  I0310077d53ae4ed9904df42e3f81c634['h02a28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01515] =  I0310077d53ae4ed9904df42e3f81c634['h02a2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01516] =  I0310077d53ae4ed9904df42e3f81c634['h02a2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01517] =  I0310077d53ae4ed9904df42e3f81c634['h02a2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01518] =  I0310077d53ae4ed9904df42e3f81c634['h02a30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01519] =  I0310077d53ae4ed9904df42e3f81c634['h02a32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0151a] =  I0310077d53ae4ed9904df42e3f81c634['h02a34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0151b] =  I0310077d53ae4ed9904df42e3f81c634['h02a36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0151c] =  I0310077d53ae4ed9904df42e3f81c634['h02a38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0151d] =  I0310077d53ae4ed9904df42e3f81c634['h02a3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0151e] =  I0310077d53ae4ed9904df42e3f81c634['h02a3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0151f] =  I0310077d53ae4ed9904df42e3f81c634['h02a3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01520] =  I0310077d53ae4ed9904df42e3f81c634['h02a40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01521] =  I0310077d53ae4ed9904df42e3f81c634['h02a42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01522] =  I0310077d53ae4ed9904df42e3f81c634['h02a44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01523] =  I0310077d53ae4ed9904df42e3f81c634['h02a46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01524] =  I0310077d53ae4ed9904df42e3f81c634['h02a48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01525] =  I0310077d53ae4ed9904df42e3f81c634['h02a4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01526] =  I0310077d53ae4ed9904df42e3f81c634['h02a4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01527] =  I0310077d53ae4ed9904df42e3f81c634['h02a4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01528] =  I0310077d53ae4ed9904df42e3f81c634['h02a50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01529] =  I0310077d53ae4ed9904df42e3f81c634['h02a52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0152a] =  I0310077d53ae4ed9904df42e3f81c634['h02a54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0152b] =  I0310077d53ae4ed9904df42e3f81c634['h02a56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0152c] =  I0310077d53ae4ed9904df42e3f81c634['h02a58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0152d] =  I0310077d53ae4ed9904df42e3f81c634['h02a5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0152e] =  I0310077d53ae4ed9904df42e3f81c634['h02a5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0152f] =  I0310077d53ae4ed9904df42e3f81c634['h02a5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01530] =  I0310077d53ae4ed9904df42e3f81c634['h02a60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01531] =  I0310077d53ae4ed9904df42e3f81c634['h02a62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01532] =  I0310077d53ae4ed9904df42e3f81c634['h02a64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01533] =  I0310077d53ae4ed9904df42e3f81c634['h02a66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01534] =  I0310077d53ae4ed9904df42e3f81c634['h02a68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01535] =  I0310077d53ae4ed9904df42e3f81c634['h02a6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01536] =  I0310077d53ae4ed9904df42e3f81c634['h02a6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01537] =  I0310077d53ae4ed9904df42e3f81c634['h02a6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01538] =  I0310077d53ae4ed9904df42e3f81c634['h02a70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01539] =  I0310077d53ae4ed9904df42e3f81c634['h02a72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0153a] =  I0310077d53ae4ed9904df42e3f81c634['h02a74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0153b] =  I0310077d53ae4ed9904df42e3f81c634['h02a76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0153c] =  I0310077d53ae4ed9904df42e3f81c634['h02a78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0153d] =  I0310077d53ae4ed9904df42e3f81c634['h02a7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0153e] =  I0310077d53ae4ed9904df42e3f81c634['h02a7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0153f] =  I0310077d53ae4ed9904df42e3f81c634['h02a7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01540] =  I0310077d53ae4ed9904df42e3f81c634['h02a80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01541] =  I0310077d53ae4ed9904df42e3f81c634['h02a82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01542] =  I0310077d53ae4ed9904df42e3f81c634['h02a84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01543] =  I0310077d53ae4ed9904df42e3f81c634['h02a86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01544] =  I0310077d53ae4ed9904df42e3f81c634['h02a88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01545] =  I0310077d53ae4ed9904df42e3f81c634['h02a8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01546] =  I0310077d53ae4ed9904df42e3f81c634['h02a8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01547] =  I0310077d53ae4ed9904df42e3f81c634['h02a8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01548] =  I0310077d53ae4ed9904df42e3f81c634['h02a90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01549] =  I0310077d53ae4ed9904df42e3f81c634['h02a92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0154a] =  I0310077d53ae4ed9904df42e3f81c634['h02a94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0154b] =  I0310077d53ae4ed9904df42e3f81c634['h02a96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0154c] =  I0310077d53ae4ed9904df42e3f81c634['h02a98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0154d] =  I0310077d53ae4ed9904df42e3f81c634['h02a9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0154e] =  I0310077d53ae4ed9904df42e3f81c634['h02a9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0154f] =  I0310077d53ae4ed9904df42e3f81c634['h02a9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01550] =  I0310077d53ae4ed9904df42e3f81c634['h02aa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01551] =  I0310077d53ae4ed9904df42e3f81c634['h02aa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01552] =  I0310077d53ae4ed9904df42e3f81c634['h02aa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01553] =  I0310077d53ae4ed9904df42e3f81c634['h02aa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01554] =  I0310077d53ae4ed9904df42e3f81c634['h02aa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01555] =  I0310077d53ae4ed9904df42e3f81c634['h02aaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01556] =  I0310077d53ae4ed9904df42e3f81c634['h02aac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01557] =  I0310077d53ae4ed9904df42e3f81c634['h02aae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01558] =  I0310077d53ae4ed9904df42e3f81c634['h02ab0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01559] =  I0310077d53ae4ed9904df42e3f81c634['h02ab2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0155a] =  I0310077d53ae4ed9904df42e3f81c634['h02ab4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0155b] =  I0310077d53ae4ed9904df42e3f81c634['h02ab6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0155c] =  I0310077d53ae4ed9904df42e3f81c634['h02ab8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0155d] =  I0310077d53ae4ed9904df42e3f81c634['h02aba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0155e] =  I0310077d53ae4ed9904df42e3f81c634['h02abc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0155f] =  I0310077d53ae4ed9904df42e3f81c634['h02abe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01560] =  I0310077d53ae4ed9904df42e3f81c634['h02ac0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01561] =  I0310077d53ae4ed9904df42e3f81c634['h02ac2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01562] =  I0310077d53ae4ed9904df42e3f81c634['h02ac4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01563] =  I0310077d53ae4ed9904df42e3f81c634['h02ac6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01564] =  I0310077d53ae4ed9904df42e3f81c634['h02ac8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01565] =  I0310077d53ae4ed9904df42e3f81c634['h02aca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01566] =  I0310077d53ae4ed9904df42e3f81c634['h02acc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01567] =  I0310077d53ae4ed9904df42e3f81c634['h02ace] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01568] =  I0310077d53ae4ed9904df42e3f81c634['h02ad0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01569] =  I0310077d53ae4ed9904df42e3f81c634['h02ad2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0156a] =  I0310077d53ae4ed9904df42e3f81c634['h02ad4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0156b] =  I0310077d53ae4ed9904df42e3f81c634['h02ad6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0156c] =  I0310077d53ae4ed9904df42e3f81c634['h02ad8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0156d] =  I0310077d53ae4ed9904df42e3f81c634['h02ada] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0156e] =  I0310077d53ae4ed9904df42e3f81c634['h02adc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0156f] =  I0310077d53ae4ed9904df42e3f81c634['h02ade] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01570] =  I0310077d53ae4ed9904df42e3f81c634['h02ae0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01571] =  I0310077d53ae4ed9904df42e3f81c634['h02ae2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01572] =  I0310077d53ae4ed9904df42e3f81c634['h02ae4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01573] =  I0310077d53ae4ed9904df42e3f81c634['h02ae6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01574] =  I0310077d53ae4ed9904df42e3f81c634['h02ae8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01575] =  I0310077d53ae4ed9904df42e3f81c634['h02aea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01576] =  I0310077d53ae4ed9904df42e3f81c634['h02aec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01577] =  I0310077d53ae4ed9904df42e3f81c634['h02aee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01578] =  I0310077d53ae4ed9904df42e3f81c634['h02af0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01579] =  I0310077d53ae4ed9904df42e3f81c634['h02af2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0157a] =  I0310077d53ae4ed9904df42e3f81c634['h02af4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0157b] =  I0310077d53ae4ed9904df42e3f81c634['h02af6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0157c] =  I0310077d53ae4ed9904df42e3f81c634['h02af8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0157d] =  I0310077d53ae4ed9904df42e3f81c634['h02afa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0157e] =  I0310077d53ae4ed9904df42e3f81c634['h02afc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0157f] =  I0310077d53ae4ed9904df42e3f81c634['h02afe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01580] =  I0310077d53ae4ed9904df42e3f81c634['h02b00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01581] =  I0310077d53ae4ed9904df42e3f81c634['h02b02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01582] =  I0310077d53ae4ed9904df42e3f81c634['h02b04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01583] =  I0310077d53ae4ed9904df42e3f81c634['h02b06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01584] =  I0310077d53ae4ed9904df42e3f81c634['h02b08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01585] =  I0310077d53ae4ed9904df42e3f81c634['h02b0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01586] =  I0310077d53ae4ed9904df42e3f81c634['h02b0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01587] =  I0310077d53ae4ed9904df42e3f81c634['h02b0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01588] =  I0310077d53ae4ed9904df42e3f81c634['h02b10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01589] =  I0310077d53ae4ed9904df42e3f81c634['h02b12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0158a] =  I0310077d53ae4ed9904df42e3f81c634['h02b14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0158b] =  I0310077d53ae4ed9904df42e3f81c634['h02b16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0158c] =  I0310077d53ae4ed9904df42e3f81c634['h02b18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0158d] =  I0310077d53ae4ed9904df42e3f81c634['h02b1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0158e] =  I0310077d53ae4ed9904df42e3f81c634['h02b1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0158f] =  I0310077d53ae4ed9904df42e3f81c634['h02b1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01590] =  I0310077d53ae4ed9904df42e3f81c634['h02b20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01591] =  I0310077d53ae4ed9904df42e3f81c634['h02b22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01592] =  I0310077d53ae4ed9904df42e3f81c634['h02b24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01593] =  I0310077d53ae4ed9904df42e3f81c634['h02b26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01594] =  I0310077d53ae4ed9904df42e3f81c634['h02b28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01595] =  I0310077d53ae4ed9904df42e3f81c634['h02b2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01596] =  I0310077d53ae4ed9904df42e3f81c634['h02b2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01597] =  I0310077d53ae4ed9904df42e3f81c634['h02b2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01598] =  I0310077d53ae4ed9904df42e3f81c634['h02b30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01599] =  I0310077d53ae4ed9904df42e3f81c634['h02b32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0159a] =  I0310077d53ae4ed9904df42e3f81c634['h02b34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0159b] =  I0310077d53ae4ed9904df42e3f81c634['h02b36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0159c] =  I0310077d53ae4ed9904df42e3f81c634['h02b38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0159d] =  I0310077d53ae4ed9904df42e3f81c634['h02b3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0159e] =  I0310077d53ae4ed9904df42e3f81c634['h02b3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0159f] =  I0310077d53ae4ed9904df42e3f81c634['h02b3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a0] =  I0310077d53ae4ed9904df42e3f81c634['h02b40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a1] =  I0310077d53ae4ed9904df42e3f81c634['h02b42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a2] =  I0310077d53ae4ed9904df42e3f81c634['h02b44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a3] =  I0310077d53ae4ed9904df42e3f81c634['h02b46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a4] =  I0310077d53ae4ed9904df42e3f81c634['h02b48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a5] =  I0310077d53ae4ed9904df42e3f81c634['h02b4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a6] =  I0310077d53ae4ed9904df42e3f81c634['h02b4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a7] =  I0310077d53ae4ed9904df42e3f81c634['h02b4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a8] =  I0310077d53ae4ed9904df42e3f81c634['h02b50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015a9] =  I0310077d53ae4ed9904df42e3f81c634['h02b52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015aa] =  I0310077d53ae4ed9904df42e3f81c634['h02b54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ab] =  I0310077d53ae4ed9904df42e3f81c634['h02b56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ac] =  I0310077d53ae4ed9904df42e3f81c634['h02b58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ad] =  I0310077d53ae4ed9904df42e3f81c634['h02b5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ae] =  I0310077d53ae4ed9904df42e3f81c634['h02b5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015af] =  I0310077d53ae4ed9904df42e3f81c634['h02b5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b0] =  I0310077d53ae4ed9904df42e3f81c634['h02b60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b1] =  I0310077d53ae4ed9904df42e3f81c634['h02b62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b2] =  I0310077d53ae4ed9904df42e3f81c634['h02b64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b3] =  I0310077d53ae4ed9904df42e3f81c634['h02b66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b4] =  I0310077d53ae4ed9904df42e3f81c634['h02b68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b5] =  I0310077d53ae4ed9904df42e3f81c634['h02b6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b6] =  I0310077d53ae4ed9904df42e3f81c634['h02b6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b7] =  I0310077d53ae4ed9904df42e3f81c634['h02b6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b8] =  I0310077d53ae4ed9904df42e3f81c634['h02b70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015b9] =  I0310077d53ae4ed9904df42e3f81c634['h02b72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ba] =  I0310077d53ae4ed9904df42e3f81c634['h02b74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015bb] =  I0310077d53ae4ed9904df42e3f81c634['h02b76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015bc] =  I0310077d53ae4ed9904df42e3f81c634['h02b78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015bd] =  I0310077d53ae4ed9904df42e3f81c634['h02b7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015be] =  I0310077d53ae4ed9904df42e3f81c634['h02b7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015bf] =  I0310077d53ae4ed9904df42e3f81c634['h02b7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c0] =  I0310077d53ae4ed9904df42e3f81c634['h02b80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c1] =  I0310077d53ae4ed9904df42e3f81c634['h02b82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c2] =  I0310077d53ae4ed9904df42e3f81c634['h02b84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c3] =  I0310077d53ae4ed9904df42e3f81c634['h02b86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c4] =  I0310077d53ae4ed9904df42e3f81c634['h02b88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c5] =  I0310077d53ae4ed9904df42e3f81c634['h02b8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c6] =  I0310077d53ae4ed9904df42e3f81c634['h02b8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c7] =  I0310077d53ae4ed9904df42e3f81c634['h02b8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c8] =  I0310077d53ae4ed9904df42e3f81c634['h02b90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015c9] =  I0310077d53ae4ed9904df42e3f81c634['h02b92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ca] =  I0310077d53ae4ed9904df42e3f81c634['h02b94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015cb] =  I0310077d53ae4ed9904df42e3f81c634['h02b96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015cc] =  I0310077d53ae4ed9904df42e3f81c634['h02b98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015cd] =  I0310077d53ae4ed9904df42e3f81c634['h02b9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ce] =  I0310077d53ae4ed9904df42e3f81c634['h02b9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015cf] =  I0310077d53ae4ed9904df42e3f81c634['h02b9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d0] =  I0310077d53ae4ed9904df42e3f81c634['h02ba0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d1] =  I0310077d53ae4ed9904df42e3f81c634['h02ba2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d2] =  I0310077d53ae4ed9904df42e3f81c634['h02ba4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d3] =  I0310077d53ae4ed9904df42e3f81c634['h02ba6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d4] =  I0310077d53ae4ed9904df42e3f81c634['h02ba8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d5] =  I0310077d53ae4ed9904df42e3f81c634['h02baa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d6] =  I0310077d53ae4ed9904df42e3f81c634['h02bac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d7] =  I0310077d53ae4ed9904df42e3f81c634['h02bae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d8] =  I0310077d53ae4ed9904df42e3f81c634['h02bb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015d9] =  I0310077d53ae4ed9904df42e3f81c634['h02bb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015da] =  I0310077d53ae4ed9904df42e3f81c634['h02bb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015db] =  I0310077d53ae4ed9904df42e3f81c634['h02bb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015dc] =  I0310077d53ae4ed9904df42e3f81c634['h02bb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015dd] =  I0310077d53ae4ed9904df42e3f81c634['h02bba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015de] =  I0310077d53ae4ed9904df42e3f81c634['h02bbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015df] =  I0310077d53ae4ed9904df42e3f81c634['h02bbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e0] =  I0310077d53ae4ed9904df42e3f81c634['h02bc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e1] =  I0310077d53ae4ed9904df42e3f81c634['h02bc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e2] =  I0310077d53ae4ed9904df42e3f81c634['h02bc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e3] =  I0310077d53ae4ed9904df42e3f81c634['h02bc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e4] =  I0310077d53ae4ed9904df42e3f81c634['h02bc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e5] =  I0310077d53ae4ed9904df42e3f81c634['h02bca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e6] =  I0310077d53ae4ed9904df42e3f81c634['h02bcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e7] =  I0310077d53ae4ed9904df42e3f81c634['h02bce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e8] =  I0310077d53ae4ed9904df42e3f81c634['h02bd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015e9] =  I0310077d53ae4ed9904df42e3f81c634['h02bd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ea] =  I0310077d53ae4ed9904df42e3f81c634['h02bd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015eb] =  I0310077d53ae4ed9904df42e3f81c634['h02bd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ec] =  I0310077d53ae4ed9904df42e3f81c634['h02bd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ed] =  I0310077d53ae4ed9904df42e3f81c634['h02bda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ee] =  I0310077d53ae4ed9904df42e3f81c634['h02bdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ef] =  I0310077d53ae4ed9904df42e3f81c634['h02bde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f0] =  I0310077d53ae4ed9904df42e3f81c634['h02be0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f1] =  I0310077d53ae4ed9904df42e3f81c634['h02be2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f2] =  I0310077d53ae4ed9904df42e3f81c634['h02be4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f3] =  I0310077d53ae4ed9904df42e3f81c634['h02be6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f4] =  I0310077d53ae4ed9904df42e3f81c634['h02be8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f5] =  I0310077d53ae4ed9904df42e3f81c634['h02bea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f6] =  I0310077d53ae4ed9904df42e3f81c634['h02bec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f7] =  I0310077d53ae4ed9904df42e3f81c634['h02bee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f8] =  I0310077d53ae4ed9904df42e3f81c634['h02bf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015f9] =  I0310077d53ae4ed9904df42e3f81c634['h02bf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015fa] =  I0310077d53ae4ed9904df42e3f81c634['h02bf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015fb] =  I0310077d53ae4ed9904df42e3f81c634['h02bf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015fc] =  I0310077d53ae4ed9904df42e3f81c634['h02bf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015fd] =  I0310077d53ae4ed9904df42e3f81c634['h02bfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015fe] =  I0310077d53ae4ed9904df42e3f81c634['h02bfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h015ff] =  I0310077d53ae4ed9904df42e3f81c634['h02bfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01600] =  I0310077d53ae4ed9904df42e3f81c634['h02c00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01601] =  I0310077d53ae4ed9904df42e3f81c634['h02c02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01602] =  I0310077d53ae4ed9904df42e3f81c634['h02c04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01603] =  I0310077d53ae4ed9904df42e3f81c634['h02c06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01604] =  I0310077d53ae4ed9904df42e3f81c634['h02c08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01605] =  I0310077d53ae4ed9904df42e3f81c634['h02c0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01606] =  I0310077d53ae4ed9904df42e3f81c634['h02c0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01607] =  I0310077d53ae4ed9904df42e3f81c634['h02c0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01608] =  I0310077d53ae4ed9904df42e3f81c634['h02c10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01609] =  I0310077d53ae4ed9904df42e3f81c634['h02c12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0160a] =  I0310077d53ae4ed9904df42e3f81c634['h02c14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0160b] =  I0310077d53ae4ed9904df42e3f81c634['h02c16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0160c] =  I0310077d53ae4ed9904df42e3f81c634['h02c18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0160d] =  I0310077d53ae4ed9904df42e3f81c634['h02c1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0160e] =  I0310077d53ae4ed9904df42e3f81c634['h02c1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0160f] =  I0310077d53ae4ed9904df42e3f81c634['h02c1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01610] =  I0310077d53ae4ed9904df42e3f81c634['h02c20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01611] =  I0310077d53ae4ed9904df42e3f81c634['h02c22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01612] =  I0310077d53ae4ed9904df42e3f81c634['h02c24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01613] =  I0310077d53ae4ed9904df42e3f81c634['h02c26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01614] =  I0310077d53ae4ed9904df42e3f81c634['h02c28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01615] =  I0310077d53ae4ed9904df42e3f81c634['h02c2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01616] =  I0310077d53ae4ed9904df42e3f81c634['h02c2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01617] =  I0310077d53ae4ed9904df42e3f81c634['h02c2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01618] =  I0310077d53ae4ed9904df42e3f81c634['h02c30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01619] =  I0310077d53ae4ed9904df42e3f81c634['h02c32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0161a] =  I0310077d53ae4ed9904df42e3f81c634['h02c34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0161b] =  I0310077d53ae4ed9904df42e3f81c634['h02c36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0161c] =  I0310077d53ae4ed9904df42e3f81c634['h02c38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0161d] =  I0310077d53ae4ed9904df42e3f81c634['h02c3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0161e] =  I0310077d53ae4ed9904df42e3f81c634['h02c3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0161f] =  I0310077d53ae4ed9904df42e3f81c634['h02c3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01620] =  I0310077d53ae4ed9904df42e3f81c634['h02c40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01621] =  I0310077d53ae4ed9904df42e3f81c634['h02c42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01622] =  I0310077d53ae4ed9904df42e3f81c634['h02c44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01623] =  I0310077d53ae4ed9904df42e3f81c634['h02c46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01624] =  I0310077d53ae4ed9904df42e3f81c634['h02c48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01625] =  I0310077d53ae4ed9904df42e3f81c634['h02c4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01626] =  I0310077d53ae4ed9904df42e3f81c634['h02c4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01627] =  I0310077d53ae4ed9904df42e3f81c634['h02c4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01628] =  I0310077d53ae4ed9904df42e3f81c634['h02c50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01629] =  I0310077d53ae4ed9904df42e3f81c634['h02c52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0162a] =  I0310077d53ae4ed9904df42e3f81c634['h02c54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0162b] =  I0310077d53ae4ed9904df42e3f81c634['h02c56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0162c] =  I0310077d53ae4ed9904df42e3f81c634['h02c58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0162d] =  I0310077d53ae4ed9904df42e3f81c634['h02c5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0162e] =  I0310077d53ae4ed9904df42e3f81c634['h02c5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0162f] =  I0310077d53ae4ed9904df42e3f81c634['h02c5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01630] =  I0310077d53ae4ed9904df42e3f81c634['h02c60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01631] =  I0310077d53ae4ed9904df42e3f81c634['h02c62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01632] =  I0310077d53ae4ed9904df42e3f81c634['h02c64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01633] =  I0310077d53ae4ed9904df42e3f81c634['h02c66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01634] =  I0310077d53ae4ed9904df42e3f81c634['h02c68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01635] =  I0310077d53ae4ed9904df42e3f81c634['h02c6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01636] =  I0310077d53ae4ed9904df42e3f81c634['h02c6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01637] =  I0310077d53ae4ed9904df42e3f81c634['h02c6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01638] =  I0310077d53ae4ed9904df42e3f81c634['h02c70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01639] =  I0310077d53ae4ed9904df42e3f81c634['h02c72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0163a] =  I0310077d53ae4ed9904df42e3f81c634['h02c74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0163b] =  I0310077d53ae4ed9904df42e3f81c634['h02c76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0163c] =  I0310077d53ae4ed9904df42e3f81c634['h02c78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0163d] =  I0310077d53ae4ed9904df42e3f81c634['h02c7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0163e] =  I0310077d53ae4ed9904df42e3f81c634['h02c7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0163f] =  I0310077d53ae4ed9904df42e3f81c634['h02c7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01640] =  I0310077d53ae4ed9904df42e3f81c634['h02c80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01641] =  I0310077d53ae4ed9904df42e3f81c634['h02c82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01642] =  I0310077d53ae4ed9904df42e3f81c634['h02c84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01643] =  I0310077d53ae4ed9904df42e3f81c634['h02c86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01644] =  I0310077d53ae4ed9904df42e3f81c634['h02c88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01645] =  I0310077d53ae4ed9904df42e3f81c634['h02c8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01646] =  I0310077d53ae4ed9904df42e3f81c634['h02c8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01647] =  I0310077d53ae4ed9904df42e3f81c634['h02c8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01648] =  I0310077d53ae4ed9904df42e3f81c634['h02c90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01649] =  I0310077d53ae4ed9904df42e3f81c634['h02c92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0164a] =  I0310077d53ae4ed9904df42e3f81c634['h02c94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0164b] =  I0310077d53ae4ed9904df42e3f81c634['h02c96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0164c] =  I0310077d53ae4ed9904df42e3f81c634['h02c98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0164d] =  I0310077d53ae4ed9904df42e3f81c634['h02c9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0164e] =  I0310077d53ae4ed9904df42e3f81c634['h02c9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0164f] =  I0310077d53ae4ed9904df42e3f81c634['h02c9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01650] =  I0310077d53ae4ed9904df42e3f81c634['h02ca0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01651] =  I0310077d53ae4ed9904df42e3f81c634['h02ca2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01652] =  I0310077d53ae4ed9904df42e3f81c634['h02ca4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01653] =  I0310077d53ae4ed9904df42e3f81c634['h02ca6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01654] =  I0310077d53ae4ed9904df42e3f81c634['h02ca8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01655] =  I0310077d53ae4ed9904df42e3f81c634['h02caa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01656] =  I0310077d53ae4ed9904df42e3f81c634['h02cac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01657] =  I0310077d53ae4ed9904df42e3f81c634['h02cae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01658] =  I0310077d53ae4ed9904df42e3f81c634['h02cb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01659] =  I0310077d53ae4ed9904df42e3f81c634['h02cb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0165a] =  I0310077d53ae4ed9904df42e3f81c634['h02cb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0165b] =  I0310077d53ae4ed9904df42e3f81c634['h02cb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0165c] =  I0310077d53ae4ed9904df42e3f81c634['h02cb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0165d] =  I0310077d53ae4ed9904df42e3f81c634['h02cba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0165e] =  I0310077d53ae4ed9904df42e3f81c634['h02cbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0165f] =  I0310077d53ae4ed9904df42e3f81c634['h02cbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01660] =  I0310077d53ae4ed9904df42e3f81c634['h02cc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01661] =  I0310077d53ae4ed9904df42e3f81c634['h02cc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01662] =  I0310077d53ae4ed9904df42e3f81c634['h02cc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01663] =  I0310077d53ae4ed9904df42e3f81c634['h02cc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01664] =  I0310077d53ae4ed9904df42e3f81c634['h02cc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01665] =  I0310077d53ae4ed9904df42e3f81c634['h02cca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01666] =  I0310077d53ae4ed9904df42e3f81c634['h02ccc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01667] =  I0310077d53ae4ed9904df42e3f81c634['h02cce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01668] =  I0310077d53ae4ed9904df42e3f81c634['h02cd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01669] =  I0310077d53ae4ed9904df42e3f81c634['h02cd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0166a] =  I0310077d53ae4ed9904df42e3f81c634['h02cd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0166b] =  I0310077d53ae4ed9904df42e3f81c634['h02cd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0166c] =  I0310077d53ae4ed9904df42e3f81c634['h02cd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0166d] =  I0310077d53ae4ed9904df42e3f81c634['h02cda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0166e] =  I0310077d53ae4ed9904df42e3f81c634['h02cdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0166f] =  I0310077d53ae4ed9904df42e3f81c634['h02cde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01670] =  I0310077d53ae4ed9904df42e3f81c634['h02ce0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01671] =  I0310077d53ae4ed9904df42e3f81c634['h02ce2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01672] =  I0310077d53ae4ed9904df42e3f81c634['h02ce4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01673] =  I0310077d53ae4ed9904df42e3f81c634['h02ce6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01674] =  I0310077d53ae4ed9904df42e3f81c634['h02ce8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01675] =  I0310077d53ae4ed9904df42e3f81c634['h02cea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01676] =  I0310077d53ae4ed9904df42e3f81c634['h02cec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01677] =  I0310077d53ae4ed9904df42e3f81c634['h02cee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01678] =  I0310077d53ae4ed9904df42e3f81c634['h02cf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01679] =  I0310077d53ae4ed9904df42e3f81c634['h02cf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0167a] =  I0310077d53ae4ed9904df42e3f81c634['h02cf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0167b] =  I0310077d53ae4ed9904df42e3f81c634['h02cf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0167c] =  I0310077d53ae4ed9904df42e3f81c634['h02cf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0167d] =  I0310077d53ae4ed9904df42e3f81c634['h02cfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0167e] =  I0310077d53ae4ed9904df42e3f81c634['h02cfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0167f] =  I0310077d53ae4ed9904df42e3f81c634['h02cfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01680] =  I0310077d53ae4ed9904df42e3f81c634['h02d00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01681] =  I0310077d53ae4ed9904df42e3f81c634['h02d02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01682] =  I0310077d53ae4ed9904df42e3f81c634['h02d04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01683] =  I0310077d53ae4ed9904df42e3f81c634['h02d06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01684] =  I0310077d53ae4ed9904df42e3f81c634['h02d08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01685] =  I0310077d53ae4ed9904df42e3f81c634['h02d0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01686] =  I0310077d53ae4ed9904df42e3f81c634['h02d0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01687] =  I0310077d53ae4ed9904df42e3f81c634['h02d0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01688] =  I0310077d53ae4ed9904df42e3f81c634['h02d10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01689] =  I0310077d53ae4ed9904df42e3f81c634['h02d12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0168a] =  I0310077d53ae4ed9904df42e3f81c634['h02d14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0168b] =  I0310077d53ae4ed9904df42e3f81c634['h02d16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0168c] =  I0310077d53ae4ed9904df42e3f81c634['h02d18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0168d] =  I0310077d53ae4ed9904df42e3f81c634['h02d1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0168e] =  I0310077d53ae4ed9904df42e3f81c634['h02d1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0168f] =  I0310077d53ae4ed9904df42e3f81c634['h02d1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01690] =  I0310077d53ae4ed9904df42e3f81c634['h02d20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01691] =  I0310077d53ae4ed9904df42e3f81c634['h02d22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01692] =  I0310077d53ae4ed9904df42e3f81c634['h02d24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01693] =  I0310077d53ae4ed9904df42e3f81c634['h02d26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01694] =  I0310077d53ae4ed9904df42e3f81c634['h02d28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01695] =  I0310077d53ae4ed9904df42e3f81c634['h02d2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01696] =  I0310077d53ae4ed9904df42e3f81c634['h02d2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01697] =  I0310077d53ae4ed9904df42e3f81c634['h02d2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01698] =  I0310077d53ae4ed9904df42e3f81c634['h02d30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01699] =  I0310077d53ae4ed9904df42e3f81c634['h02d32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0169a] =  I0310077d53ae4ed9904df42e3f81c634['h02d34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0169b] =  I0310077d53ae4ed9904df42e3f81c634['h02d36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0169c] =  I0310077d53ae4ed9904df42e3f81c634['h02d38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0169d] =  I0310077d53ae4ed9904df42e3f81c634['h02d3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0169e] =  I0310077d53ae4ed9904df42e3f81c634['h02d3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0169f] =  I0310077d53ae4ed9904df42e3f81c634['h02d3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a0] =  I0310077d53ae4ed9904df42e3f81c634['h02d40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a1] =  I0310077d53ae4ed9904df42e3f81c634['h02d42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a2] =  I0310077d53ae4ed9904df42e3f81c634['h02d44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a3] =  I0310077d53ae4ed9904df42e3f81c634['h02d46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a4] =  I0310077d53ae4ed9904df42e3f81c634['h02d48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a5] =  I0310077d53ae4ed9904df42e3f81c634['h02d4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a6] =  I0310077d53ae4ed9904df42e3f81c634['h02d4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a7] =  I0310077d53ae4ed9904df42e3f81c634['h02d4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a8] =  I0310077d53ae4ed9904df42e3f81c634['h02d50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016a9] =  I0310077d53ae4ed9904df42e3f81c634['h02d52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016aa] =  I0310077d53ae4ed9904df42e3f81c634['h02d54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ab] =  I0310077d53ae4ed9904df42e3f81c634['h02d56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ac] =  I0310077d53ae4ed9904df42e3f81c634['h02d58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ad] =  I0310077d53ae4ed9904df42e3f81c634['h02d5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ae] =  I0310077d53ae4ed9904df42e3f81c634['h02d5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016af] =  I0310077d53ae4ed9904df42e3f81c634['h02d5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b0] =  I0310077d53ae4ed9904df42e3f81c634['h02d60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b1] =  I0310077d53ae4ed9904df42e3f81c634['h02d62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b2] =  I0310077d53ae4ed9904df42e3f81c634['h02d64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b3] =  I0310077d53ae4ed9904df42e3f81c634['h02d66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b4] =  I0310077d53ae4ed9904df42e3f81c634['h02d68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b5] =  I0310077d53ae4ed9904df42e3f81c634['h02d6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b6] =  I0310077d53ae4ed9904df42e3f81c634['h02d6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b7] =  I0310077d53ae4ed9904df42e3f81c634['h02d6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b8] =  I0310077d53ae4ed9904df42e3f81c634['h02d70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016b9] =  I0310077d53ae4ed9904df42e3f81c634['h02d72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ba] =  I0310077d53ae4ed9904df42e3f81c634['h02d74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016bb] =  I0310077d53ae4ed9904df42e3f81c634['h02d76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016bc] =  I0310077d53ae4ed9904df42e3f81c634['h02d78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016bd] =  I0310077d53ae4ed9904df42e3f81c634['h02d7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016be] =  I0310077d53ae4ed9904df42e3f81c634['h02d7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016bf] =  I0310077d53ae4ed9904df42e3f81c634['h02d7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c0] =  I0310077d53ae4ed9904df42e3f81c634['h02d80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c1] =  I0310077d53ae4ed9904df42e3f81c634['h02d82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c2] =  I0310077d53ae4ed9904df42e3f81c634['h02d84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c3] =  I0310077d53ae4ed9904df42e3f81c634['h02d86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c4] =  I0310077d53ae4ed9904df42e3f81c634['h02d88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c5] =  I0310077d53ae4ed9904df42e3f81c634['h02d8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c6] =  I0310077d53ae4ed9904df42e3f81c634['h02d8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c7] =  I0310077d53ae4ed9904df42e3f81c634['h02d8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c8] =  I0310077d53ae4ed9904df42e3f81c634['h02d90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016c9] =  I0310077d53ae4ed9904df42e3f81c634['h02d92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ca] =  I0310077d53ae4ed9904df42e3f81c634['h02d94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016cb] =  I0310077d53ae4ed9904df42e3f81c634['h02d96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016cc] =  I0310077d53ae4ed9904df42e3f81c634['h02d98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016cd] =  I0310077d53ae4ed9904df42e3f81c634['h02d9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ce] =  I0310077d53ae4ed9904df42e3f81c634['h02d9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016cf] =  I0310077d53ae4ed9904df42e3f81c634['h02d9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d0] =  I0310077d53ae4ed9904df42e3f81c634['h02da0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d1] =  I0310077d53ae4ed9904df42e3f81c634['h02da2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d2] =  I0310077d53ae4ed9904df42e3f81c634['h02da4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d3] =  I0310077d53ae4ed9904df42e3f81c634['h02da6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d4] =  I0310077d53ae4ed9904df42e3f81c634['h02da8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d5] =  I0310077d53ae4ed9904df42e3f81c634['h02daa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d6] =  I0310077d53ae4ed9904df42e3f81c634['h02dac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d7] =  I0310077d53ae4ed9904df42e3f81c634['h02dae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d8] =  I0310077d53ae4ed9904df42e3f81c634['h02db0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016d9] =  I0310077d53ae4ed9904df42e3f81c634['h02db2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016da] =  I0310077d53ae4ed9904df42e3f81c634['h02db4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016db] =  I0310077d53ae4ed9904df42e3f81c634['h02db6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016dc] =  I0310077d53ae4ed9904df42e3f81c634['h02db8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016dd] =  I0310077d53ae4ed9904df42e3f81c634['h02dba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016de] =  I0310077d53ae4ed9904df42e3f81c634['h02dbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016df] =  I0310077d53ae4ed9904df42e3f81c634['h02dbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e0] =  I0310077d53ae4ed9904df42e3f81c634['h02dc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e1] =  I0310077d53ae4ed9904df42e3f81c634['h02dc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e2] =  I0310077d53ae4ed9904df42e3f81c634['h02dc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e3] =  I0310077d53ae4ed9904df42e3f81c634['h02dc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e4] =  I0310077d53ae4ed9904df42e3f81c634['h02dc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e5] =  I0310077d53ae4ed9904df42e3f81c634['h02dca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e6] =  I0310077d53ae4ed9904df42e3f81c634['h02dcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e7] =  I0310077d53ae4ed9904df42e3f81c634['h02dce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e8] =  I0310077d53ae4ed9904df42e3f81c634['h02dd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016e9] =  I0310077d53ae4ed9904df42e3f81c634['h02dd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ea] =  I0310077d53ae4ed9904df42e3f81c634['h02dd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016eb] =  I0310077d53ae4ed9904df42e3f81c634['h02dd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ec] =  I0310077d53ae4ed9904df42e3f81c634['h02dd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ed] =  I0310077d53ae4ed9904df42e3f81c634['h02dda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ee] =  I0310077d53ae4ed9904df42e3f81c634['h02ddc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ef] =  I0310077d53ae4ed9904df42e3f81c634['h02dde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f0] =  I0310077d53ae4ed9904df42e3f81c634['h02de0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f1] =  I0310077d53ae4ed9904df42e3f81c634['h02de2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f2] =  I0310077d53ae4ed9904df42e3f81c634['h02de4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f3] =  I0310077d53ae4ed9904df42e3f81c634['h02de6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f4] =  I0310077d53ae4ed9904df42e3f81c634['h02de8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f5] =  I0310077d53ae4ed9904df42e3f81c634['h02dea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f6] =  I0310077d53ae4ed9904df42e3f81c634['h02dec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f7] =  I0310077d53ae4ed9904df42e3f81c634['h02dee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f8] =  I0310077d53ae4ed9904df42e3f81c634['h02df0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016f9] =  I0310077d53ae4ed9904df42e3f81c634['h02df2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016fa] =  I0310077d53ae4ed9904df42e3f81c634['h02df4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016fb] =  I0310077d53ae4ed9904df42e3f81c634['h02df6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016fc] =  I0310077d53ae4ed9904df42e3f81c634['h02df8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016fd] =  I0310077d53ae4ed9904df42e3f81c634['h02dfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016fe] =  I0310077d53ae4ed9904df42e3f81c634['h02dfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h016ff] =  I0310077d53ae4ed9904df42e3f81c634['h02dfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01700] =  I0310077d53ae4ed9904df42e3f81c634['h02e00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01701] =  I0310077d53ae4ed9904df42e3f81c634['h02e02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01702] =  I0310077d53ae4ed9904df42e3f81c634['h02e04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01703] =  I0310077d53ae4ed9904df42e3f81c634['h02e06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01704] =  I0310077d53ae4ed9904df42e3f81c634['h02e08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01705] =  I0310077d53ae4ed9904df42e3f81c634['h02e0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01706] =  I0310077d53ae4ed9904df42e3f81c634['h02e0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01707] =  I0310077d53ae4ed9904df42e3f81c634['h02e0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01708] =  I0310077d53ae4ed9904df42e3f81c634['h02e10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01709] =  I0310077d53ae4ed9904df42e3f81c634['h02e12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0170a] =  I0310077d53ae4ed9904df42e3f81c634['h02e14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0170b] =  I0310077d53ae4ed9904df42e3f81c634['h02e16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0170c] =  I0310077d53ae4ed9904df42e3f81c634['h02e18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0170d] =  I0310077d53ae4ed9904df42e3f81c634['h02e1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0170e] =  I0310077d53ae4ed9904df42e3f81c634['h02e1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0170f] =  I0310077d53ae4ed9904df42e3f81c634['h02e1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01710] =  I0310077d53ae4ed9904df42e3f81c634['h02e20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01711] =  I0310077d53ae4ed9904df42e3f81c634['h02e22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01712] =  I0310077d53ae4ed9904df42e3f81c634['h02e24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01713] =  I0310077d53ae4ed9904df42e3f81c634['h02e26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01714] =  I0310077d53ae4ed9904df42e3f81c634['h02e28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01715] =  I0310077d53ae4ed9904df42e3f81c634['h02e2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01716] =  I0310077d53ae4ed9904df42e3f81c634['h02e2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01717] =  I0310077d53ae4ed9904df42e3f81c634['h02e2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01718] =  I0310077d53ae4ed9904df42e3f81c634['h02e30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01719] =  I0310077d53ae4ed9904df42e3f81c634['h02e32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0171a] =  I0310077d53ae4ed9904df42e3f81c634['h02e34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0171b] =  I0310077d53ae4ed9904df42e3f81c634['h02e36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0171c] =  I0310077d53ae4ed9904df42e3f81c634['h02e38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0171d] =  I0310077d53ae4ed9904df42e3f81c634['h02e3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0171e] =  I0310077d53ae4ed9904df42e3f81c634['h02e3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0171f] =  I0310077d53ae4ed9904df42e3f81c634['h02e3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01720] =  I0310077d53ae4ed9904df42e3f81c634['h02e40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01721] =  I0310077d53ae4ed9904df42e3f81c634['h02e42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01722] =  I0310077d53ae4ed9904df42e3f81c634['h02e44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01723] =  I0310077d53ae4ed9904df42e3f81c634['h02e46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01724] =  I0310077d53ae4ed9904df42e3f81c634['h02e48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01725] =  I0310077d53ae4ed9904df42e3f81c634['h02e4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01726] =  I0310077d53ae4ed9904df42e3f81c634['h02e4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01727] =  I0310077d53ae4ed9904df42e3f81c634['h02e4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01728] =  I0310077d53ae4ed9904df42e3f81c634['h02e50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01729] =  I0310077d53ae4ed9904df42e3f81c634['h02e52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0172a] =  I0310077d53ae4ed9904df42e3f81c634['h02e54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0172b] =  I0310077d53ae4ed9904df42e3f81c634['h02e56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0172c] =  I0310077d53ae4ed9904df42e3f81c634['h02e58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0172d] =  I0310077d53ae4ed9904df42e3f81c634['h02e5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0172e] =  I0310077d53ae4ed9904df42e3f81c634['h02e5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0172f] =  I0310077d53ae4ed9904df42e3f81c634['h02e5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01730] =  I0310077d53ae4ed9904df42e3f81c634['h02e60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01731] =  I0310077d53ae4ed9904df42e3f81c634['h02e62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01732] =  I0310077d53ae4ed9904df42e3f81c634['h02e64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01733] =  I0310077d53ae4ed9904df42e3f81c634['h02e66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01734] =  I0310077d53ae4ed9904df42e3f81c634['h02e68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01735] =  I0310077d53ae4ed9904df42e3f81c634['h02e6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01736] =  I0310077d53ae4ed9904df42e3f81c634['h02e6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01737] =  I0310077d53ae4ed9904df42e3f81c634['h02e6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01738] =  I0310077d53ae4ed9904df42e3f81c634['h02e70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01739] =  I0310077d53ae4ed9904df42e3f81c634['h02e72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0173a] =  I0310077d53ae4ed9904df42e3f81c634['h02e74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0173b] =  I0310077d53ae4ed9904df42e3f81c634['h02e76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0173c] =  I0310077d53ae4ed9904df42e3f81c634['h02e78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0173d] =  I0310077d53ae4ed9904df42e3f81c634['h02e7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0173e] =  I0310077d53ae4ed9904df42e3f81c634['h02e7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0173f] =  I0310077d53ae4ed9904df42e3f81c634['h02e7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01740] =  I0310077d53ae4ed9904df42e3f81c634['h02e80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01741] =  I0310077d53ae4ed9904df42e3f81c634['h02e82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01742] =  I0310077d53ae4ed9904df42e3f81c634['h02e84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01743] =  I0310077d53ae4ed9904df42e3f81c634['h02e86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01744] =  I0310077d53ae4ed9904df42e3f81c634['h02e88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01745] =  I0310077d53ae4ed9904df42e3f81c634['h02e8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01746] =  I0310077d53ae4ed9904df42e3f81c634['h02e8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01747] =  I0310077d53ae4ed9904df42e3f81c634['h02e8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01748] =  I0310077d53ae4ed9904df42e3f81c634['h02e90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01749] =  I0310077d53ae4ed9904df42e3f81c634['h02e92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0174a] =  I0310077d53ae4ed9904df42e3f81c634['h02e94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0174b] =  I0310077d53ae4ed9904df42e3f81c634['h02e96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0174c] =  I0310077d53ae4ed9904df42e3f81c634['h02e98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0174d] =  I0310077d53ae4ed9904df42e3f81c634['h02e9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0174e] =  I0310077d53ae4ed9904df42e3f81c634['h02e9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0174f] =  I0310077d53ae4ed9904df42e3f81c634['h02e9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01750] =  I0310077d53ae4ed9904df42e3f81c634['h02ea0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01751] =  I0310077d53ae4ed9904df42e3f81c634['h02ea2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01752] =  I0310077d53ae4ed9904df42e3f81c634['h02ea4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01753] =  I0310077d53ae4ed9904df42e3f81c634['h02ea6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01754] =  I0310077d53ae4ed9904df42e3f81c634['h02ea8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01755] =  I0310077d53ae4ed9904df42e3f81c634['h02eaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01756] =  I0310077d53ae4ed9904df42e3f81c634['h02eac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01757] =  I0310077d53ae4ed9904df42e3f81c634['h02eae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01758] =  I0310077d53ae4ed9904df42e3f81c634['h02eb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01759] =  I0310077d53ae4ed9904df42e3f81c634['h02eb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0175a] =  I0310077d53ae4ed9904df42e3f81c634['h02eb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0175b] =  I0310077d53ae4ed9904df42e3f81c634['h02eb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0175c] =  I0310077d53ae4ed9904df42e3f81c634['h02eb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0175d] =  I0310077d53ae4ed9904df42e3f81c634['h02eba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0175e] =  I0310077d53ae4ed9904df42e3f81c634['h02ebc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0175f] =  I0310077d53ae4ed9904df42e3f81c634['h02ebe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01760] =  I0310077d53ae4ed9904df42e3f81c634['h02ec0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01761] =  I0310077d53ae4ed9904df42e3f81c634['h02ec2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01762] =  I0310077d53ae4ed9904df42e3f81c634['h02ec4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01763] =  I0310077d53ae4ed9904df42e3f81c634['h02ec6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01764] =  I0310077d53ae4ed9904df42e3f81c634['h02ec8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01765] =  I0310077d53ae4ed9904df42e3f81c634['h02eca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01766] =  I0310077d53ae4ed9904df42e3f81c634['h02ecc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01767] =  I0310077d53ae4ed9904df42e3f81c634['h02ece] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01768] =  I0310077d53ae4ed9904df42e3f81c634['h02ed0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01769] =  I0310077d53ae4ed9904df42e3f81c634['h02ed2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0176a] =  I0310077d53ae4ed9904df42e3f81c634['h02ed4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0176b] =  I0310077d53ae4ed9904df42e3f81c634['h02ed6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0176c] =  I0310077d53ae4ed9904df42e3f81c634['h02ed8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0176d] =  I0310077d53ae4ed9904df42e3f81c634['h02eda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0176e] =  I0310077d53ae4ed9904df42e3f81c634['h02edc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0176f] =  I0310077d53ae4ed9904df42e3f81c634['h02ede] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01770] =  I0310077d53ae4ed9904df42e3f81c634['h02ee0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01771] =  I0310077d53ae4ed9904df42e3f81c634['h02ee2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01772] =  I0310077d53ae4ed9904df42e3f81c634['h02ee4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01773] =  I0310077d53ae4ed9904df42e3f81c634['h02ee6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01774] =  I0310077d53ae4ed9904df42e3f81c634['h02ee8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01775] =  I0310077d53ae4ed9904df42e3f81c634['h02eea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01776] =  I0310077d53ae4ed9904df42e3f81c634['h02eec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01777] =  I0310077d53ae4ed9904df42e3f81c634['h02eee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01778] =  I0310077d53ae4ed9904df42e3f81c634['h02ef0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01779] =  I0310077d53ae4ed9904df42e3f81c634['h02ef2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0177a] =  I0310077d53ae4ed9904df42e3f81c634['h02ef4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0177b] =  I0310077d53ae4ed9904df42e3f81c634['h02ef6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0177c] =  I0310077d53ae4ed9904df42e3f81c634['h02ef8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0177d] =  I0310077d53ae4ed9904df42e3f81c634['h02efa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0177e] =  I0310077d53ae4ed9904df42e3f81c634['h02efc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0177f] =  I0310077d53ae4ed9904df42e3f81c634['h02efe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01780] =  I0310077d53ae4ed9904df42e3f81c634['h02f00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01781] =  I0310077d53ae4ed9904df42e3f81c634['h02f02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01782] =  I0310077d53ae4ed9904df42e3f81c634['h02f04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01783] =  I0310077d53ae4ed9904df42e3f81c634['h02f06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01784] =  I0310077d53ae4ed9904df42e3f81c634['h02f08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01785] =  I0310077d53ae4ed9904df42e3f81c634['h02f0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01786] =  I0310077d53ae4ed9904df42e3f81c634['h02f0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01787] =  I0310077d53ae4ed9904df42e3f81c634['h02f0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01788] =  I0310077d53ae4ed9904df42e3f81c634['h02f10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01789] =  I0310077d53ae4ed9904df42e3f81c634['h02f12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0178a] =  I0310077d53ae4ed9904df42e3f81c634['h02f14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0178b] =  I0310077d53ae4ed9904df42e3f81c634['h02f16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0178c] =  I0310077d53ae4ed9904df42e3f81c634['h02f18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0178d] =  I0310077d53ae4ed9904df42e3f81c634['h02f1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0178e] =  I0310077d53ae4ed9904df42e3f81c634['h02f1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0178f] =  I0310077d53ae4ed9904df42e3f81c634['h02f1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01790] =  I0310077d53ae4ed9904df42e3f81c634['h02f20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01791] =  I0310077d53ae4ed9904df42e3f81c634['h02f22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01792] =  I0310077d53ae4ed9904df42e3f81c634['h02f24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01793] =  I0310077d53ae4ed9904df42e3f81c634['h02f26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01794] =  I0310077d53ae4ed9904df42e3f81c634['h02f28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01795] =  I0310077d53ae4ed9904df42e3f81c634['h02f2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01796] =  I0310077d53ae4ed9904df42e3f81c634['h02f2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01797] =  I0310077d53ae4ed9904df42e3f81c634['h02f2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01798] =  I0310077d53ae4ed9904df42e3f81c634['h02f30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01799] =  I0310077d53ae4ed9904df42e3f81c634['h02f32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0179a] =  I0310077d53ae4ed9904df42e3f81c634['h02f34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0179b] =  I0310077d53ae4ed9904df42e3f81c634['h02f36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0179c] =  I0310077d53ae4ed9904df42e3f81c634['h02f38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0179d] =  I0310077d53ae4ed9904df42e3f81c634['h02f3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0179e] =  I0310077d53ae4ed9904df42e3f81c634['h02f3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0179f] =  I0310077d53ae4ed9904df42e3f81c634['h02f3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a0] =  I0310077d53ae4ed9904df42e3f81c634['h02f40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a1] =  I0310077d53ae4ed9904df42e3f81c634['h02f42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a2] =  I0310077d53ae4ed9904df42e3f81c634['h02f44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a3] =  I0310077d53ae4ed9904df42e3f81c634['h02f46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a4] =  I0310077d53ae4ed9904df42e3f81c634['h02f48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a5] =  I0310077d53ae4ed9904df42e3f81c634['h02f4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a6] =  I0310077d53ae4ed9904df42e3f81c634['h02f4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a7] =  I0310077d53ae4ed9904df42e3f81c634['h02f4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a8] =  I0310077d53ae4ed9904df42e3f81c634['h02f50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017a9] =  I0310077d53ae4ed9904df42e3f81c634['h02f52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017aa] =  I0310077d53ae4ed9904df42e3f81c634['h02f54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ab] =  I0310077d53ae4ed9904df42e3f81c634['h02f56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ac] =  I0310077d53ae4ed9904df42e3f81c634['h02f58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ad] =  I0310077d53ae4ed9904df42e3f81c634['h02f5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ae] =  I0310077d53ae4ed9904df42e3f81c634['h02f5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017af] =  I0310077d53ae4ed9904df42e3f81c634['h02f5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b0] =  I0310077d53ae4ed9904df42e3f81c634['h02f60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b1] =  I0310077d53ae4ed9904df42e3f81c634['h02f62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b2] =  I0310077d53ae4ed9904df42e3f81c634['h02f64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b3] =  I0310077d53ae4ed9904df42e3f81c634['h02f66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b4] =  I0310077d53ae4ed9904df42e3f81c634['h02f68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b5] =  I0310077d53ae4ed9904df42e3f81c634['h02f6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b6] =  I0310077d53ae4ed9904df42e3f81c634['h02f6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b7] =  I0310077d53ae4ed9904df42e3f81c634['h02f6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b8] =  I0310077d53ae4ed9904df42e3f81c634['h02f70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017b9] =  I0310077d53ae4ed9904df42e3f81c634['h02f72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ba] =  I0310077d53ae4ed9904df42e3f81c634['h02f74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017bb] =  I0310077d53ae4ed9904df42e3f81c634['h02f76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017bc] =  I0310077d53ae4ed9904df42e3f81c634['h02f78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017bd] =  I0310077d53ae4ed9904df42e3f81c634['h02f7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017be] =  I0310077d53ae4ed9904df42e3f81c634['h02f7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017bf] =  I0310077d53ae4ed9904df42e3f81c634['h02f7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c0] =  I0310077d53ae4ed9904df42e3f81c634['h02f80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c1] =  I0310077d53ae4ed9904df42e3f81c634['h02f82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c2] =  I0310077d53ae4ed9904df42e3f81c634['h02f84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c3] =  I0310077d53ae4ed9904df42e3f81c634['h02f86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c4] =  I0310077d53ae4ed9904df42e3f81c634['h02f88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c5] =  I0310077d53ae4ed9904df42e3f81c634['h02f8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c6] =  I0310077d53ae4ed9904df42e3f81c634['h02f8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c7] =  I0310077d53ae4ed9904df42e3f81c634['h02f8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c8] =  I0310077d53ae4ed9904df42e3f81c634['h02f90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017c9] =  I0310077d53ae4ed9904df42e3f81c634['h02f92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ca] =  I0310077d53ae4ed9904df42e3f81c634['h02f94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017cb] =  I0310077d53ae4ed9904df42e3f81c634['h02f96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017cc] =  I0310077d53ae4ed9904df42e3f81c634['h02f98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017cd] =  I0310077d53ae4ed9904df42e3f81c634['h02f9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ce] =  I0310077d53ae4ed9904df42e3f81c634['h02f9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017cf] =  I0310077d53ae4ed9904df42e3f81c634['h02f9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d0] =  I0310077d53ae4ed9904df42e3f81c634['h02fa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d1] =  I0310077d53ae4ed9904df42e3f81c634['h02fa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d2] =  I0310077d53ae4ed9904df42e3f81c634['h02fa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d3] =  I0310077d53ae4ed9904df42e3f81c634['h02fa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d4] =  I0310077d53ae4ed9904df42e3f81c634['h02fa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d5] =  I0310077d53ae4ed9904df42e3f81c634['h02faa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d6] =  I0310077d53ae4ed9904df42e3f81c634['h02fac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d7] =  I0310077d53ae4ed9904df42e3f81c634['h02fae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d8] =  I0310077d53ae4ed9904df42e3f81c634['h02fb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017d9] =  I0310077d53ae4ed9904df42e3f81c634['h02fb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017da] =  I0310077d53ae4ed9904df42e3f81c634['h02fb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017db] =  I0310077d53ae4ed9904df42e3f81c634['h02fb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017dc] =  I0310077d53ae4ed9904df42e3f81c634['h02fb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017dd] =  I0310077d53ae4ed9904df42e3f81c634['h02fba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017de] =  I0310077d53ae4ed9904df42e3f81c634['h02fbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017df] =  I0310077d53ae4ed9904df42e3f81c634['h02fbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e0] =  I0310077d53ae4ed9904df42e3f81c634['h02fc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e1] =  I0310077d53ae4ed9904df42e3f81c634['h02fc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e2] =  I0310077d53ae4ed9904df42e3f81c634['h02fc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e3] =  I0310077d53ae4ed9904df42e3f81c634['h02fc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e4] =  I0310077d53ae4ed9904df42e3f81c634['h02fc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e5] =  I0310077d53ae4ed9904df42e3f81c634['h02fca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e6] =  I0310077d53ae4ed9904df42e3f81c634['h02fcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e7] =  I0310077d53ae4ed9904df42e3f81c634['h02fce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e8] =  I0310077d53ae4ed9904df42e3f81c634['h02fd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017e9] =  I0310077d53ae4ed9904df42e3f81c634['h02fd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ea] =  I0310077d53ae4ed9904df42e3f81c634['h02fd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017eb] =  I0310077d53ae4ed9904df42e3f81c634['h02fd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ec] =  I0310077d53ae4ed9904df42e3f81c634['h02fd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ed] =  I0310077d53ae4ed9904df42e3f81c634['h02fda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ee] =  I0310077d53ae4ed9904df42e3f81c634['h02fdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ef] =  I0310077d53ae4ed9904df42e3f81c634['h02fde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f0] =  I0310077d53ae4ed9904df42e3f81c634['h02fe0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f1] =  I0310077d53ae4ed9904df42e3f81c634['h02fe2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f2] =  I0310077d53ae4ed9904df42e3f81c634['h02fe4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f3] =  I0310077d53ae4ed9904df42e3f81c634['h02fe6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f4] =  I0310077d53ae4ed9904df42e3f81c634['h02fe8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f5] =  I0310077d53ae4ed9904df42e3f81c634['h02fea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f6] =  I0310077d53ae4ed9904df42e3f81c634['h02fec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f7] =  I0310077d53ae4ed9904df42e3f81c634['h02fee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f8] =  I0310077d53ae4ed9904df42e3f81c634['h02ff0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017f9] =  I0310077d53ae4ed9904df42e3f81c634['h02ff2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017fa] =  I0310077d53ae4ed9904df42e3f81c634['h02ff4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017fb] =  I0310077d53ae4ed9904df42e3f81c634['h02ff6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017fc] =  I0310077d53ae4ed9904df42e3f81c634['h02ff8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017fd] =  I0310077d53ae4ed9904df42e3f81c634['h02ffa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017fe] =  I0310077d53ae4ed9904df42e3f81c634['h02ffc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h017ff] =  I0310077d53ae4ed9904df42e3f81c634['h02ffe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01800] =  I0310077d53ae4ed9904df42e3f81c634['h03000] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01801] =  I0310077d53ae4ed9904df42e3f81c634['h03002] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01802] =  I0310077d53ae4ed9904df42e3f81c634['h03004] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01803] =  I0310077d53ae4ed9904df42e3f81c634['h03006] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01804] =  I0310077d53ae4ed9904df42e3f81c634['h03008] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01805] =  I0310077d53ae4ed9904df42e3f81c634['h0300a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01806] =  I0310077d53ae4ed9904df42e3f81c634['h0300c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01807] =  I0310077d53ae4ed9904df42e3f81c634['h0300e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01808] =  I0310077d53ae4ed9904df42e3f81c634['h03010] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01809] =  I0310077d53ae4ed9904df42e3f81c634['h03012] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0180a] =  I0310077d53ae4ed9904df42e3f81c634['h03014] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0180b] =  I0310077d53ae4ed9904df42e3f81c634['h03016] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0180c] =  I0310077d53ae4ed9904df42e3f81c634['h03018] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0180d] =  I0310077d53ae4ed9904df42e3f81c634['h0301a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0180e] =  I0310077d53ae4ed9904df42e3f81c634['h0301c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0180f] =  I0310077d53ae4ed9904df42e3f81c634['h0301e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01810] =  I0310077d53ae4ed9904df42e3f81c634['h03020] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01811] =  I0310077d53ae4ed9904df42e3f81c634['h03022] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01812] =  I0310077d53ae4ed9904df42e3f81c634['h03024] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01813] =  I0310077d53ae4ed9904df42e3f81c634['h03026] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01814] =  I0310077d53ae4ed9904df42e3f81c634['h03028] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01815] =  I0310077d53ae4ed9904df42e3f81c634['h0302a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01816] =  I0310077d53ae4ed9904df42e3f81c634['h0302c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01817] =  I0310077d53ae4ed9904df42e3f81c634['h0302e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01818] =  I0310077d53ae4ed9904df42e3f81c634['h03030] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01819] =  I0310077d53ae4ed9904df42e3f81c634['h03032] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0181a] =  I0310077d53ae4ed9904df42e3f81c634['h03034] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0181b] =  I0310077d53ae4ed9904df42e3f81c634['h03036] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0181c] =  I0310077d53ae4ed9904df42e3f81c634['h03038] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0181d] =  I0310077d53ae4ed9904df42e3f81c634['h0303a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0181e] =  I0310077d53ae4ed9904df42e3f81c634['h0303c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0181f] =  I0310077d53ae4ed9904df42e3f81c634['h0303e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01820] =  I0310077d53ae4ed9904df42e3f81c634['h03040] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01821] =  I0310077d53ae4ed9904df42e3f81c634['h03042] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01822] =  I0310077d53ae4ed9904df42e3f81c634['h03044] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01823] =  I0310077d53ae4ed9904df42e3f81c634['h03046] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01824] =  I0310077d53ae4ed9904df42e3f81c634['h03048] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01825] =  I0310077d53ae4ed9904df42e3f81c634['h0304a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01826] =  I0310077d53ae4ed9904df42e3f81c634['h0304c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01827] =  I0310077d53ae4ed9904df42e3f81c634['h0304e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01828] =  I0310077d53ae4ed9904df42e3f81c634['h03050] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01829] =  I0310077d53ae4ed9904df42e3f81c634['h03052] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0182a] =  I0310077d53ae4ed9904df42e3f81c634['h03054] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0182b] =  I0310077d53ae4ed9904df42e3f81c634['h03056] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0182c] =  I0310077d53ae4ed9904df42e3f81c634['h03058] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0182d] =  I0310077d53ae4ed9904df42e3f81c634['h0305a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0182e] =  I0310077d53ae4ed9904df42e3f81c634['h0305c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0182f] =  I0310077d53ae4ed9904df42e3f81c634['h0305e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01830] =  I0310077d53ae4ed9904df42e3f81c634['h03060] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01831] =  I0310077d53ae4ed9904df42e3f81c634['h03062] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01832] =  I0310077d53ae4ed9904df42e3f81c634['h03064] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01833] =  I0310077d53ae4ed9904df42e3f81c634['h03066] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01834] =  I0310077d53ae4ed9904df42e3f81c634['h03068] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01835] =  I0310077d53ae4ed9904df42e3f81c634['h0306a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01836] =  I0310077d53ae4ed9904df42e3f81c634['h0306c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01837] =  I0310077d53ae4ed9904df42e3f81c634['h0306e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01838] =  I0310077d53ae4ed9904df42e3f81c634['h03070] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01839] =  I0310077d53ae4ed9904df42e3f81c634['h03072] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0183a] =  I0310077d53ae4ed9904df42e3f81c634['h03074] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0183b] =  I0310077d53ae4ed9904df42e3f81c634['h03076] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0183c] =  I0310077d53ae4ed9904df42e3f81c634['h03078] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0183d] =  I0310077d53ae4ed9904df42e3f81c634['h0307a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0183e] =  I0310077d53ae4ed9904df42e3f81c634['h0307c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0183f] =  I0310077d53ae4ed9904df42e3f81c634['h0307e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01840] =  I0310077d53ae4ed9904df42e3f81c634['h03080] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01841] =  I0310077d53ae4ed9904df42e3f81c634['h03082] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01842] =  I0310077d53ae4ed9904df42e3f81c634['h03084] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01843] =  I0310077d53ae4ed9904df42e3f81c634['h03086] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01844] =  I0310077d53ae4ed9904df42e3f81c634['h03088] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01845] =  I0310077d53ae4ed9904df42e3f81c634['h0308a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01846] =  I0310077d53ae4ed9904df42e3f81c634['h0308c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01847] =  I0310077d53ae4ed9904df42e3f81c634['h0308e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01848] =  I0310077d53ae4ed9904df42e3f81c634['h03090] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01849] =  I0310077d53ae4ed9904df42e3f81c634['h03092] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0184a] =  I0310077d53ae4ed9904df42e3f81c634['h03094] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0184b] =  I0310077d53ae4ed9904df42e3f81c634['h03096] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0184c] =  I0310077d53ae4ed9904df42e3f81c634['h03098] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0184d] =  I0310077d53ae4ed9904df42e3f81c634['h0309a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0184e] =  I0310077d53ae4ed9904df42e3f81c634['h0309c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0184f] =  I0310077d53ae4ed9904df42e3f81c634['h0309e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01850] =  I0310077d53ae4ed9904df42e3f81c634['h030a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01851] =  I0310077d53ae4ed9904df42e3f81c634['h030a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01852] =  I0310077d53ae4ed9904df42e3f81c634['h030a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01853] =  I0310077d53ae4ed9904df42e3f81c634['h030a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01854] =  I0310077d53ae4ed9904df42e3f81c634['h030a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01855] =  I0310077d53ae4ed9904df42e3f81c634['h030aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01856] =  I0310077d53ae4ed9904df42e3f81c634['h030ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01857] =  I0310077d53ae4ed9904df42e3f81c634['h030ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01858] =  I0310077d53ae4ed9904df42e3f81c634['h030b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01859] =  I0310077d53ae4ed9904df42e3f81c634['h030b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0185a] =  I0310077d53ae4ed9904df42e3f81c634['h030b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0185b] =  I0310077d53ae4ed9904df42e3f81c634['h030b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0185c] =  I0310077d53ae4ed9904df42e3f81c634['h030b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0185d] =  I0310077d53ae4ed9904df42e3f81c634['h030ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0185e] =  I0310077d53ae4ed9904df42e3f81c634['h030bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0185f] =  I0310077d53ae4ed9904df42e3f81c634['h030be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01860] =  I0310077d53ae4ed9904df42e3f81c634['h030c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01861] =  I0310077d53ae4ed9904df42e3f81c634['h030c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01862] =  I0310077d53ae4ed9904df42e3f81c634['h030c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01863] =  I0310077d53ae4ed9904df42e3f81c634['h030c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01864] =  I0310077d53ae4ed9904df42e3f81c634['h030c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01865] =  I0310077d53ae4ed9904df42e3f81c634['h030ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01866] =  I0310077d53ae4ed9904df42e3f81c634['h030cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01867] =  I0310077d53ae4ed9904df42e3f81c634['h030ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01868] =  I0310077d53ae4ed9904df42e3f81c634['h030d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01869] =  I0310077d53ae4ed9904df42e3f81c634['h030d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0186a] =  I0310077d53ae4ed9904df42e3f81c634['h030d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0186b] =  I0310077d53ae4ed9904df42e3f81c634['h030d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0186c] =  I0310077d53ae4ed9904df42e3f81c634['h030d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0186d] =  I0310077d53ae4ed9904df42e3f81c634['h030da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0186e] =  I0310077d53ae4ed9904df42e3f81c634['h030dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0186f] =  I0310077d53ae4ed9904df42e3f81c634['h030de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01870] =  I0310077d53ae4ed9904df42e3f81c634['h030e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01871] =  I0310077d53ae4ed9904df42e3f81c634['h030e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01872] =  I0310077d53ae4ed9904df42e3f81c634['h030e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01873] =  I0310077d53ae4ed9904df42e3f81c634['h030e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01874] =  I0310077d53ae4ed9904df42e3f81c634['h030e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01875] =  I0310077d53ae4ed9904df42e3f81c634['h030ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01876] =  I0310077d53ae4ed9904df42e3f81c634['h030ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01877] =  I0310077d53ae4ed9904df42e3f81c634['h030ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01878] =  I0310077d53ae4ed9904df42e3f81c634['h030f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01879] =  I0310077d53ae4ed9904df42e3f81c634['h030f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0187a] =  I0310077d53ae4ed9904df42e3f81c634['h030f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0187b] =  I0310077d53ae4ed9904df42e3f81c634['h030f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0187c] =  I0310077d53ae4ed9904df42e3f81c634['h030f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0187d] =  I0310077d53ae4ed9904df42e3f81c634['h030fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0187e] =  I0310077d53ae4ed9904df42e3f81c634['h030fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0187f] =  I0310077d53ae4ed9904df42e3f81c634['h030fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01880] =  I0310077d53ae4ed9904df42e3f81c634['h03100] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01881] =  I0310077d53ae4ed9904df42e3f81c634['h03102] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01882] =  I0310077d53ae4ed9904df42e3f81c634['h03104] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01883] =  I0310077d53ae4ed9904df42e3f81c634['h03106] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01884] =  I0310077d53ae4ed9904df42e3f81c634['h03108] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01885] =  I0310077d53ae4ed9904df42e3f81c634['h0310a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01886] =  I0310077d53ae4ed9904df42e3f81c634['h0310c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01887] =  I0310077d53ae4ed9904df42e3f81c634['h0310e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01888] =  I0310077d53ae4ed9904df42e3f81c634['h03110] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01889] =  I0310077d53ae4ed9904df42e3f81c634['h03112] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0188a] =  I0310077d53ae4ed9904df42e3f81c634['h03114] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0188b] =  I0310077d53ae4ed9904df42e3f81c634['h03116] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0188c] =  I0310077d53ae4ed9904df42e3f81c634['h03118] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0188d] =  I0310077d53ae4ed9904df42e3f81c634['h0311a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0188e] =  I0310077d53ae4ed9904df42e3f81c634['h0311c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0188f] =  I0310077d53ae4ed9904df42e3f81c634['h0311e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01890] =  I0310077d53ae4ed9904df42e3f81c634['h03120] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01891] =  I0310077d53ae4ed9904df42e3f81c634['h03122] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01892] =  I0310077d53ae4ed9904df42e3f81c634['h03124] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01893] =  I0310077d53ae4ed9904df42e3f81c634['h03126] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01894] =  I0310077d53ae4ed9904df42e3f81c634['h03128] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01895] =  I0310077d53ae4ed9904df42e3f81c634['h0312a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01896] =  I0310077d53ae4ed9904df42e3f81c634['h0312c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01897] =  I0310077d53ae4ed9904df42e3f81c634['h0312e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01898] =  I0310077d53ae4ed9904df42e3f81c634['h03130] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01899] =  I0310077d53ae4ed9904df42e3f81c634['h03132] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0189a] =  I0310077d53ae4ed9904df42e3f81c634['h03134] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0189b] =  I0310077d53ae4ed9904df42e3f81c634['h03136] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0189c] =  I0310077d53ae4ed9904df42e3f81c634['h03138] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0189d] =  I0310077d53ae4ed9904df42e3f81c634['h0313a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0189e] =  I0310077d53ae4ed9904df42e3f81c634['h0313c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0189f] =  I0310077d53ae4ed9904df42e3f81c634['h0313e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a0] =  I0310077d53ae4ed9904df42e3f81c634['h03140] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a1] =  I0310077d53ae4ed9904df42e3f81c634['h03142] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a2] =  I0310077d53ae4ed9904df42e3f81c634['h03144] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a3] =  I0310077d53ae4ed9904df42e3f81c634['h03146] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a4] =  I0310077d53ae4ed9904df42e3f81c634['h03148] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a5] =  I0310077d53ae4ed9904df42e3f81c634['h0314a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a6] =  I0310077d53ae4ed9904df42e3f81c634['h0314c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a7] =  I0310077d53ae4ed9904df42e3f81c634['h0314e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a8] =  I0310077d53ae4ed9904df42e3f81c634['h03150] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018a9] =  I0310077d53ae4ed9904df42e3f81c634['h03152] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018aa] =  I0310077d53ae4ed9904df42e3f81c634['h03154] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ab] =  I0310077d53ae4ed9904df42e3f81c634['h03156] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ac] =  I0310077d53ae4ed9904df42e3f81c634['h03158] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ad] =  I0310077d53ae4ed9904df42e3f81c634['h0315a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ae] =  I0310077d53ae4ed9904df42e3f81c634['h0315c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018af] =  I0310077d53ae4ed9904df42e3f81c634['h0315e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b0] =  I0310077d53ae4ed9904df42e3f81c634['h03160] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b1] =  I0310077d53ae4ed9904df42e3f81c634['h03162] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b2] =  I0310077d53ae4ed9904df42e3f81c634['h03164] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b3] =  I0310077d53ae4ed9904df42e3f81c634['h03166] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b4] =  I0310077d53ae4ed9904df42e3f81c634['h03168] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b5] =  I0310077d53ae4ed9904df42e3f81c634['h0316a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b6] =  I0310077d53ae4ed9904df42e3f81c634['h0316c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b7] =  I0310077d53ae4ed9904df42e3f81c634['h0316e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b8] =  I0310077d53ae4ed9904df42e3f81c634['h03170] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018b9] =  I0310077d53ae4ed9904df42e3f81c634['h03172] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ba] =  I0310077d53ae4ed9904df42e3f81c634['h03174] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018bb] =  I0310077d53ae4ed9904df42e3f81c634['h03176] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018bc] =  I0310077d53ae4ed9904df42e3f81c634['h03178] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018bd] =  I0310077d53ae4ed9904df42e3f81c634['h0317a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018be] =  I0310077d53ae4ed9904df42e3f81c634['h0317c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018bf] =  I0310077d53ae4ed9904df42e3f81c634['h0317e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c0] =  I0310077d53ae4ed9904df42e3f81c634['h03180] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c1] =  I0310077d53ae4ed9904df42e3f81c634['h03182] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c2] =  I0310077d53ae4ed9904df42e3f81c634['h03184] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c3] =  I0310077d53ae4ed9904df42e3f81c634['h03186] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c4] =  I0310077d53ae4ed9904df42e3f81c634['h03188] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c5] =  I0310077d53ae4ed9904df42e3f81c634['h0318a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c6] =  I0310077d53ae4ed9904df42e3f81c634['h0318c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c7] =  I0310077d53ae4ed9904df42e3f81c634['h0318e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c8] =  I0310077d53ae4ed9904df42e3f81c634['h03190] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018c9] =  I0310077d53ae4ed9904df42e3f81c634['h03192] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ca] =  I0310077d53ae4ed9904df42e3f81c634['h03194] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018cb] =  I0310077d53ae4ed9904df42e3f81c634['h03196] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018cc] =  I0310077d53ae4ed9904df42e3f81c634['h03198] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018cd] =  I0310077d53ae4ed9904df42e3f81c634['h0319a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ce] =  I0310077d53ae4ed9904df42e3f81c634['h0319c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018cf] =  I0310077d53ae4ed9904df42e3f81c634['h0319e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d0] =  I0310077d53ae4ed9904df42e3f81c634['h031a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d1] =  I0310077d53ae4ed9904df42e3f81c634['h031a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d2] =  I0310077d53ae4ed9904df42e3f81c634['h031a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d3] =  I0310077d53ae4ed9904df42e3f81c634['h031a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d4] =  I0310077d53ae4ed9904df42e3f81c634['h031a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d5] =  I0310077d53ae4ed9904df42e3f81c634['h031aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d6] =  I0310077d53ae4ed9904df42e3f81c634['h031ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d7] =  I0310077d53ae4ed9904df42e3f81c634['h031ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d8] =  I0310077d53ae4ed9904df42e3f81c634['h031b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018d9] =  I0310077d53ae4ed9904df42e3f81c634['h031b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018da] =  I0310077d53ae4ed9904df42e3f81c634['h031b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018db] =  I0310077d53ae4ed9904df42e3f81c634['h031b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018dc] =  I0310077d53ae4ed9904df42e3f81c634['h031b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018dd] =  I0310077d53ae4ed9904df42e3f81c634['h031ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018de] =  I0310077d53ae4ed9904df42e3f81c634['h031bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018df] =  I0310077d53ae4ed9904df42e3f81c634['h031be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e0] =  I0310077d53ae4ed9904df42e3f81c634['h031c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e1] =  I0310077d53ae4ed9904df42e3f81c634['h031c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e2] =  I0310077d53ae4ed9904df42e3f81c634['h031c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e3] =  I0310077d53ae4ed9904df42e3f81c634['h031c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e4] =  I0310077d53ae4ed9904df42e3f81c634['h031c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e5] =  I0310077d53ae4ed9904df42e3f81c634['h031ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e6] =  I0310077d53ae4ed9904df42e3f81c634['h031cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e7] =  I0310077d53ae4ed9904df42e3f81c634['h031ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e8] =  I0310077d53ae4ed9904df42e3f81c634['h031d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018e9] =  I0310077d53ae4ed9904df42e3f81c634['h031d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ea] =  I0310077d53ae4ed9904df42e3f81c634['h031d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018eb] =  I0310077d53ae4ed9904df42e3f81c634['h031d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ec] =  I0310077d53ae4ed9904df42e3f81c634['h031d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ed] =  I0310077d53ae4ed9904df42e3f81c634['h031da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ee] =  I0310077d53ae4ed9904df42e3f81c634['h031dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ef] =  I0310077d53ae4ed9904df42e3f81c634['h031de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f0] =  I0310077d53ae4ed9904df42e3f81c634['h031e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f1] =  I0310077d53ae4ed9904df42e3f81c634['h031e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f2] =  I0310077d53ae4ed9904df42e3f81c634['h031e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f3] =  I0310077d53ae4ed9904df42e3f81c634['h031e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f4] =  I0310077d53ae4ed9904df42e3f81c634['h031e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f5] =  I0310077d53ae4ed9904df42e3f81c634['h031ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f6] =  I0310077d53ae4ed9904df42e3f81c634['h031ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f7] =  I0310077d53ae4ed9904df42e3f81c634['h031ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f8] =  I0310077d53ae4ed9904df42e3f81c634['h031f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018f9] =  I0310077d53ae4ed9904df42e3f81c634['h031f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018fa] =  I0310077d53ae4ed9904df42e3f81c634['h031f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018fb] =  I0310077d53ae4ed9904df42e3f81c634['h031f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018fc] =  I0310077d53ae4ed9904df42e3f81c634['h031f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018fd] =  I0310077d53ae4ed9904df42e3f81c634['h031fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018fe] =  I0310077d53ae4ed9904df42e3f81c634['h031fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h018ff] =  I0310077d53ae4ed9904df42e3f81c634['h031fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01900] =  I0310077d53ae4ed9904df42e3f81c634['h03200] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01901] =  I0310077d53ae4ed9904df42e3f81c634['h03202] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01902] =  I0310077d53ae4ed9904df42e3f81c634['h03204] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01903] =  I0310077d53ae4ed9904df42e3f81c634['h03206] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01904] =  I0310077d53ae4ed9904df42e3f81c634['h03208] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01905] =  I0310077d53ae4ed9904df42e3f81c634['h0320a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01906] =  I0310077d53ae4ed9904df42e3f81c634['h0320c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01907] =  I0310077d53ae4ed9904df42e3f81c634['h0320e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01908] =  I0310077d53ae4ed9904df42e3f81c634['h03210] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01909] =  I0310077d53ae4ed9904df42e3f81c634['h03212] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0190a] =  I0310077d53ae4ed9904df42e3f81c634['h03214] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0190b] =  I0310077d53ae4ed9904df42e3f81c634['h03216] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0190c] =  I0310077d53ae4ed9904df42e3f81c634['h03218] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0190d] =  I0310077d53ae4ed9904df42e3f81c634['h0321a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0190e] =  I0310077d53ae4ed9904df42e3f81c634['h0321c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0190f] =  I0310077d53ae4ed9904df42e3f81c634['h0321e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01910] =  I0310077d53ae4ed9904df42e3f81c634['h03220] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01911] =  I0310077d53ae4ed9904df42e3f81c634['h03222] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01912] =  I0310077d53ae4ed9904df42e3f81c634['h03224] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01913] =  I0310077d53ae4ed9904df42e3f81c634['h03226] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01914] =  I0310077d53ae4ed9904df42e3f81c634['h03228] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01915] =  I0310077d53ae4ed9904df42e3f81c634['h0322a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01916] =  I0310077d53ae4ed9904df42e3f81c634['h0322c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01917] =  I0310077d53ae4ed9904df42e3f81c634['h0322e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01918] =  I0310077d53ae4ed9904df42e3f81c634['h03230] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01919] =  I0310077d53ae4ed9904df42e3f81c634['h03232] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0191a] =  I0310077d53ae4ed9904df42e3f81c634['h03234] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0191b] =  I0310077d53ae4ed9904df42e3f81c634['h03236] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0191c] =  I0310077d53ae4ed9904df42e3f81c634['h03238] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0191d] =  I0310077d53ae4ed9904df42e3f81c634['h0323a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0191e] =  I0310077d53ae4ed9904df42e3f81c634['h0323c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0191f] =  I0310077d53ae4ed9904df42e3f81c634['h0323e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01920] =  I0310077d53ae4ed9904df42e3f81c634['h03240] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01921] =  I0310077d53ae4ed9904df42e3f81c634['h03242] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01922] =  I0310077d53ae4ed9904df42e3f81c634['h03244] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01923] =  I0310077d53ae4ed9904df42e3f81c634['h03246] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01924] =  I0310077d53ae4ed9904df42e3f81c634['h03248] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01925] =  I0310077d53ae4ed9904df42e3f81c634['h0324a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01926] =  I0310077d53ae4ed9904df42e3f81c634['h0324c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01927] =  I0310077d53ae4ed9904df42e3f81c634['h0324e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01928] =  I0310077d53ae4ed9904df42e3f81c634['h03250] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01929] =  I0310077d53ae4ed9904df42e3f81c634['h03252] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0192a] =  I0310077d53ae4ed9904df42e3f81c634['h03254] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0192b] =  I0310077d53ae4ed9904df42e3f81c634['h03256] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0192c] =  I0310077d53ae4ed9904df42e3f81c634['h03258] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0192d] =  I0310077d53ae4ed9904df42e3f81c634['h0325a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0192e] =  I0310077d53ae4ed9904df42e3f81c634['h0325c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0192f] =  I0310077d53ae4ed9904df42e3f81c634['h0325e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01930] =  I0310077d53ae4ed9904df42e3f81c634['h03260] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01931] =  I0310077d53ae4ed9904df42e3f81c634['h03262] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01932] =  I0310077d53ae4ed9904df42e3f81c634['h03264] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01933] =  I0310077d53ae4ed9904df42e3f81c634['h03266] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01934] =  I0310077d53ae4ed9904df42e3f81c634['h03268] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01935] =  I0310077d53ae4ed9904df42e3f81c634['h0326a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01936] =  I0310077d53ae4ed9904df42e3f81c634['h0326c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01937] =  I0310077d53ae4ed9904df42e3f81c634['h0326e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01938] =  I0310077d53ae4ed9904df42e3f81c634['h03270] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01939] =  I0310077d53ae4ed9904df42e3f81c634['h03272] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0193a] =  I0310077d53ae4ed9904df42e3f81c634['h03274] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0193b] =  I0310077d53ae4ed9904df42e3f81c634['h03276] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0193c] =  I0310077d53ae4ed9904df42e3f81c634['h03278] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0193d] =  I0310077d53ae4ed9904df42e3f81c634['h0327a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0193e] =  I0310077d53ae4ed9904df42e3f81c634['h0327c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0193f] =  I0310077d53ae4ed9904df42e3f81c634['h0327e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01940] =  I0310077d53ae4ed9904df42e3f81c634['h03280] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01941] =  I0310077d53ae4ed9904df42e3f81c634['h03282] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01942] =  I0310077d53ae4ed9904df42e3f81c634['h03284] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01943] =  I0310077d53ae4ed9904df42e3f81c634['h03286] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01944] =  I0310077d53ae4ed9904df42e3f81c634['h03288] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01945] =  I0310077d53ae4ed9904df42e3f81c634['h0328a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01946] =  I0310077d53ae4ed9904df42e3f81c634['h0328c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01947] =  I0310077d53ae4ed9904df42e3f81c634['h0328e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01948] =  I0310077d53ae4ed9904df42e3f81c634['h03290] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01949] =  I0310077d53ae4ed9904df42e3f81c634['h03292] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0194a] =  I0310077d53ae4ed9904df42e3f81c634['h03294] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0194b] =  I0310077d53ae4ed9904df42e3f81c634['h03296] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0194c] =  I0310077d53ae4ed9904df42e3f81c634['h03298] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0194d] =  I0310077d53ae4ed9904df42e3f81c634['h0329a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0194e] =  I0310077d53ae4ed9904df42e3f81c634['h0329c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0194f] =  I0310077d53ae4ed9904df42e3f81c634['h0329e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01950] =  I0310077d53ae4ed9904df42e3f81c634['h032a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01951] =  I0310077d53ae4ed9904df42e3f81c634['h032a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01952] =  I0310077d53ae4ed9904df42e3f81c634['h032a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01953] =  I0310077d53ae4ed9904df42e3f81c634['h032a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01954] =  I0310077d53ae4ed9904df42e3f81c634['h032a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01955] =  I0310077d53ae4ed9904df42e3f81c634['h032aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01956] =  I0310077d53ae4ed9904df42e3f81c634['h032ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01957] =  I0310077d53ae4ed9904df42e3f81c634['h032ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01958] =  I0310077d53ae4ed9904df42e3f81c634['h032b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01959] =  I0310077d53ae4ed9904df42e3f81c634['h032b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0195a] =  I0310077d53ae4ed9904df42e3f81c634['h032b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0195b] =  I0310077d53ae4ed9904df42e3f81c634['h032b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0195c] =  I0310077d53ae4ed9904df42e3f81c634['h032b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0195d] =  I0310077d53ae4ed9904df42e3f81c634['h032ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0195e] =  I0310077d53ae4ed9904df42e3f81c634['h032bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0195f] =  I0310077d53ae4ed9904df42e3f81c634['h032be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01960] =  I0310077d53ae4ed9904df42e3f81c634['h032c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01961] =  I0310077d53ae4ed9904df42e3f81c634['h032c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01962] =  I0310077d53ae4ed9904df42e3f81c634['h032c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01963] =  I0310077d53ae4ed9904df42e3f81c634['h032c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01964] =  I0310077d53ae4ed9904df42e3f81c634['h032c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01965] =  I0310077d53ae4ed9904df42e3f81c634['h032ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01966] =  I0310077d53ae4ed9904df42e3f81c634['h032cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01967] =  I0310077d53ae4ed9904df42e3f81c634['h032ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01968] =  I0310077d53ae4ed9904df42e3f81c634['h032d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01969] =  I0310077d53ae4ed9904df42e3f81c634['h032d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0196a] =  I0310077d53ae4ed9904df42e3f81c634['h032d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0196b] =  I0310077d53ae4ed9904df42e3f81c634['h032d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0196c] =  I0310077d53ae4ed9904df42e3f81c634['h032d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0196d] =  I0310077d53ae4ed9904df42e3f81c634['h032da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0196e] =  I0310077d53ae4ed9904df42e3f81c634['h032dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0196f] =  I0310077d53ae4ed9904df42e3f81c634['h032de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01970] =  I0310077d53ae4ed9904df42e3f81c634['h032e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01971] =  I0310077d53ae4ed9904df42e3f81c634['h032e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01972] =  I0310077d53ae4ed9904df42e3f81c634['h032e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01973] =  I0310077d53ae4ed9904df42e3f81c634['h032e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01974] =  I0310077d53ae4ed9904df42e3f81c634['h032e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01975] =  I0310077d53ae4ed9904df42e3f81c634['h032ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01976] =  I0310077d53ae4ed9904df42e3f81c634['h032ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01977] =  I0310077d53ae4ed9904df42e3f81c634['h032ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01978] =  I0310077d53ae4ed9904df42e3f81c634['h032f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01979] =  I0310077d53ae4ed9904df42e3f81c634['h032f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0197a] =  I0310077d53ae4ed9904df42e3f81c634['h032f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0197b] =  I0310077d53ae4ed9904df42e3f81c634['h032f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0197c] =  I0310077d53ae4ed9904df42e3f81c634['h032f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0197d] =  I0310077d53ae4ed9904df42e3f81c634['h032fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0197e] =  I0310077d53ae4ed9904df42e3f81c634['h032fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0197f] =  I0310077d53ae4ed9904df42e3f81c634['h032fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01980] =  I0310077d53ae4ed9904df42e3f81c634['h03300] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01981] =  I0310077d53ae4ed9904df42e3f81c634['h03302] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01982] =  I0310077d53ae4ed9904df42e3f81c634['h03304] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01983] =  I0310077d53ae4ed9904df42e3f81c634['h03306] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01984] =  I0310077d53ae4ed9904df42e3f81c634['h03308] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01985] =  I0310077d53ae4ed9904df42e3f81c634['h0330a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01986] =  I0310077d53ae4ed9904df42e3f81c634['h0330c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01987] =  I0310077d53ae4ed9904df42e3f81c634['h0330e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01988] =  I0310077d53ae4ed9904df42e3f81c634['h03310] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01989] =  I0310077d53ae4ed9904df42e3f81c634['h03312] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0198a] =  I0310077d53ae4ed9904df42e3f81c634['h03314] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0198b] =  I0310077d53ae4ed9904df42e3f81c634['h03316] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0198c] =  I0310077d53ae4ed9904df42e3f81c634['h03318] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0198d] =  I0310077d53ae4ed9904df42e3f81c634['h0331a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0198e] =  I0310077d53ae4ed9904df42e3f81c634['h0331c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0198f] =  I0310077d53ae4ed9904df42e3f81c634['h0331e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01990] =  I0310077d53ae4ed9904df42e3f81c634['h03320] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01991] =  I0310077d53ae4ed9904df42e3f81c634['h03322] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01992] =  I0310077d53ae4ed9904df42e3f81c634['h03324] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01993] =  I0310077d53ae4ed9904df42e3f81c634['h03326] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01994] =  I0310077d53ae4ed9904df42e3f81c634['h03328] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01995] =  I0310077d53ae4ed9904df42e3f81c634['h0332a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01996] =  I0310077d53ae4ed9904df42e3f81c634['h0332c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01997] =  I0310077d53ae4ed9904df42e3f81c634['h0332e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01998] =  I0310077d53ae4ed9904df42e3f81c634['h03330] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01999] =  I0310077d53ae4ed9904df42e3f81c634['h03332] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0199a] =  I0310077d53ae4ed9904df42e3f81c634['h03334] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0199b] =  I0310077d53ae4ed9904df42e3f81c634['h03336] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0199c] =  I0310077d53ae4ed9904df42e3f81c634['h03338] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0199d] =  I0310077d53ae4ed9904df42e3f81c634['h0333a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0199e] =  I0310077d53ae4ed9904df42e3f81c634['h0333c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h0199f] =  I0310077d53ae4ed9904df42e3f81c634['h0333e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a0] =  I0310077d53ae4ed9904df42e3f81c634['h03340] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a1] =  I0310077d53ae4ed9904df42e3f81c634['h03342] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a2] =  I0310077d53ae4ed9904df42e3f81c634['h03344] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a3] =  I0310077d53ae4ed9904df42e3f81c634['h03346] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a4] =  I0310077d53ae4ed9904df42e3f81c634['h03348] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a5] =  I0310077d53ae4ed9904df42e3f81c634['h0334a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a6] =  I0310077d53ae4ed9904df42e3f81c634['h0334c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a7] =  I0310077d53ae4ed9904df42e3f81c634['h0334e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a8] =  I0310077d53ae4ed9904df42e3f81c634['h03350] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019a9] =  I0310077d53ae4ed9904df42e3f81c634['h03352] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019aa] =  I0310077d53ae4ed9904df42e3f81c634['h03354] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ab] =  I0310077d53ae4ed9904df42e3f81c634['h03356] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ac] =  I0310077d53ae4ed9904df42e3f81c634['h03358] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ad] =  I0310077d53ae4ed9904df42e3f81c634['h0335a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ae] =  I0310077d53ae4ed9904df42e3f81c634['h0335c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019af] =  I0310077d53ae4ed9904df42e3f81c634['h0335e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b0] =  I0310077d53ae4ed9904df42e3f81c634['h03360] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b1] =  I0310077d53ae4ed9904df42e3f81c634['h03362] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b2] =  I0310077d53ae4ed9904df42e3f81c634['h03364] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b3] =  I0310077d53ae4ed9904df42e3f81c634['h03366] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b4] =  I0310077d53ae4ed9904df42e3f81c634['h03368] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b5] =  I0310077d53ae4ed9904df42e3f81c634['h0336a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b6] =  I0310077d53ae4ed9904df42e3f81c634['h0336c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b7] =  I0310077d53ae4ed9904df42e3f81c634['h0336e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b8] =  I0310077d53ae4ed9904df42e3f81c634['h03370] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019b9] =  I0310077d53ae4ed9904df42e3f81c634['h03372] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ba] =  I0310077d53ae4ed9904df42e3f81c634['h03374] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019bb] =  I0310077d53ae4ed9904df42e3f81c634['h03376] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019bc] =  I0310077d53ae4ed9904df42e3f81c634['h03378] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019bd] =  I0310077d53ae4ed9904df42e3f81c634['h0337a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019be] =  I0310077d53ae4ed9904df42e3f81c634['h0337c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019bf] =  I0310077d53ae4ed9904df42e3f81c634['h0337e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c0] =  I0310077d53ae4ed9904df42e3f81c634['h03380] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c1] =  I0310077d53ae4ed9904df42e3f81c634['h03382] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c2] =  I0310077d53ae4ed9904df42e3f81c634['h03384] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c3] =  I0310077d53ae4ed9904df42e3f81c634['h03386] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c4] =  I0310077d53ae4ed9904df42e3f81c634['h03388] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c5] =  I0310077d53ae4ed9904df42e3f81c634['h0338a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c6] =  I0310077d53ae4ed9904df42e3f81c634['h0338c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c7] =  I0310077d53ae4ed9904df42e3f81c634['h0338e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c8] =  I0310077d53ae4ed9904df42e3f81c634['h03390] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019c9] =  I0310077d53ae4ed9904df42e3f81c634['h03392] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ca] =  I0310077d53ae4ed9904df42e3f81c634['h03394] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019cb] =  I0310077d53ae4ed9904df42e3f81c634['h03396] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019cc] =  I0310077d53ae4ed9904df42e3f81c634['h03398] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019cd] =  I0310077d53ae4ed9904df42e3f81c634['h0339a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ce] =  I0310077d53ae4ed9904df42e3f81c634['h0339c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019cf] =  I0310077d53ae4ed9904df42e3f81c634['h0339e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d0] =  I0310077d53ae4ed9904df42e3f81c634['h033a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d1] =  I0310077d53ae4ed9904df42e3f81c634['h033a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d2] =  I0310077d53ae4ed9904df42e3f81c634['h033a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d3] =  I0310077d53ae4ed9904df42e3f81c634['h033a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d4] =  I0310077d53ae4ed9904df42e3f81c634['h033a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d5] =  I0310077d53ae4ed9904df42e3f81c634['h033aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d6] =  I0310077d53ae4ed9904df42e3f81c634['h033ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d7] =  I0310077d53ae4ed9904df42e3f81c634['h033ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d8] =  I0310077d53ae4ed9904df42e3f81c634['h033b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019d9] =  I0310077d53ae4ed9904df42e3f81c634['h033b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019da] =  I0310077d53ae4ed9904df42e3f81c634['h033b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019db] =  I0310077d53ae4ed9904df42e3f81c634['h033b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019dc] =  I0310077d53ae4ed9904df42e3f81c634['h033b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019dd] =  I0310077d53ae4ed9904df42e3f81c634['h033ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019de] =  I0310077d53ae4ed9904df42e3f81c634['h033bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019df] =  I0310077d53ae4ed9904df42e3f81c634['h033be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e0] =  I0310077d53ae4ed9904df42e3f81c634['h033c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e1] =  I0310077d53ae4ed9904df42e3f81c634['h033c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e2] =  I0310077d53ae4ed9904df42e3f81c634['h033c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e3] =  I0310077d53ae4ed9904df42e3f81c634['h033c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e4] =  I0310077d53ae4ed9904df42e3f81c634['h033c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e5] =  I0310077d53ae4ed9904df42e3f81c634['h033ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e6] =  I0310077d53ae4ed9904df42e3f81c634['h033cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e7] =  I0310077d53ae4ed9904df42e3f81c634['h033ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e8] =  I0310077d53ae4ed9904df42e3f81c634['h033d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019e9] =  I0310077d53ae4ed9904df42e3f81c634['h033d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ea] =  I0310077d53ae4ed9904df42e3f81c634['h033d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019eb] =  I0310077d53ae4ed9904df42e3f81c634['h033d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ec] =  I0310077d53ae4ed9904df42e3f81c634['h033d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ed] =  I0310077d53ae4ed9904df42e3f81c634['h033da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ee] =  I0310077d53ae4ed9904df42e3f81c634['h033dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ef] =  I0310077d53ae4ed9904df42e3f81c634['h033de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f0] =  I0310077d53ae4ed9904df42e3f81c634['h033e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f1] =  I0310077d53ae4ed9904df42e3f81c634['h033e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f2] =  I0310077d53ae4ed9904df42e3f81c634['h033e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f3] =  I0310077d53ae4ed9904df42e3f81c634['h033e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f4] =  I0310077d53ae4ed9904df42e3f81c634['h033e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f5] =  I0310077d53ae4ed9904df42e3f81c634['h033ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f6] =  I0310077d53ae4ed9904df42e3f81c634['h033ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f7] =  I0310077d53ae4ed9904df42e3f81c634['h033ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f8] =  I0310077d53ae4ed9904df42e3f81c634['h033f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019f9] =  I0310077d53ae4ed9904df42e3f81c634['h033f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019fa] =  I0310077d53ae4ed9904df42e3f81c634['h033f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019fb] =  I0310077d53ae4ed9904df42e3f81c634['h033f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019fc] =  I0310077d53ae4ed9904df42e3f81c634['h033f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019fd] =  I0310077d53ae4ed9904df42e3f81c634['h033fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019fe] =  I0310077d53ae4ed9904df42e3f81c634['h033fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h019ff] =  I0310077d53ae4ed9904df42e3f81c634['h033fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a00] =  I0310077d53ae4ed9904df42e3f81c634['h03400] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a01] =  I0310077d53ae4ed9904df42e3f81c634['h03402] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a02] =  I0310077d53ae4ed9904df42e3f81c634['h03404] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a03] =  I0310077d53ae4ed9904df42e3f81c634['h03406] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a04] =  I0310077d53ae4ed9904df42e3f81c634['h03408] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a05] =  I0310077d53ae4ed9904df42e3f81c634['h0340a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a06] =  I0310077d53ae4ed9904df42e3f81c634['h0340c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a07] =  I0310077d53ae4ed9904df42e3f81c634['h0340e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a08] =  I0310077d53ae4ed9904df42e3f81c634['h03410] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a09] =  I0310077d53ae4ed9904df42e3f81c634['h03412] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a0a] =  I0310077d53ae4ed9904df42e3f81c634['h03414] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a0b] =  I0310077d53ae4ed9904df42e3f81c634['h03416] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a0c] =  I0310077d53ae4ed9904df42e3f81c634['h03418] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a0d] =  I0310077d53ae4ed9904df42e3f81c634['h0341a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a0e] =  I0310077d53ae4ed9904df42e3f81c634['h0341c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a0f] =  I0310077d53ae4ed9904df42e3f81c634['h0341e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a10] =  I0310077d53ae4ed9904df42e3f81c634['h03420] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a11] =  I0310077d53ae4ed9904df42e3f81c634['h03422] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a12] =  I0310077d53ae4ed9904df42e3f81c634['h03424] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a13] =  I0310077d53ae4ed9904df42e3f81c634['h03426] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a14] =  I0310077d53ae4ed9904df42e3f81c634['h03428] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a15] =  I0310077d53ae4ed9904df42e3f81c634['h0342a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a16] =  I0310077d53ae4ed9904df42e3f81c634['h0342c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a17] =  I0310077d53ae4ed9904df42e3f81c634['h0342e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a18] =  I0310077d53ae4ed9904df42e3f81c634['h03430] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a19] =  I0310077d53ae4ed9904df42e3f81c634['h03432] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a1a] =  I0310077d53ae4ed9904df42e3f81c634['h03434] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a1b] =  I0310077d53ae4ed9904df42e3f81c634['h03436] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a1c] =  I0310077d53ae4ed9904df42e3f81c634['h03438] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a1d] =  I0310077d53ae4ed9904df42e3f81c634['h0343a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a1e] =  I0310077d53ae4ed9904df42e3f81c634['h0343c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a1f] =  I0310077d53ae4ed9904df42e3f81c634['h0343e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a20] =  I0310077d53ae4ed9904df42e3f81c634['h03440] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a21] =  I0310077d53ae4ed9904df42e3f81c634['h03442] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a22] =  I0310077d53ae4ed9904df42e3f81c634['h03444] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a23] =  I0310077d53ae4ed9904df42e3f81c634['h03446] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a24] =  I0310077d53ae4ed9904df42e3f81c634['h03448] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a25] =  I0310077d53ae4ed9904df42e3f81c634['h0344a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a26] =  I0310077d53ae4ed9904df42e3f81c634['h0344c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a27] =  I0310077d53ae4ed9904df42e3f81c634['h0344e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a28] =  I0310077d53ae4ed9904df42e3f81c634['h03450] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a29] =  I0310077d53ae4ed9904df42e3f81c634['h03452] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a2a] =  I0310077d53ae4ed9904df42e3f81c634['h03454] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a2b] =  I0310077d53ae4ed9904df42e3f81c634['h03456] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a2c] =  I0310077d53ae4ed9904df42e3f81c634['h03458] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a2d] =  I0310077d53ae4ed9904df42e3f81c634['h0345a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a2e] =  I0310077d53ae4ed9904df42e3f81c634['h0345c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a2f] =  I0310077d53ae4ed9904df42e3f81c634['h0345e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a30] =  I0310077d53ae4ed9904df42e3f81c634['h03460] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a31] =  I0310077d53ae4ed9904df42e3f81c634['h03462] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a32] =  I0310077d53ae4ed9904df42e3f81c634['h03464] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a33] =  I0310077d53ae4ed9904df42e3f81c634['h03466] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a34] =  I0310077d53ae4ed9904df42e3f81c634['h03468] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a35] =  I0310077d53ae4ed9904df42e3f81c634['h0346a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a36] =  I0310077d53ae4ed9904df42e3f81c634['h0346c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a37] =  I0310077d53ae4ed9904df42e3f81c634['h0346e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a38] =  I0310077d53ae4ed9904df42e3f81c634['h03470] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a39] =  I0310077d53ae4ed9904df42e3f81c634['h03472] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a3a] =  I0310077d53ae4ed9904df42e3f81c634['h03474] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a3b] =  I0310077d53ae4ed9904df42e3f81c634['h03476] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a3c] =  I0310077d53ae4ed9904df42e3f81c634['h03478] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a3d] =  I0310077d53ae4ed9904df42e3f81c634['h0347a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a3e] =  I0310077d53ae4ed9904df42e3f81c634['h0347c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a3f] =  I0310077d53ae4ed9904df42e3f81c634['h0347e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a40] =  I0310077d53ae4ed9904df42e3f81c634['h03480] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a41] =  I0310077d53ae4ed9904df42e3f81c634['h03482] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a42] =  I0310077d53ae4ed9904df42e3f81c634['h03484] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a43] =  I0310077d53ae4ed9904df42e3f81c634['h03486] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a44] =  I0310077d53ae4ed9904df42e3f81c634['h03488] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a45] =  I0310077d53ae4ed9904df42e3f81c634['h0348a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a46] =  I0310077d53ae4ed9904df42e3f81c634['h0348c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a47] =  I0310077d53ae4ed9904df42e3f81c634['h0348e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a48] =  I0310077d53ae4ed9904df42e3f81c634['h03490] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a49] =  I0310077d53ae4ed9904df42e3f81c634['h03492] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a4a] =  I0310077d53ae4ed9904df42e3f81c634['h03494] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a4b] =  I0310077d53ae4ed9904df42e3f81c634['h03496] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a4c] =  I0310077d53ae4ed9904df42e3f81c634['h03498] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a4d] =  I0310077d53ae4ed9904df42e3f81c634['h0349a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a4e] =  I0310077d53ae4ed9904df42e3f81c634['h0349c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a4f] =  I0310077d53ae4ed9904df42e3f81c634['h0349e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a50] =  I0310077d53ae4ed9904df42e3f81c634['h034a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a51] =  I0310077d53ae4ed9904df42e3f81c634['h034a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a52] =  I0310077d53ae4ed9904df42e3f81c634['h034a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a53] =  I0310077d53ae4ed9904df42e3f81c634['h034a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a54] =  I0310077d53ae4ed9904df42e3f81c634['h034a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a55] =  I0310077d53ae4ed9904df42e3f81c634['h034aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a56] =  I0310077d53ae4ed9904df42e3f81c634['h034ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a57] =  I0310077d53ae4ed9904df42e3f81c634['h034ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a58] =  I0310077d53ae4ed9904df42e3f81c634['h034b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a59] =  I0310077d53ae4ed9904df42e3f81c634['h034b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a5a] =  I0310077d53ae4ed9904df42e3f81c634['h034b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a5b] =  I0310077d53ae4ed9904df42e3f81c634['h034b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a5c] =  I0310077d53ae4ed9904df42e3f81c634['h034b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a5d] =  I0310077d53ae4ed9904df42e3f81c634['h034ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a5e] =  I0310077d53ae4ed9904df42e3f81c634['h034bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a5f] =  I0310077d53ae4ed9904df42e3f81c634['h034be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a60] =  I0310077d53ae4ed9904df42e3f81c634['h034c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a61] =  I0310077d53ae4ed9904df42e3f81c634['h034c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a62] =  I0310077d53ae4ed9904df42e3f81c634['h034c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a63] =  I0310077d53ae4ed9904df42e3f81c634['h034c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a64] =  I0310077d53ae4ed9904df42e3f81c634['h034c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a65] =  I0310077d53ae4ed9904df42e3f81c634['h034ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a66] =  I0310077d53ae4ed9904df42e3f81c634['h034cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a67] =  I0310077d53ae4ed9904df42e3f81c634['h034ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a68] =  I0310077d53ae4ed9904df42e3f81c634['h034d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a69] =  I0310077d53ae4ed9904df42e3f81c634['h034d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a6a] =  I0310077d53ae4ed9904df42e3f81c634['h034d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a6b] =  I0310077d53ae4ed9904df42e3f81c634['h034d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a6c] =  I0310077d53ae4ed9904df42e3f81c634['h034d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a6d] =  I0310077d53ae4ed9904df42e3f81c634['h034da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a6e] =  I0310077d53ae4ed9904df42e3f81c634['h034dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a6f] =  I0310077d53ae4ed9904df42e3f81c634['h034de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a70] =  I0310077d53ae4ed9904df42e3f81c634['h034e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a71] =  I0310077d53ae4ed9904df42e3f81c634['h034e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a72] =  I0310077d53ae4ed9904df42e3f81c634['h034e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a73] =  I0310077d53ae4ed9904df42e3f81c634['h034e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a74] =  I0310077d53ae4ed9904df42e3f81c634['h034e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a75] =  I0310077d53ae4ed9904df42e3f81c634['h034ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a76] =  I0310077d53ae4ed9904df42e3f81c634['h034ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a77] =  I0310077d53ae4ed9904df42e3f81c634['h034ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a78] =  I0310077d53ae4ed9904df42e3f81c634['h034f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a79] =  I0310077d53ae4ed9904df42e3f81c634['h034f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a7a] =  I0310077d53ae4ed9904df42e3f81c634['h034f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a7b] =  I0310077d53ae4ed9904df42e3f81c634['h034f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a7c] =  I0310077d53ae4ed9904df42e3f81c634['h034f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a7d] =  I0310077d53ae4ed9904df42e3f81c634['h034fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a7e] =  I0310077d53ae4ed9904df42e3f81c634['h034fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a7f] =  I0310077d53ae4ed9904df42e3f81c634['h034fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a80] =  I0310077d53ae4ed9904df42e3f81c634['h03500] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a81] =  I0310077d53ae4ed9904df42e3f81c634['h03502] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a82] =  I0310077d53ae4ed9904df42e3f81c634['h03504] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a83] =  I0310077d53ae4ed9904df42e3f81c634['h03506] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a84] =  I0310077d53ae4ed9904df42e3f81c634['h03508] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a85] =  I0310077d53ae4ed9904df42e3f81c634['h0350a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a86] =  I0310077d53ae4ed9904df42e3f81c634['h0350c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a87] =  I0310077d53ae4ed9904df42e3f81c634['h0350e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a88] =  I0310077d53ae4ed9904df42e3f81c634['h03510] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a89] =  I0310077d53ae4ed9904df42e3f81c634['h03512] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a8a] =  I0310077d53ae4ed9904df42e3f81c634['h03514] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a8b] =  I0310077d53ae4ed9904df42e3f81c634['h03516] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a8c] =  I0310077d53ae4ed9904df42e3f81c634['h03518] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a8d] =  I0310077d53ae4ed9904df42e3f81c634['h0351a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a8e] =  I0310077d53ae4ed9904df42e3f81c634['h0351c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a8f] =  I0310077d53ae4ed9904df42e3f81c634['h0351e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a90] =  I0310077d53ae4ed9904df42e3f81c634['h03520] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a91] =  I0310077d53ae4ed9904df42e3f81c634['h03522] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a92] =  I0310077d53ae4ed9904df42e3f81c634['h03524] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a93] =  I0310077d53ae4ed9904df42e3f81c634['h03526] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a94] =  I0310077d53ae4ed9904df42e3f81c634['h03528] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a95] =  I0310077d53ae4ed9904df42e3f81c634['h0352a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a96] =  I0310077d53ae4ed9904df42e3f81c634['h0352c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a97] =  I0310077d53ae4ed9904df42e3f81c634['h0352e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a98] =  I0310077d53ae4ed9904df42e3f81c634['h03530] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a99] =  I0310077d53ae4ed9904df42e3f81c634['h03532] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a9a] =  I0310077d53ae4ed9904df42e3f81c634['h03534] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a9b] =  I0310077d53ae4ed9904df42e3f81c634['h03536] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a9c] =  I0310077d53ae4ed9904df42e3f81c634['h03538] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a9d] =  I0310077d53ae4ed9904df42e3f81c634['h0353a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a9e] =  I0310077d53ae4ed9904df42e3f81c634['h0353c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01a9f] =  I0310077d53ae4ed9904df42e3f81c634['h0353e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa0] =  I0310077d53ae4ed9904df42e3f81c634['h03540] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa1] =  I0310077d53ae4ed9904df42e3f81c634['h03542] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa2] =  I0310077d53ae4ed9904df42e3f81c634['h03544] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa3] =  I0310077d53ae4ed9904df42e3f81c634['h03546] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa4] =  I0310077d53ae4ed9904df42e3f81c634['h03548] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa5] =  I0310077d53ae4ed9904df42e3f81c634['h0354a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa6] =  I0310077d53ae4ed9904df42e3f81c634['h0354c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa7] =  I0310077d53ae4ed9904df42e3f81c634['h0354e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa8] =  I0310077d53ae4ed9904df42e3f81c634['h03550] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aa9] =  I0310077d53ae4ed9904df42e3f81c634['h03552] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aaa] =  I0310077d53ae4ed9904df42e3f81c634['h03554] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aab] =  I0310077d53ae4ed9904df42e3f81c634['h03556] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aac] =  I0310077d53ae4ed9904df42e3f81c634['h03558] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aad] =  I0310077d53ae4ed9904df42e3f81c634['h0355a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aae] =  I0310077d53ae4ed9904df42e3f81c634['h0355c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aaf] =  I0310077d53ae4ed9904df42e3f81c634['h0355e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab0] =  I0310077d53ae4ed9904df42e3f81c634['h03560] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab1] =  I0310077d53ae4ed9904df42e3f81c634['h03562] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab2] =  I0310077d53ae4ed9904df42e3f81c634['h03564] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab3] =  I0310077d53ae4ed9904df42e3f81c634['h03566] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab4] =  I0310077d53ae4ed9904df42e3f81c634['h03568] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab5] =  I0310077d53ae4ed9904df42e3f81c634['h0356a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab6] =  I0310077d53ae4ed9904df42e3f81c634['h0356c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab7] =  I0310077d53ae4ed9904df42e3f81c634['h0356e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab8] =  I0310077d53ae4ed9904df42e3f81c634['h03570] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ab9] =  I0310077d53ae4ed9904df42e3f81c634['h03572] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aba] =  I0310077d53ae4ed9904df42e3f81c634['h03574] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01abb] =  I0310077d53ae4ed9904df42e3f81c634['h03576] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01abc] =  I0310077d53ae4ed9904df42e3f81c634['h03578] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01abd] =  I0310077d53ae4ed9904df42e3f81c634['h0357a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01abe] =  I0310077d53ae4ed9904df42e3f81c634['h0357c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01abf] =  I0310077d53ae4ed9904df42e3f81c634['h0357e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac0] =  I0310077d53ae4ed9904df42e3f81c634['h03580] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac1] =  I0310077d53ae4ed9904df42e3f81c634['h03582] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac2] =  I0310077d53ae4ed9904df42e3f81c634['h03584] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac3] =  I0310077d53ae4ed9904df42e3f81c634['h03586] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac4] =  I0310077d53ae4ed9904df42e3f81c634['h03588] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac5] =  I0310077d53ae4ed9904df42e3f81c634['h0358a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac6] =  I0310077d53ae4ed9904df42e3f81c634['h0358c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac7] =  I0310077d53ae4ed9904df42e3f81c634['h0358e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac8] =  I0310077d53ae4ed9904df42e3f81c634['h03590] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ac9] =  I0310077d53ae4ed9904df42e3f81c634['h03592] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aca] =  I0310077d53ae4ed9904df42e3f81c634['h03594] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01acb] =  I0310077d53ae4ed9904df42e3f81c634['h03596] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01acc] =  I0310077d53ae4ed9904df42e3f81c634['h03598] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01acd] =  I0310077d53ae4ed9904df42e3f81c634['h0359a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ace] =  I0310077d53ae4ed9904df42e3f81c634['h0359c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01acf] =  I0310077d53ae4ed9904df42e3f81c634['h0359e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad0] =  I0310077d53ae4ed9904df42e3f81c634['h035a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad1] =  I0310077d53ae4ed9904df42e3f81c634['h035a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad2] =  I0310077d53ae4ed9904df42e3f81c634['h035a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad3] =  I0310077d53ae4ed9904df42e3f81c634['h035a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad4] =  I0310077d53ae4ed9904df42e3f81c634['h035a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad5] =  I0310077d53ae4ed9904df42e3f81c634['h035aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad6] =  I0310077d53ae4ed9904df42e3f81c634['h035ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad7] =  I0310077d53ae4ed9904df42e3f81c634['h035ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad8] =  I0310077d53ae4ed9904df42e3f81c634['h035b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ad9] =  I0310077d53ae4ed9904df42e3f81c634['h035b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ada] =  I0310077d53ae4ed9904df42e3f81c634['h035b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01adb] =  I0310077d53ae4ed9904df42e3f81c634['h035b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01adc] =  I0310077d53ae4ed9904df42e3f81c634['h035b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01add] =  I0310077d53ae4ed9904df42e3f81c634['h035ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ade] =  I0310077d53ae4ed9904df42e3f81c634['h035bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01adf] =  I0310077d53ae4ed9904df42e3f81c634['h035be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae0] =  I0310077d53ae4ed9904df42e3f81c634['h035c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae1] =  I0310077d53ae4ed9904df42e3f81c634['h035c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae2] =  I0310077d53ae4ed9904df42e3f81c634['h035c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae3] =  I0310077d53ae4ed9904df42e3f81c634['h035c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae4] =  I0310077d53ae4ed9904df42e3f81c634['h035c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae5] =  I0310077d53ae4ed9904df42e3f81c634['h035ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae6] =  I0310077d53ae4ed9904df42e3f81c634['h035cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae7] =  I0310077d53ae4ed9904df42e3f81c634['h035ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae8] =  I0310077d53ae4ed9904df42e3f81c634['h035d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ae9] =  I0310077d53ae4ed9904df42e3f81c634['h035d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aea] =  I0310077d53ae4ed9904df42e3f81c634['h035d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aeb] =  I0310077d53ae4ed9904df42e3f81c634['h035d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aec] =  I0310077d53ae4ed9904df42e3f81c634['h035d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aed] =  I0310077d53ae4ed9904df42e3f81c634['h035da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aee] =  I0310077d53ae4ed9904df42e3f81c634['h035dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aef] =  I0310077d53ae4ed9904df42e3f81c634['h035de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af0] =  I0310077d53ae4ed9904df42e3f81c634['h035e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af1] =  I0310077d53ae4ed9904df42e3f81c634['h035e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af2] =  I0310077d53ae4ed9904df42e3f81c634['h035e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af3] =  I0310077d53ae4ed9904df42e3f81c634['h035e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af4] =  I0310077d53ae4ed9904df42e3f81c634['h035e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af5] =  I0310077d53ae4ed9904df42e3f81c634['h035ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af6] =  I0310077d53ae4ed9904df42e3f81c634['h035ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af7] =  I0310077d53ae4ed9904df42e3f81c634['h035ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af8] =  I0310077d53ae4ed9904df42e3f81c634['h035f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01af9] =  I0310077d53ae4ed9904df42e3f81c634['h035f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01afa] =  I0310077d53ae4ed9904df42e3f81c634['h035f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01afb] =  I0310077d53ae4ed9904df42e3f81c634['h035f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01afc] =  I0310077d53ae4ed9904df42e3f81c634['h035f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01afd] =  I0310077d53ae4ed9904df42e3f81c634['h035fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01afe] =  I0310077d53ae4ed9904df42e3f81c634['h035fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01aff] =  I0310077d53ae4ed9904df42e3f81c634['h035fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b00] =  I0310077d53ae4ed9904df42e3f81c634['h03600] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b01] =  I0310077d53ae4ed9904df42e3f81c634['h03602] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b02] =  I0310077d53ae4ed9904df42e3f81c634['h03604] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b03] =  I0310077d53ae4ed9904df42e3f81c634['h03606] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b04] =  I0310077d53ae4ed9904df42e3f81c634['h03608] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b05] =  I0310077d53ae4ed9904df42e3f81c634['h0360a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b06] =  I0310077d53ae4ed9904df42e3f81c634['h0360c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b07] =  I0310077d53ae4ed9904df42e3f81c634['h0360e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b08] =  I0310077d53ae4ed9904df42e3f81c634['h03610] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b09] =  I0310077d53ae4ed9904df42e3f81c634['h03612] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b0a] =  I0310077d53ae4ed9904df42e3f81c634['h03614] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b0b] =  I0310077d53ae4ed9904df42e3f81c634['h03616] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b0c] =  I0310077d53ae4ed9904df42e3f81c634['h03618] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b0d] =  I0310077d53ae4ed9904df42e3f81c634['h0361a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b0e] =  I0310077d53ae4ed9904df42e3f81c634['h0361c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b0f] =  I0310077d53ae4ed9904df42e3f81c634['h0361e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b10] =  I0310077d53ae4ed9904df42e3f81c634['h03620] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b11] =  I0310077d53ae4ed9904df42e3f81c634['h03622] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b12] =  I0310077d53ae4ed9904df42e3f81c634['h03624] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b13] =  I0310077d53ae4ed9904df42e3f81c634['h03626] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b14] =  I0310077d53ae4ed9904df42e3f81c634['h03628] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b15] =  I0310077d53ae4ed9904df42e3f81c634['h0362a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b16] =  I0310077d53ae4ed9904df42e3f81c634['h0362c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b17] =  I0310077d53ae4ed9904df42e3f81c634['h0362e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b18] =  I0310077d53ae4ed9904df42e3f81c634['h03630] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b19] =  I0310077d53ae4ed9904df42e3f81c634['h03632] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b1a] =  I0310077d53ae4ed9904df42e3f81c634['h03634] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b1b] =  I0310077d53ae4ed9904df42e3f81c634['h03636] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b1c] =  I0310077d53ae4ed9904df42e3f81c634['h03638] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b1d] =  I0310077d53ae4ed9904df42e3f81c634['h0363a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b1e] =  I0310077d53ae4ed9904df42e3f81c634['h0363c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b1f] =  I0310077d53ae4ed9904df42e3f81c634['h0363e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b20] =  I0310077d53ae4ed9904df42e3f81c634['h03640] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b21] =  I0310077d53ae4ed9904df42e3f81c634['h03642] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b22] =  I0310077d53ae4ed9904df42e3f81c634['h03644] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b23] =  I0310077d53ae4ed9904df42e3f81c634['h03646] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b24] =  I0310077d53ae4ed9904df42e3f81c634['h03648] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b25] =  I0310077d53ae4ed9904df42e3f81c634['h0364a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b26] =  I0310077d53ae4ed9904df42e3f81c634['h0364c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b27] =  I0310077d53ae4ed9904df42e3f81c634['h0364e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b28] =  I0310077d53ae4ed9904df42e3f81c634['h03650] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b29] =  I0310077d53ae4ed9904df42e3f81c634['h03652] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b2a] =  I0310077d53ae4ed9904df42e3f81c634['h03654] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b2b] =  I0310077d53ae4ed9904df42e3f81c634['h03656] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b2c] =  I0310077d53ae4ed9904df42e3f81c634['h03658] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b2d] =  I0310077d53ae4ed9904df42e3f81c634['h0365a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b2e] =  I0310077d53ae4ed9904df42e3f81c634['h0365c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b2f] =  I0310077d53ae4ed9904df42e3f81c634['h0365e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b30] =  I0310077d53ae4ed9904df42e3f81c634['h03660] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b31] =  I0310077d53ae4ed9904df42e3f81c634['h03662] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b32] =  I0310077d53ae4ed9904df42e3f81c634['h03664] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b33] =  I0310077d53ae4ed9904df42e3f81c634['h03666] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b34] =  I0310077d53ae4ed9904df42e3f81c634['h03668] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b35] =  I0310077d53ae4ed9904df42e3f81c634['h0366a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b36] =  I0310077d53ae4ed9904df42e3f81c634['h0366c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b37] =  I0310077d53ae4ed9904df42e3f81c634['h0366e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b38] =  I0310077d53ae4ed9904df42e3f81c634['h03670] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b39] =  I0310077d53ae4ed9904df42e3f81c634['h03672] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b3a] =  I0310077d53ae4ed9904df42e3f81c634['h03674] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b3b] =  I0310077d53ae4ed9904df42e3f81c634['h03676] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b3c] =  I0310077d53ae4ed9904df42e3f81c634['h03678] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b3d] =  I0310077d53ae4ed9904df42e3f81c634['h0367a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b3e] =  I0310077d53ae4ed9904df42e3f81c634['h0367c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b3f] =  I0310077d53ae4ed9904df42e3f81c634['h0367e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b40] =  I0310077d53ae4ed9904df42e3f81c634['h03680] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b41] =  I0310077d53ae4ed9904df42e3f81c634['h03682] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b42] =  I0310077d53ae4ed9904df42e3f81c634['h03684] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b43] =  I0310077d53ae4ed9904df42e3f81c634['h03686] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b44] =  I0310077d53ae4ed9904df42e3f81c634['h03688] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b45] =  I0310077d53ae4ed9904df42e3f81c634['h0368a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b46] =  I0310077d53ae4ed9904df42e3f81c634['h0368c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b47] =  I0310077d53ae4ed9904df42e3f81c634['h0368e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b48] =  I0310077d53ae4ed9904df42e3f81c634['h03690] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b49] =  I0310077d53ae4ed9904df42e3f81c634['h03692] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b4a] =  I0310077d53ae4ed9904df42e3f81c634['h03694] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b4b] =  I0310077d53ae4ed9904df42e3f81c634['h03696] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b4c] =  I0310077d53ae4ed9904df42e3f81c634['h03698] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b4d] =  I0310077d53ae4ed9904df42e3f81c634['h0369a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b4e] =  I0310077d53ae4ed9904df42e3f81c634['h0369c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b4f] =  I0310077d53ae4ed9904df42e3f81c634['h0369e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b50] =  I0310077d53ae4ed9904df42e3f81c634['h036a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b51] =  I0310077d53ae4ed9904df42e3f81c634['h036a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b52] =  I0310077d53ae4ed9904df42e3f81c634['h036a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b53] =  I0310077d53ae4ed9904df42e3f81c634['h036a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b54] =  I0310077d53ae4ed9904df42e3f81c634['h036a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b55] =  I0310077d53ae4ed9904df42e3f81c634['h036aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b56] =  I0310077d53ae4ed9904df42e3f81c634['h036ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b57] =  I0310077d53ae4ed9904df42e3f81c634['h036ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b58] =  I0310077d53ae4ed9904df42e3f81c634['h036b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b59] =  I0310077d53ae4ed9904df42e3f81c634['h036b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b5a] =  I0310077d53ae4ed9904df42e3f81c634['h036b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b5b] =  I0310077d53ae4ed9904df42e3f81c634['h036b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b5c] =  I0310077d53ae4ed9904df42e3f81c634['h036b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b5d] =  I0310077d53ae4ed9904df42e3f81c634['h036ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b5e] =  I0310077d53ae4ed9904df42e3f81c634['h036bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b5f] =  I0310077d53ae4ed9904df42e3f81c634['h036be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b60] =  I0310077d53ae4ed9904df42e3f81c634['h036c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b61] =  I0310077d53ae4ed9904df42e3f81c634['h036c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b62] =  I0310077d53ae4ed9904df42e3f81c634['h036c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b63] =  I0310077d53ae4ed9904df42e3f81c634['h036c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b64] =  I0310077d53ae4ed9904df42e3f81c634['h036c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b65] =  I0310077d53ae4ed9904df42e3f81c634['h036ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b66] =  I0310077d53ae4ed9904df42e3f81c634['h036cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b67] =  I0310077d53ae4ed9904df42e3f81c634['h036ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b68] =  I0310077d53ae4ed9904df42e3f81c634['h036d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b69] =  I0310077d53ae4ed9904df42e3f81c634['h036d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b6a] =  I0310077d53ae4ed9904df42e3f81c634['h036d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b6b] =  I0310077d53ae4ed9904df42e3f81c634['h036d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b6c] =  I0310077d53ae4ed9904df42e3f81c634['h036d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b6d] =  I0310077d53ae4ed9904df42e3f81c634['h036da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b6e] =  I0310077d53ae4ed9904df42e3f81c634['h036dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b6f] =  I0310077d53ae4ed9904df42e3f81c634['h036de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b70] =  I0310077d53ae4ed9904df42e3f81c634['h036e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b71] =  I0310077d53ae4ed9904df42e3f81c634['h036e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b72] =  I0310077d53ae4ed9904df42e3f81c634['h036e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b73] =  I0310077d53ae4ed9904df42e3f81c634['h036e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b74] =  I0310077d53ae4ed9904df42e3f81c634['h036e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b75] =  I0310077d53ae4ed9904df42e3f81c634['h036ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b76] =  I0310077d53ae4ed9904df42e3f81c634['h036ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b77] =  I0310077d53ae4ed9904df42e3f81c634['h036ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b78] =  I0310077d53ae4ed9904df42e3f81c634['h036f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b79] =  I0310077d53ae4ed9904df42e3f81c634['h036f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b7a] =  I0310077d53ae4ed9904df42e3f81c634['h036f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b7b] =  I0310077d53ae4ed9904df42e3f81c634['h036f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b7c] =  I0310077d53ae4ed9904df42e3f81c634['h036f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b7d] =  I0310077d53ae4ed9904df42e3f81c634['h036fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b7e] =  I0310077d53ae4ed9904df42e3f81c634['h036fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b7f] =  I0310077d53ae4ed9904df42e3f81c634['h036fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b80] =  I0310077d53ae4ed9904df42e3f81c634['h03700] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b81] =  I0310077d53ae4ed9904df42e3f81c634['h03702] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b82] =  I0310077d53ae4ed9904df42e3f81c634['h03704] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b83] =  I0310077d53ae4ed9904df42e3f81c634['h03706] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b84] =  I0310077d53ae4ed9904df42e3f81c634['h03708] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b85] =  I0310077d53ae4ed9904df42e3f81c634['h0370a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b86] =  I0310077d53ae4ed9904df42e3f81c634['h0370c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b87] =  I0310077d53ae4ed9904df42e3f81c634['h0370e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b88] =  I0310077d53ae4ed9904df42e3f81c634['h03710] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b89] =  I0310077d53ae4ed9904df42e3f81c634['h03712] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b8a] =  I0310077d53ae4ed9904df42e3f81c634['h03714] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b8b] =  I0310077d53ae4ed9904df42e3f81c634['h03716] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b8c] =  I0310077d53ae4ed9904df42e3f81c634['h03718] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b8d] =  I0310077d53ae4ed9904df42e3f81c634['h0371a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b8e] =  I0310077d53ae4ed9904df42e3f81c634['h0371c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b8f] =  I0310077d53ae4ed9904df42e3f81c634['h0371e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b90] =  I0310077d53ae4ed9904df42e3f81c634['h03720] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b91] =  I0310077d53ae4ed9904df42e3f81c634['h03722] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b92] =  I0310077d53ae4ed9904df42e3f81c634['h03724] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b93] =  I0310077d53ae4ed9904df42e3f81c634['h03726] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b94] =  I0310077d53ae4ed9904df42e3f81c634['h03728] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b95] =  I0310077d53ae4ed9904df42e3f81c634['h0372a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b96] =  I0310077d53ae4ed9904df42e3f81c634['h0372c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b97] =  I0310077d53ae4ed9904df42e3f81c634['h0372e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b98] =  I0310077d53ae4ed9904df42e3f81c634['h03730] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b99] =  I0310077d53ae4ed9904df42e3f81c634['h03732] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b9a] =  I0310077d53ae4ed9904df42e3f81c634['h03734] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b9b] =  I0310077d53ae4ed9904df42e3f81c634['h03736] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b9c] =  I0310077d53ae4ed9904df42e3f81c634['h03738] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b9d] =  I0310077d53ae4ed9904df42e3f81c634['h0373a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b9e] =  I0310077d53ae4ed9904df42e3f81c634['h0373c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01b9f] =  I0310077d53ae4ed9904df42e3f81c634['h0373e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba0] =  I0310077d53ae4ed9904df42e3f81c634['h03740] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba1] =  I0310077d53ae4ed9904df42e3f81c634['h03742] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba2] =  I0310077d53ae4ed9904df42e3f81c634['h03744] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba3] =  I0310077d53ae4ed9904df42e3f81c634['h03746] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba4] =  I0310077d53ae4ed9904df42e3f81c634['h03748] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba5] =  I0310077d53ae4ed9904df42e3f81c634['h0374a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba6] =  I0310077d53ae4ed9904df42e3f81c634['h0374c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba7] =  I0310077d53ae4ed9904df42e3f81c634['h0374e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba8] =  I0310077d53ae4ed9904df42e3f81c634['h03750] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ba9] =  I0310077d53ae4ed9904df42e3f81c634['h03752] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01baa] =  I0310077d53ae4ed9904df42e3f81c634['h03754] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bab] =  I0310077d53ae4ed9904df42e3f81c634['h03756] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bac] =  I0310077d53ae4ed9904df42e3f81c634['h03758] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bad] =  I0310077d53ae4ed9904df42e3f81c634['h0375a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bae] =  I0310077d53ae4ed9904df42e3f81c634['h0375c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01baf] =  I0310077d53ae4ed9904df42e3f81c634['h0375e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb0] =  I0310077d53ae4ed9904df42e3f81c634['h03760] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb1] =  I0310077d53ae4ed9904df42e3f81c634['h03762] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb2] =  I0310077d53ae4ed9904df42e3f81c634['h03764] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb3] =  I0310077d53ae4ed9904df42e3f81c634['h03766] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb4] =  I0310077d53ae4ed9904df42e3f81c634['h03768] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb5] =  I0310077d53ae4ed9904df42e3f81c634['h0376a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb6] =  I0310077d53ae4ed9904df42e3f81c634['h0376c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb7] =  I0310077d53ae4ed9904df42e3f81c634['h0376e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb8] =  I0310077d53ae4ed9904df42e3f81c634['h03770] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bb9] =  I0310077d53ae4ed9904df42e3f81c634['h03772] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bba] =  I0310077d53ae4ed9904df42e3f81c634['h03774] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bbb] =  I0310077d53ae4ed9904df42e3f81c634['h03776] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bbc] =  I0310077d53ae4ed9904df42e3f81c634['h03778] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bbd] =  I0310077d53ae4ed9904df42e3f81c634['h0377a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bbe] =  I0310077d53ae4ed9904df42e3f81c634['h0377c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bbf] =  I0310077d53ae4ed9904df42e3f81c634['h0377e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc0] =  I0310077d53ae4ed9904df42e3f81c634['h03780] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc1] =  I0310077d53ae4ed9904df42e3f81c634['h03782] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc2] =  I0310077d53ae4ed9904df42e3f81c634['h03784] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc3] =  I0310077d53ae4ed9904df42e3f81c634['h03786] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc4] =  I0310077d53ae4ed9904df42e3f81c634['h03788] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc5] =  I0310077d53ae4ed9904df42e3f81c634['h0378a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc6] =  I0310077d53ae4ed9904df42e3f81c634['h0378c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc7] =  I0310077d53ae4ed9904df42e3f81c634['h0378e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc8] =  I0310077d53ae4ed9904df42e3f81c634['h03790] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bc9] =  I0310077d53ae4ed9904df42e3f81c634['h03792] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bca] =  I0310077d53ae4ed9904df42e3f81c634['h03794] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bcb] =  I0310077d53ae4ed9904df42e3f81c634['h03796] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bcc] =  I0310077d53ae4ed9904df42e3f81c634['h03798] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bcd] =  I0310077d53ae4ed9904df42e3f81c634['h0379a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bce] =  I0310077d53ae4ed9904df42e3f81c634['h0379c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bcf] =  I0310077d53ae4ed9904df42e3f81c634['h0379e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd0] =  I0310077d53ae4ed9904df42e3f81c634['h037a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd1] =  I0310077d53ae4ed9904df42e3f81c634['h037a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd2] =  I0310077d53ae4ed9904df42e3f81c634['h037a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd3] =  I0310077d53ae4ed9904df42e3f81c634['h037a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd4] =  I0310077d53ae4ed9904df42e3f81c634['h037a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd5] =  I0310077d53ae4ed9904df42e3f81c634['h037aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd6] =  I0310077d53ae4ed9904df42e3f81c634['h037ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd7] =  I0310077d53ae4ed9904df42e3f81c634['h037ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd8] =  I0310077d53ae4ed9904df42e3f81c634['h037b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bd9] =  I0310077d53ae4ed9904df42e3f81c634['h037b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bda] =  I0310077d53ae4ed9904df42e3f81c634['h037b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bdb] =  I0310077d53ae4ed9904df42e3f81c634['h037b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bdc] =  I0310077d53ae4ed9904df42e3f81c634['h037b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bdd] =  I0310077d53ae4ed9904df42e3f81c634['h037ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bde] =  I0310077d53ae4ed9904df42e3f81c634['h037bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bdf] =  I0310077d53ae4ed9904df42e3f81c634['h037be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be0] =  I0310077d53ae4ed9904df42e3f81c634['h037c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be1] =  I0310077d53ae4ed9904df42e3f81c634['h037c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be2] =  I0310077d53ae4ed9904df42e3f81c634['h037c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be3] =  I0310077d53ae4ed9904df42e3f81c634['h037c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be4] =  I0310077d53ae4ed9904df42e3f81c634['h037c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be5] =  I0310077d53ae4ed9904df42e3f81c634['h037ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be6] =  I0310077d53ae4ed9904df42e3f81c634['h037cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be7] =  I0310077d53ae4ed9904df42e3f81c634['h037ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be8] =  I0310077d53ae4ed9904df42e3f81c634['h037d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01be9] =  I0310077d53ae4ed9904df42e3f81c634['h037d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bea] =  I0310077d53ae4ed9904df42e3f81c634['h037d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01beb] =  I0310077d53ae4ed9904df42e3f81c634['h037d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bec] =  I0310077d53ae4ed9904df42e3f81c634['h037d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bed] =  I0310077d53ae4ed9904df42e3f81c634['h037da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bee] =  I0310077d53ae4ed9904df42e3f81c634['h037dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bef] =  I0310077d53ae4ed9904df42e3f81c634['h037de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf0] =  I0310077d53ae4ed9904df42e3f81c634['h037e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf1] =  I0310077d53ae4ed9904df42e3f81c634['h037e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf2] =  I0310077d53ae4ed9904df42e3f81c634['h037e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf3] =  I0310077d53ae4ed9904df42e3f81c634['h037e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf4] =  I0310077d53ae4ed9904df42e3f81c634['h037e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf5] =  I0310077d53ae4ed9904df42e3f81c634['h037ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf6] =  I0310077d53ae4ed9904df42e3f81c634['h037ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf7] =  I0310077d53ae4ed9904df42e3f81c634['h037ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf8] =  I0310077d53ae4ed9904df42e3f81c634['h037f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bf9] =  I0310077d53ae4ed9904df42e3f81c634['h037f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bfa] =  I0310077d53ae4ed9904df42e3f81c634['h037f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bfb] =  I0310077d53ae4ed9904df42e3f81c634['h037f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bfc] =  I0310077d53ae4ed9904df42e3f81c634['h037f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bfd] =  I0310077d53ae4ed9904df42e3f81c634['h037fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bfe] =  I0310077d53ae4ed9904df42e3f81c634['h037fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01bff] =  I0310077d53ae4ed9904df42e3f81c634['h037fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c00] =  I0310077d53ae4ed9904df42e3f81c634['h03800] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c01] =  I0310077d53ae4ed9904df42e3f81c634['h03802] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c02] =  I0310077d53ae4ed9904df42e3f81c634['h03804] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c03] =  I0310077d53ae4ed9904df42e3f81c634['h03806] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c04] =  I0310077d53ae4ed9904df42e3f81c634['h03808] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c05] =  I0310077d53ae4ed9904df42e3f81c634['h0380a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c06] =  I0310077d53ae4ed9904df42e3f81c634['h0380c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c07] =  I0310077d53ae4ed9904df42e3f81c634['h0380e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c08] =  I0310077d53ae4ed9904df42e3f81c634['h03810] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c09] =  I0310077d53ae4ed9904df42e3f81c634['h03812] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c0a] =  I0310077d53ae4ed9904df42e3f81c634['h03814] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c0b] =  I0310077d53ae4ed9904df42e3f81c634['h03816] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c0c] =  I0310077d53ae4ed9904df42e3f81c634['h03818] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c0d] =  I0310077d53ae4ed9904df42e3f81c634['h0381a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c0e] =  I0310077d53ae4ed9904df42e3f81c634['h0381c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c0f] =  I0310077d53ae4ed9904df42e3f81c634['h0381e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c10] =  I0310077d53ae4ed9904df42e3f81c634['h03820] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c11] =  I0310077d53ae4ed9904df42e3f81c634['h03822] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c12] =  I0310077d53ae4ed9904df42e3f81c634['h03824] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c13] =  I0310077d53ae4ed9904df42e3f81c634['h03826] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c14] =  I0310077d53ae4ed9904df42e3f81c634['h03828] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c15] =  I0310077d53ae4ed9904df42e3f81c634['h0382a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c16] =  I0310077d53ae4ed9904df42e3f81c634['h0382c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c17] =  I0310077d53ae4ed9904df42e3f81c634['h0382e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c18] =  I0310077d53ae4ed9904df42e3f81c634['h03830] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c19] =  I0310077d53ae4ed9904df42e3f81c634['h03832] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c1a] =  I0310077d53ae4ed9904df42e3f81c634['h03834] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c1b] =  I0310077d53ae4ed9904df42e3f81c634['h03836] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c1c] =  I0310077d53ae4ed9904df42e3f81c634['h03838] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c1d] =  I0310077d53ae4ed9904df42e3f81c634['h0383a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c1e] =  I0310077d53ae4ed9904df42e3f81c634['h0383c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c1f] =  I0310077d53ae4ed9904df42e3f81c634['h0383e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c20] =  I0310077d53ae4ed9904df42e3f81c634['h03840] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c21] =  I0310077d53ae4ed9904df42e3f81c634['h03842] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c22] =  I0310077d53ae4ed9904df42e3f81c634['h03844] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c23] =  I0310077d53ae4ed9904df42e3f81c634['h03846] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c24] =  I0310077d53ae4ed9904df42e3f81c634['h03848] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c25] =  I0310077d53ae4ed9904df42e3f81c634['h0384a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c26] =  I0310077d53ae4ed9904df42e3f81c634['h0384c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c27] =  I0310077d53ae4ed9904df42e3f81c634['h0384e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c28] =  I0310077d53ae4ed9904df42e3f81c634['h03850] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c29] =  I0310077d53ae4ed9904df42e3f81c634['h03852] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c2a] =  I0310077d53ae4ed9904df42e3f81c634['h03854] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c2b] =  I0310077d53ae4ed9904df42e3f81c634['h03856] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c2c] =  I0310077d53ae4ed9904df42e3f81c634['h03858] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c2d] =  I0310077d53ae4ed9904df42e3f81c634['h0385a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c2e] =  I0310077d53ae4ed9904df42e3f81c634['h0385c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c2f] =  I0310077d53ae4ed9904df42e3f81c634['h0385e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c30] =  I0310077d53ae4ed9904df42e3f81c634['h03860] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c31] =  I0310077d53ae4ed9904df42e3f81c634['h03862] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c32] =  I0310077d53ae4ed9904df42e3f81c634['h03864] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c33] =  I0310077d53ae4ed9904df42e3f81c634['h03866] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c34] =  I0310077d53ae4ed9904df42e3f81c634['h03868] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c35] =  I0310077d53ae4ed9904df42e3f81c634['h0386a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c36] =  I0310077d53ae4ed9904df42e3f81c634['h0386c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c37] =  I0310077d53ae4ed9904df42e3f81c634['h0386e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c38] =  I0310077d53ae4ed9904df42e3f81c634['h03870] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c39] =  I0310077d53ae4ed9904df42e3f81c634['h03872] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c3a] =  I0310077d53ae4ed9904df42e3f81c634['h03874] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c3b] =  I0310077d53ae4ed9904df42e3f81c634['h03876] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c3c] =  I0310077d53ae4ed9904df42e3f81c634['h03878] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c3d] =  I0310077d53ae4ed9904df42e3f81c634['h0387a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c3e] =  I0310077d53ae4ed9904df42e3f81c634['h0387c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c3f] =  I0310077d53ae4ed9904df42e3f81c634['h0387e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c40] =  I0310077d53ae4ed9904df42e3f81c634['h03880] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c41] =  I0310077d53ae4ed9904df42e3f81c634['h03882] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c42] =  I0310077d53ae4ed9904df42e3f81c634['h03884] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c43] =  I0310077d53ae4ed9904df42e3f81c634['h03886] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c44] =  I0310077d53ae4ed9904df42e3f81c634['h03888] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c45] =  I0310077d53ae4ed9904df42e3f81c634['h0388a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c46] =  I0310077d53ae4ed9904df42e3f81c634['h0388c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c47] =  I0310077d53ae4ed9904df42e3f81c634['h0388e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c48] =  I0310077d53ae4ed9904df42e3f81c634['h03890] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c49] =  I0310077d53ae4ed9904df42e3f81c634['h03892] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c4a] =  I0310077d53ae4ed9904df42e3f81c634['h03894] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c4b] =  I0310077d53ae4ed9904df42e3f81c634['h03896] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c4c] =  I0310077d53ae4ed9904df42e3f81c634['h03898] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c4d] =  I0310077d53ae4ed9904df42e3f81c634['h0389a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c4e] =  I0310077d53ae4ed9904df42e3f81c634['h0389c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c4f] =  I0310077d53ae4ed9904df42e3f81c634['h0389e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c50] =  I0310077d53ae4ed9904df42e3f81c634['h038a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c51] =  I0310077d53ae4ed9904df42e3f81c634['h038a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c52] =  I0310077d53ae4ed9904df42e3f81c634['h038a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c53] =  I0310077d53ae4ed9904df42e3f81c634['h038a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c54] =  I0310077d53ae4ed9904df42e3f81c634['h038a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c55] =  I0310077d53ae4ed9904df42e3f81c634['h038aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c56] =  I0310077d53ae4ed9904df42e3f81c634['h038ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c57] =  I0310077d53ae4ed9904df42e3f81c634['h038ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c58] =  I0310077d53ae4ed9904df42e3f81c634['h038b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c59] =  I0310077d53ae4ed9904df42e3f81c634['h038b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c5a] =  I0310077d53ae4ed9904df42e3f81c634['h038b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c5b] =  I0310077d53ae4ed9904df42e3f81c634['h038b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c5c] =  I0310077d53ae4ed9904df42e3f81c634['h038b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c5d] =  I0310077d53ae4ed9904df42e3f81c634['h038ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c5e] =  I0310077d53ae4ed9904df42e3f81c634['h038bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c5f] =  I0310077d53ae4ed9904df42e3f81c634['h038be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c60] =  I0310077d53ae4ed9904df42e3f81c634['h038c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c61] =  I0310077d53ae4ed9904df42e3f81c634['h038c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c62] =  I0310077d53ae4ed9904df42e3f81c634['h038c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c63] =  I0310077d53ae4ed9904df42e3f81c634['h038c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c64] =  I0310077d53ae4ed9904df42e3f81c634['h038c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c65] =  I0310077d53ae4ed9904df42e3f81c634['h038ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c66] =  I0310077d53ae4ed9904df42e3f81c634['h038cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c67] =  I0310077d53ae4ed9904df42e3f81c634['h038ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c68] =  I0310077d53ae4ed9904df42e3f81c634['h038d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c69] =  I0310077d53ae4ed9904df42e3f81c634['h038d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c6a] =  I0310077d53ae4ed9904df42e3f81c634['h038d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c6b] =  I0310077d53ae4ed9904df42e3f81c634['h038d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c6c] =  I0310077d53ae4ed9904df42e3f81c634['h038d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c6d] =  I0310077d53ae4ed9904df42e3f81c634['h038da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c6e] =  I0310077d53ae4ed9904df42e3f81c634['h038dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c6f] =  I0310077d53ae4ed9904df42e3f81c634['h038de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c70] =  I0310077d53ae4ed9904df42e3f81c634['h038e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c71] =  I0310077d53ae4ed9904df42e3f81c634['h038e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c72] =  I0310077d53ae4ed9904df42e3f81c634['h038e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c73] =  I0310077d53ae4ed9904df42e3f81c634['h038e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c74] =  I0310077d53ae4ed9904df42e3f81c634['h038e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c75] =  I0310077d53ae4ed9904df42e3f81c634['h038ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c76] =  I0310077d53ae4ed9904df42e3f81c634['h038ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c77] =  I0310077d53ae4ed9904df42e3f81c634['h038ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c78] =  I0310077d53ae4ed9904df42e3f81c634['h038f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c79] =  I0310077d53ae4ed9904df42e3f81c634['h038f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c7a] =  I0310077d53ae4ed9904df42e3f81c634['h038f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c7b] =  I0310077d53ae4ed9904df42e3f81c634['h038f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c7c] =  I0310077d53ae4ed9904df42e3f81c634['h038f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c7d] =  I0310077d53ae4ed9904df42e3f81c634['h038fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c7e] =  I0310077d53ae4ed9904df42e3f81c634['h038fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c7f] =  I0310077d53ae4ed9904df42e3f81c634['h038fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c80] =  I0310077d53ae4ed9904df42e3f81c634['h03900] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c81] =  I0310077d53ae4ed9904df42e3f81c634['h03902] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c82] =  I0310077d53ae4ed9904df42e3f81c634['h03904] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c83] =  I0310077d53ae4ed9904df42e3f81c634['h03906] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c84] =  I0310077d53ae4ed9904df42e3f81c634['h03908] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c85] =  I0310077d53ae4ed9904df42e3f81c634['h0390a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c86] =  I0310077d53ae4ed9904df42e3f81c634['h0390c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c87] =  I0310077d53ae4ed9904df42e3f81c634['h0390e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c88] =  I0310077d53ae4ed9904df42e3f81c634['h03910] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c89] =  I0310077d53ae4ed9904df42e3f81c634['h03912] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c8a] =  I0310077d53ae4ed9904df42e3f81c634['h03914] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c8b] =  I0310077d53ae4ed9904df42e3f81c634['h03916] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c8c] =  I0310077d53ae4ed9904df42e3f81c634['h03918] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c8d] =  I0310077d53ae4ed9904df42e3f81c634['h0391a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c8e] =  I0310077d53ae4ed9904df42e3f81c634['h0391c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c8f] =  I0310077d53ae4ed9904df42e3f81c634['h0391e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c90] =  I0310077d53ae4ed9904df42e3f81c634['h03920] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c91] =  I0310077d53ae4ed9904df42e3f81c634['h03922] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c92] =  I0310077d53ae4ed9904df42e3f81c634['h03924] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c93] =  I0310077d53ae4ed9904df42e3f81c634['h03926] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c94] =  I0310077d53ae4ed9904df42e3f81c634['h03928] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c95] =  I0310077d53ae4ed9904df42e3f81c634['h0392a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c96] =  I0310077d53ae4ed9904df42e3f81c634['h0392c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c97] =  I0310077d53ae4ed9904df42e3f81c634['h0392e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c98] =  I0310077d53ae4ed9904df42e3f81c634['h03930] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c99] =  I0310077d53ae4ed9904df42e3f81c634['h03932] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c9a] =  I0310077d53ae4ed9904df42e3f81c634['h03934] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c9b] =  I0310077d53ae4ed9904df42e3f81c634['h03936] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c9c] =  I0310077d53ae4ed9904df42e3f81c634['h03938] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c9d] =  I0310077d53ae4ed9904df42e3f81c634['h0393a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c9e] =  I0310077d53ae4ed9904df42e3f81c634['h0393c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01c9f] =  I0310077d53ae4ed9904df42e3f81c634['h0393e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca0] =  I0310077d53ae4ed9904df42e3f81c634['h03940] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca1] =  I0310077d53ae4ed9904df42e3f81c634['h03942] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca2] =  I0310077d53ae4ed9904df42e3f81c634['h03944] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca3] =  I0310077d53ae4ed9904df42e3f81c634['h03946] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca4] =  I0310077d53ae4ed9904df42e3f81c634['h03948] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca5] =  I0310077d53ae4ed9904df42e3f81c634['h0394a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca6] =  I0310077d53ae4ed9904df42e3f81c634['h0394c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca7] =  I0310077d53ae4ed9904df42e3f81c634['h0394e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca8] =  I0310077d53ae4ed9904df42e3f81c634['h03950] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ca9] =  I0310077d53ae4ed9904df42e3f81c634['h03952] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01caa] =  I0310077d53ae4ed9904df42e3f81c634['h03954] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cab] =  I0310077d53ae4ed9904df42e3f81c634['h03956] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cac] =  I0310077d53ae4ed9904df42e3f81c634['h03958] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cad] =  I0310077d53ae4ed9904df42e3f81c634['h0395a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cae] =  I0310077d53ae4ed9904df42e3f81c634['h0395c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01caf] =  I0310077d53ae4ed9904df42e3f81c634['h0395e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb0] =  I0310077d53ae4ed9904df42e3f81c634['h03960] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb1] =  I0310077d53ae4ed9904df42e3f81c634['h03962] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb2] =  I0310077d53ae4ed9904df42e3f81c634['h03964] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb3] =  I0310077d53ae4ed9904df42e3f81c634['h03966] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb4] =  I0310077d53ae4ed9904df42e3f81c634['h03968] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb5] =  I0310077d53ae4ed9904df42e3f81c634['h0396a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb6] =  I0310077d53ae4ed9904df42e3f81c634['h0396c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb7] =  I0310077d53ae4ed9904df42e3f81c634['h0396e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb8] =  I0310077d53ae4ed9904df42e3f81c634['h03970] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cb9] =  I0310077d53ae4ed9904df42e3f81c634['h03972] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cba] =  I0310077d53ae4ed9904df42e3f81c634['h03974] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cbb] =  I0310077d53ae4ed9904df42e3f81c634['h03976] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cbc] =  I0310077d53ae4ed9904df42e3f81c634['h03978] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cbd] =  I0310077d53ae4ed9904df42e3f81c634['h0397a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cbe] =  I0310077d53ae4ed9904df42e3f81c634['h0397c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cbf] =  I0310077d53ae4ed9904df42e3f81c634['h0397e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc0] =  I0310077d53ae4ed9904df42e3f81c634['h03980] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc1] =  I0310077d53ae4ed9904df42e3f81c634['h03982] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc2] =  I0310077d53ae4ed9904df42e3f81c634['h03984] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc3] =  I0310077d53ae4ed9904df42e3f81c634['h03986] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc4] =  I0310077d53ae4ed9904df42e3f81c634['h03988] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc5] =  I0310077d53ae4ed9904df42e3f81c634['h0398a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc6] =  I0310077d53ae4ed9904df42e3f81c634['h0398c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc7] =  I0310077d53ae4ed9904df42e3f81c634['h0398e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc8] =  I0310077d53ae4ed9904df42e3f81c634['h03990] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cc9] =  I0310077d53ae4ed9904df42e3f81c634['h03992] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cca] =  I0310077d53ae4ed9904df42e3f81c634['h03994] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ccb] =  I0310077d53ae4ed9904df42e3f81c634['h03996] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ccc] =  I0310077d53ae4ed9904df42e3f81c634['h03998] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ccd] =  I0310077d53ae4ed9904df42e3f81c634['h0399a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cce] =  I0310077d53ae4ed9904df42e3f81c634['h0399c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ccf] =  I0310077d53ae4ed9904df42e3f81c634['h0399e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd0] =  I0310077d53ae4ed9904df42e3f81c634['h039a0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd1] =  I0310077d53ae4ed9904df42e3f81c634['h039a2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd2] =  I0310077d53ae4ed9904df42e3f81c634['h039a4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd3] =  I0310077d53ae4ed9904df42e3f81c634['h039a6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd4] =  I0310077d53ae4ed9904df42e3f81c634['h039a8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd5] =  I0310077d53ae4ed9904df42e3f81c634['h039aa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd6] =  I0310077d53ae4ed9904df42e3f81c634['h039ac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd7] =  I0310077d53ae4ed9904df42e3f81c634['h039ae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd8] =  I0310077d53ae4ed9904df42e3f81c634['h039b0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cd9] =  I0310077d53ae4ed9904df42e3f81c634['h039b2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cda] =  I0310077d53ae4ed9904df42e3f81c634['h039b4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cdb] =  I0310077d53ae4ed9904df42e3f81c634['h039b6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cdc] =  I0310077d53ae4ed9904df42e3f81c634['h039b8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cdd] =  I0310077d53ae4ed9904df42e3f81c634['h039ba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cde] =  I0310077d53ae4ed9904df42e3f81c634['h039bc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cdf] =  I0310077d53ae4ed9904df42e3f81c634['h039be] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce0] =  I0310077d53ae4ed9904df42e3f81c634['h039c0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce1] =  I0310077d53ae4ed9904df42e3f81c634['h039c2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce2] =  I0310077d53ae4ed9904df42e3f81c634['h039c4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce3] =  I0310077d53ae4ed9904df42e3f81c634['h039c6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce4] =  I0310077d53ae4ed9904df42e3f81c634['h039c8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce5] =  I0310077d53ae4ed9904df42e3f81c634['h039ca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce6] =  I0310077d53ae4ed9904df42e3f81c634['h039cc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce7] =  I0310077d53ae4ed9904df42e3f81c634['h039ce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce8] =  I0310077d53ae4ed9904df42e3f81c634['h039d0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ce9] =  I0310077d53ae4ed9904df42e3f81c634['h039d2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cea] =  I0310077d53ae4ed9904df42e3f81c634['h039d4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ceb] =  I0310077d53ae4ed9904df42e3f81c634['h039d6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cec] =  I0310077d53ae4ed9904df42e3f81c634['h039d8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ced] =  I0310077d53ae4ed9904df42e3f81c634['h039da] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cee] =  I0310077d53ae4ed9904df42e3f81c634['h039dc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cef] =  I0310077d53ae4ed9904df42e3f81c634['h039de] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf0] =  I0310077d53ae4ed9904df42e3f81c634['h039e0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf1] =  I0310077d53ae4ed9904df42e3f81c634['h039e2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf2] =  I0310077d53ae4ed9904df42e3f81c634['h039e4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf3] =  I0310077d53ae4ed9904df42e3f81c634['h039e6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf4] =  I0310077d53ae4ed9904df42e3f81c634['h039e8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf5] =  I0310077d53ae4ed9904df42e3f81c634['h039ea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf6] =  I0310077d53ae4ed9904df42e3f81c634['h039ec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf7] =  I0310077d53ae4ed9904df42e3f81c634['h039ee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf8] =  I0310077d53ae4ed9904df42e3f81c634['h039f0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cf9] =  I0310077d53ae4ed9904df42e3f81c634['h039f2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cfa] =  I0310077d53ae4ed9904df42e3f81c634['h039f4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cfb] =  I0310077d53ae4ed9904df42e3f81c634['h039f6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cfc] =  I0310077d53ae4ed9904df42e3f81c634['h039f8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cfd] =  I0310077d53ae4ed9904df42e3f81c634['h039fa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cfe] =  I0310077d53ae4ed9904df42e3f81c634['h039fc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01cff] =  I0310077d53ae4ed9904df42e3f81c634['h039fe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d00] =  I0310077d53ae4ed9904df42e3f81c634['h03a00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d01] =  I0310077d53ae4ed9904df42e3f81c634['h03a02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d02] =  I0310077d53ae4ed9904df42e3f81c634['h03a04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d03] =  I0310077d53ae4ed9904df42e3f81c634['h03a06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d04] =  I0310077d53ae4ed9904df42e3f81c634['h03a08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d05] =  I0310077d53ae4ed9904df42e3f81c634['h03a0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d06] =  I0310077d53ae4ed9904df42e3f81c634['h03a0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d07] =  I0310077d53ae4ed9904df42e3f81c634['h03a0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d08] =  I0310077d53ae4ed9904df42e3f81c634['h03a10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d09] =  I0310077d53ae4ed9904df42e3f81c634['h03a12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d0a] =  I0310077d53ae4ed9904df42e3f81c634['h03a14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d0b] =  I0310077d53ae4ed9904df42e3f81c634['h03a16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d0c] =  I0310077d53ae4ed9904df42e3f81c634['h03a18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d0d] =  I0310077d53ae4ed9904df42e3f81c634['h03a1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d0e] =  I0310077d53ae4ed9904df42e3f81c634['h03a1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d0f] =  I0310077d53ae4ed9904df42e3f81c634['h03a1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d10] =  I0310077d53ae4ed9904df42e3f81c634['h03a20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d11] =  I0310077d53ae4ed9904df42e3f81c634['h03a22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d12] =  I0310077d53ae4ed9904df42e3f81c634['h03a24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d13] =  I0310077d53ae4ed9904df42e3f81c634['h03a26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d14] =  I0310077d53ae4ed9904df42e3f81c634['h03a28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d15] =  I0310077d53ae4ed9904df42e3f81c634['h03a2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d16] =  I0310077d53ae4ed9904df42e3f81c634['h03a2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d17] =  I0310077d53ae4ed9904df42e3f81c634['h03a2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d18] =  I0310077d53ae4ed9904df42e3f81c634['h03a30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d19] =  I0310077d53ae4ed9904df42e3f81c634['h03a32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d1a] =  I0310077d53ae4ed9904df42e3f81c634['h03a34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d1b] =  I0310077d53ae4ed9904df42e3f81c634['h03a36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d1c] =  I0310077d53ae4ed9904df42e3f81c634['h03a38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d1d] =  I0310077d53ae4ed9904df42e3f81c634['h03a3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d1e] =  I0310077d53ae4ed9904df42e3f81c634['h03a3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d1f] =  I0310077d53ae4ed9904df42e3f81c634['h03a3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d20] =  I0310077d53ae4ed9904df42e3f81c634['h03a40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d21] =  I0310077d53ae4ed9904df42e3f81c634['h03a42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d22] =  I0310077d53ae4ed9904df42e3f81c634['h03a44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d23] =  I0310077d53ae4ed9904df42e3f81c634['h03a46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d24] =  I0310077d53ae4ed9904df42e3f81c634['h03a48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d25] =  I0310077d53ae4ed9904df42e3f81c634['h03a4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d26] =  I0310077d53ae4ed9904df42e3f81c634['h03a4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d27] =  I0310077d53ae4ed9904df42e3f81c634['h03a4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d28] =  I0310077d53ae4ed9904df42e3f81c634['h03a50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d29] =  I0310077d53ae4ed9904df42e3f81c634['h03a52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d2a] =  I0310077d53ae4ed9904df42e3f81c634['h03a54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d2b] =  I0310077d53ae4ed9904df42e3f81c634['h03a56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d2c] =  I0310077d53ae4ed9904df42e3f81c634['h03a58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d2d] =  I0310077d53ae4ed9904df42e3f81c634['h03a5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d2e] =  I0310077d53ae4ed9904df42e3f81c634['h03a5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d2f] =  I0310077d53ae4ed9904df42e3f81c634['h03a5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d30] =  I0310077d53ae4ed9904df42e3f81c634['h03a60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d31] =  I0310077d53ae4ed9904df42e3f81c634['h03a62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d32] =  I0310077d53ae4ed9904df42e3f81c634['h03a64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d33] =  I0310077d53ae4ed9904df42e3f81c634['h03a66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d34] =  I0310077d53ae4ed9904df42e3f81c634['h03a68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d35] =  I0310077d53ae4ed9904df42e3f81c634['h03a6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d36] =  I0310077d53ae4ed9904df42e3f81c634['h03a6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d37] =  I0310077d53ae4ed9904df42e3f81c634['h03a6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d38] =  I0310077d53ae4ed9904df42e3f81c634['h03a70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d39] =  I0310077d53ae4ed9904df42e3f81c634['h03a72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d3a] =  I0310077d53ae4ed9904df42e3f81c634['h03a74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d3b] =  I0310077d53ae4ed9904df42e3f81c634['h03a76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d3c] =  I0310077d53ae4ed9904df42e3f81c634['h03a78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d3d] =  I0310077d53ae4ed9904df42e3f81c634['h03a7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d3e] =  I0310077d53ae4ed9904df42e3f81c634['h03a7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d3f] =  I0310077d53ae4ed9904df42e3f81c634['h03a7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d40] =  I0310077d53ae4ed9904df42e3f81c634['h03a80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d41] =  I0310077d53ae4ed9904df42e3f81c634['h03a82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d42] =  I0310077d53ae4ed9904df42e3f81c634['h03a84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d43] =  I0310077d53ae4ed9904df42e3f81c634['h03a86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d44] =  I0310077d53ae4ed9904df42e3f81c634['h03a88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d45] =  I0310077d53ae4ed9904df42e3f81c634['h03a8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d46] =  I0310077d53ae4ed9904df42e3f81c634['h03a8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d47] =  I0310077d53ae4ed9904df42e3f81c634['h03a8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d48] =  I0310077d53ae4ed9904df42e3f81c634['h03a90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d49] =  I0310077d53ae4ed9904df42e3f81c634['h03a92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d4a] =  I0310077d53ae4ed9904df42e3f81c634['h03a94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d4b] =  I0310077d53ae4ed9904df42e3f81c634['h03a96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d4c] =  I0310077d53ae4ed9904df42e3f81c634['h03a98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d4d] =  I0310077d53ae4ed9904df42e3f81c634['h03a9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d4e] =  I0310077d53ae4ed9904df42e3f81c634['h03a9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d4f] =  I0310077d53ae4ed9904df42e3f81c634['h03a9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d50] =  I0310077d53ae4ed9904df42e3f81c634['h03aa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d51] =  I0310077d53ae4ed9904df42e3f81c634['h03aa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d52] =  I0310077d53ae4ed9904df42e3f81c634['h03aa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d53] =  I0310077d53ae4ed9904df42e3f81c634['h03aa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d54] =  I0310077d53ae4ed9904df42e3f81c634['h03aa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d55] =  I0310077d53ae4ed9904df42e3f81c634['h03aaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d56] =  I0310077d53ae4ed9904df42e3f81c634['h03aac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d57] =  I0310077d53ae4ed9904df42e3f81c634['h03aae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d58] =  I0310077d53ae4ed9904df42e3f81c634['h03ab0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d59] =  I0310077d53ae4ed9904df42e3f81c634['h03ab2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d5a] =  I0310077d53ae4ed9904df42e3f81c634['h03ab4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d5b] =  I0310077d53ae4ed9904df42e3f81c634['h03ab6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d5c] =  I0310077d53ae4ed9904df42e3f81c634['h03ab8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d5d] =  I0310077d53ae4ed9904df42e3f81c634['h03aba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d5e] =  I0310077d53ae4ed9904df42e3f81c634['h03abc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d5f] =  I0310077d53ae4ed9904df42e3f81c634['h03abe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d60] =  I0310077d53ae4ed9904df42e3f81c634['h03ac0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d61] =  I0310077d53ae4ed9904df42e3f81c634['h03ac2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d62] =  I0310077d53ae4ed9904df42e3f81c634['h03ac4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d63] =  I0310077d53ae4ed9904df42e3f81c634['h03ac6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d64] =  I0310077d53ae4ed9904df42e3f81c634['h03ac8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d65] =  I0310077d53ae4ed9904df42e3f81c634['h03aca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d66] =  I0310077d53ae4ed9904df42e3f81c634['h03acc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d67] =  I0310077d53ae4ed9904df42e3f81c634['h03ace] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d68] =  I0310077d53ae4ed9904df42e3f81c634['h03ad0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d69] =  I0310077d53ae4ed9904df42e3f81c634['h03ad2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d6a] =  I0310077d53ae4ed9904df42e3f81c634['h03ad4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d6b] =  I0310077d53ae4ed9904df42e3f81c634['h03ad6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d6c] =  I0310077d53ae4ed9904df42e3f81c634['h03ad8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d6d] =  I0310077d53ae4ed9904df42e3f81c634['h03ada] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d6e] =  I0310077d53ae4ed9904df42e3f81c634['h03adc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d6f] =  I0310077d53ae4ed9904df42e3f81c634['h03ade] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d70] =  I0310077d53ae4ed9904df42e3f81c634['h03ae0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d71] =  I0310077d53ae4ed9904df42e3f81c634['h03ae2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d72] =  I0310077d53ae4ed9904df42e3f81c634['h03ae4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d73] =  I0310077d53ae4ed9904df42e3f81c634['h03ae6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d74] =  I0310077d53ae4ed9904df42e3f81c634['h03ae8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d75] =  I0310077d53ae4ed9904df42e3f81c634['h03aea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d76] =  I0310077d53ae4ed9904df42e3f81c634['h03aec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d77] =  I0310077d53ae4ed9904df42e3f81c634['h03aee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d78] =  I0310077d53ae4ed9904df42e3f81c634['h03af0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d79] =  I0310077d53ae4ed9904df42e3f81c634['h03af2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d7a] =  I0310077d53ae4ed9904df42e3f81c634['h03af4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d7b] =  I0310077d53ae4ed9904df42e3f81c634['h03af6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d7c] =  I0310077d53ae4ed9904df42e3f81c634['h03af8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d7d] =  I0310077d53ae4ed9904df42e3f81c634['h03afa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d7e] =  I0310077d53ae4ed9904df42e3f81c634['h03afc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d7f] =  I0310077d53ae4ed9904df42e3f81c634['h03afe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d80] =  I0310077d53ae4ed9904df42e3f81c634['h03b00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d81] =  I0310077d53ae4ed9904df42e3f81c634['h03b02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d82] =  I0310077d53ae4ed9904df42e3f81c634['h03b04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d83] =  I0310077d53ae4ed9904df42e3f81c634['h03b06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d84] =  I0310077d53ae4ed9904df42e3f81c634['h03b08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d85] =  I0310077d53ae4ed9904df42e3f81c634['h03b0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d86] =  I0310077d53ae4ed9904df42e3f81c634['h03b0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d87] =  I0310077d53ae4ed9904df42e3f81c634['h03b0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d88] =  I0310077d53ae4ed9904df42e3f81c634['h03b10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d89] =  I0310077d53ae4ed9904df42e3f81c634['h03b12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d8a] =  I0310077d53ae4ed9904df42e3f81c634['h03b14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d8b] =  I0310077d53ae4ed9904df42e3f81c634['h03b16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d8c] =  I0310077d53ae4ed9904df42e3f81c634['h03b18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d8d] =  I0310077d53ae4ed9904df42e3f81c634['h03b1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d8e] =  I0310077d53ae4ed9904df42e3f81c634['h03b1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d8f] =  I0310077d53ae4ed9904df42e3f81c634['h03b1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d90] =  I0310077d53ae4ed9904df42e3f81c634['h03b20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d91] =  I0310077d53ae4ed9904df42e3f81c634['h03b22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d92] =  I0310077d53ae4ed9904df42e3f81c634['h03b24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d93] =  I0310077d53ae4ed9904df42e3f81c634['h03b26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d94] =  I0310077d53ae4ed9904df42e3f81c634['h03b28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d95] =  I0310077d53ae4ed9904df42e3f81c634['h03b2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d96] =  I0310077d53ae4ed9904df42e3f81c634['h03b2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d97] =  I0310077d53ae4ed9904df42e3f81c634['h03b2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d98] =  I0310077d53ae4ed9904df42e3f81c634['h03b30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d99] =  I0310077d53ae4ed9904df42e3f81c634['h03b32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d9a] =  I0310077d53ae4ed9904df42e3f81c634['h03b34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d9b] =  I0310077d53ae4ed9904df42e3f81c634['h03b36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d9c] =  I0310077d53ae4ed9904df42e3f81c634['h03b38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d9d] =  I0310077d53ae4ed9904df42e3f81c634['h03b3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d9e] =  I0310077d53ae4ed9904df42e3f81c634['h03b3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01d9f] =  I0310077d53ae4ed9904df42e3f81c634['h03b3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da0] =  I0310077d53ae4ed9904df42e3f81c634['h03b40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da1] =  I0310077d53ae4ed9904df42e3f81c634['h03b42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da2] =  I0310077d53ae4ed9904df42e3f81c634['h03b44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da3] =  I0310077d53ae4ed9904df42e3f81c634['h03b46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da4] =  I0310077d53ae4ed9904df42e3f81c634['h03b48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da5] =  I0310077d53ae4ed9904df42e3f81c634['h03b4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da6] =  I0310077d53ae4ed9904df42e3f81c634['h03b4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da7] =  I0310077d53ae4ed9904df42e3f81c634['h03b4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da8] =  I0310077d53ae4ed9904df42e3f81c634['h03b50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01da9] =  I0310077d53ae4ed9904df42e3f81c634['h03b52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01daa] =  I0310077d53ae4ed9904df42e3f81c634['h03b54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dab] =  I0310077d53ae4ed9904df42e3f81c634['h03b56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dac] =  I0310077d53ae4ed9904df42e3f81c634['h03b58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dad] =  I0310077d53ae4ed9904df42e3f81c634['h03b5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dae] =  I0310077d53ae4ed9904df42e3f81c634['h03b5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01daf] =  I0310077d53ae4ed9904df42e3f81c634['h03b5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db0] =  I0310077d53ae4ed9904df42e3f81c634['h03b60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db1] =  I0310077d53ae4ed9904df42e3f81c634['h03b62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db2] =  I0310077d53ae4ed9904df42e3f81c634['h03b64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db3] =  I0310077d53ae4ed9904df42e3f81c634['h03b66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db4] =  I0310077d53ae4ed9904df42e3f81c634['h03b68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db5] =  I0310077d53ae4ed9904df42e3f81c634['h03b6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db6] =  I0310077d53ae4ed9904df42e3f81c634['h03b6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db7] =  I0310077d53ae4ed9904df42e3f81c634['h03b6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db8] =  I0310077d53ae4ed9904df42e3f81c634['h03b70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01db9] =  I0310077d53ae4ed9904df42e3f81c634['h03b72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dba] =  I0310077d53ae4ed9904df42e3f81c634['h03b74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dbb] =  I0310077d53ae4ed9904df42e3f81c634['h03b76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dbc] =  I0310077d53ae4ed9904df42e3f81c634['h03b78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dbd] =  I0310077d53ae4ed9904df42e3f81c634['h03b7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dbe] =  I0310077d53ae4ed9904df42e3f81c634['h03b7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dbf] =  I0310077d53ae4ed9904df42e3f81c634['h03b7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc0] =  I0310077d53ae4ed9904df42e3f81c634['h03b80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc1] =  I0310077d53ae4ed9904df42e3f81c634['h03b82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc2] =  I0310077d53ae4ed9904df42e3f81c634['h03b84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc3] =  I0310077d53ae4ed9904df42e3f81c634['h03b86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc4] =  I0310077d53ae4ed9904df42e3f81c634['h03b88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc5] =  I0310077d53ae4ed9904df42e3f81c634['h03b8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc6] =  I0310077d53ae4ed9904df42e3f81c634['h03b8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc7] =  I0310077d53ae4ed9904df42e3f81c634['h03b8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc8] =  I0310077d53ae4ed9904df42e3f81c634['h03b90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dc9] =  I0310077d53ae4ed9904df42e3f81c634['h03b92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dca] =  I0310077d53ae4ed9904df42e3f81c634['h03b94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dcb] =  I0310077d53ae4ed9904df42e3f81c634['h03b96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dcc] =  I0310077d53ae4ed9904df42e3f81c634['h03b98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dcd] =  I0310077d53ae4ed9904df42e3f81c634['h03b9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dce] =  I0310077d53ae4ed9904df42e3f81c634['h03b9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dcf] =  I0310077d53ae4ed9904df42e3f81c634['h03b9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd0] =  I0310077d53ae4ed9904df42e3f81c634['h03ba0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd1] =  I0310077d53ae4ed9904df42e3f81c634['h03ba2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd2] =  I0310077d53ae4ed9904df42e3f81c634['h03ba4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd3] =  I0310077d53ae4ed9904df42e3f81c634['h03ba6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd4] =  I0310077d53ae4ed9904df42e3f81c634['h03ba8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd5] =  I0310077d53ae4ed9904df42e3f81c634['h03baa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd6] =  I0310077d53ae4ed9904df42e3f81c634['h03bac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd7] =  I0310077d53ae4ed9904df42e3f81c634['h03bae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd8] =  I0310077d53ae4ed9904df42e3f81c634['h03bb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dd9] =  I0310077d53ae4ed9904df42e3f81c634['h03bb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dda] =  I0310077d53ae4ed9904df42e3f81c634['h03bb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ddb] =  I0310077d53ae4ed9904df42e3f81c634['h03bb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ddc] =  I0310077d53ae4ed9904df42e3f81c634['h03bb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ddd] =  I0310077d53ae4ed9904df42e3f81c634['h03bba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dde] =  I0310077d53ae4ed9904df42e3f81c634['h03bbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ddf] =  I0310077d53ae4ed9904df42e3f81c634['h03bbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de0] =  I0310077d53ae4ed9904df42e3f81c634['h03bc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de1] =  I0310077d53ae4ed9904df42e3f81c634['h03bc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de2] =  I0310077d53ae4ed9904df42e3f81c634['h03bc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de3] =  I0310077d53ae4ed9904df42e3f81c634['h03bc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de4] =  I0310077d53ae4ed9904df42e3f81c634['h03bc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de5] =  I0310077d53ae4ed9904df42e3f81c634['h03bca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de6] =  I0310077d53ae4ed9904df42e3f81c634['h03bcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de7] =  I0310077d53ae4ed9904df42e3f81c634['h03bce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de8] =  I0310077d53ae4ed9904df42e3f81c634['h03bd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01de9] =  I0310077d53ae4ed9904df42e3f81c634['h03bd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dea] =  I0310077d53ae4ed9904df42e3f81c634['h03bd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01deb] =  I0310077d53ae4ed9904df42e3f81c634['h03bd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dec] =  I0310077d53ae4ed9904df42e3f81c634['h03bd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ded] =  I0310077d53ae4ed9904df42e3f81c634['h03bda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dee] =  I0310077d53ae4ed9904df42e3f81c634['h03bdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01def] =  I0310077d53ae4ed9904df42e3f81c634['h03bde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df0] =  I0310077d53ae4ed9904df42e3f81c634['h03be0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df1] =  I0310077d53ae4ed9904df42e3f81c634['h03be2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df2] =  I0310077d53ae4ed9904df42e3f81c634['h03be4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df3] =  I0310077d53ae4ed9904df42e3f81c634['h03be6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df4] =  I0310077d53ae4ed9904df42e3f81c634['h03be8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df5] =  I0310077d53ae4ed9904df42e3f81c634['h03bea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df6] =  I0310077d53ae4ed9904df42e3f81c634['h03bec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df7] =  I0310077d53ae4ed9904df42e3f81c634['h03bee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df8] =  I0310077d53ae4ed9904df42e3f81c634['h03bf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01df9] =  I0310077d53ae4ed9904df42e3f81c634['h03bf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dfa] =  I0310077d53ae4ed9904df42e3f81c634['h03bf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dfb] =  I0310077d53ae4ed9904df42e3f81c634['h03bf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dfc] =  I0310077d53ae4ed9904df42e3f81c634['h03bf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dfd] =  I0310077d53ae4ed9904df42e3f81c634['h03bfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dfe] =  I0310077d53ae4ed9904df42e3f81c634['h03bfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01dff] =  I0310077d53ae4ed9904df42e3f81c634['h03bfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e00] =  I0310077d53ae4ed9904df42e3f81c634['h03c00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e01] =  I0310077d53ae4ed9904df42e3f81c634['h03c02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e02] =  I0310077d53ae4ed9904df42e3f81c634['h03c04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e03] =  I0310077d53ae4ed9904df42e3f81c634['h03c06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e04] =  I0310077d53ae4ed9904df42e3f81c634['h03c08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e05] =  I0310077d53ae4ed9904df42e3f81c634['h03c0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e06] =  I0310077d53ae4ed9904df42e3f81c634['h03c0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e07] =  I0310077d53ae4ed9904df42e3f81c634['h03c0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e08] =  I0310077d53ae4ed9904df42e3f81c634['h03c10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e09] =  I0310077d53ae4ed9904df42e3f81c634['h03c12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e0a] =  I0310077d53ae4ed9904df42e3f81c634['h03c14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e0b] =  I0310077d53ae4ed9904df42e3f81c634['h03c16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e0c] =  I0310077d53ae4ed9904df42e3f81c634['h03c18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e0d] =  I0310077d53ae4ed9904df42e3f81c634['h03c1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e0e] =  I0310077d53ae4ed9904df42e3f81c634['h03c1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e0f] =  I0310077d53ae4ed9904df42e3f81c634['h03c1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e10] =  I0310077d53ae4ed9904df42e3f81c634['h03c20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e11] =  I0310077d53ae4ed9904df42e3f81c634['h03c22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e12] =  I0310077d53ae4ed9904df42e3f81c634['h03c24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e13] =  I0310077d53ae4ed9904df42e3f81c634['h03c26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e14] =  I0310077d53ae4ed9904df42e3f81c634['h03c28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e15] =  I0310077d53ae4ed9904df42e3f81c634['h03c2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e16] =  I0310077d53ae4ed9904df42e3f81c634['h03c2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e17] =  I0310077d53ae4ed9904df42e3f81c634['h03c2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e18] =  I0310077d53ae4ed9904df42e3f81c634['h03c30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e19] =  I0310077d53ae4ed9904df42e3f81c634['h03c32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e1a] =  I0310077d53ae4ed9904df42e3f81c634['h03c34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e1b] =  I0310077d53ae4ed9904df42e3f81c634['h03c36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e1c] =  I0310077d53ae4ed9904df42e3f81c634['h03c38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e1d] =  I0310077d53ae4ed9904df42e3f81c634['h03c3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e1e] =  I0310077d53ae4ed9904df42e3f81c634['h03c3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e1f] =  I0310077d53ae4ed9904df42e3f81c634['h03c3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e20] =  I0310077d53ae4ed9904df42e3f81c634['h03c40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e21] =  I0310077d53ae4ed9904df42e3f81c634['h03c42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e22] =  I0310077d53ae4ed9904df42e3f81c634['h03c44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e23] =  I0310077d53ae4ed9904df42e3f81c634['h03c46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e24] =  I0310077d53ae4ed9904df42e3f81c634['h03c48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e25] =  I0310077d53ae4ed9904df42e3f81c634['h03c4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e26] =  I0310077d53ae4ed9904df42e3f81c634['h03c4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e27] =  I0310077d53ae4ed9904df42e3f81c634['h03c4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e28] =  I0310077d53ae4ed9904df42e3f81c634['h03c50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e29] =  I0310077d53ae4ed9904df42e3f81c634['h03c52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e2a] =  I0310077d53ae4ed9904df42e3f81c634['h03c54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e2b] =  I0310077d53ae4ed9904df42e3f81c634['h03c56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e2c] =  I0310077d53ae4ed9904df42e3f81c634['h03c58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e2d] =  I0310077d53ae4ed9904df42e3f81c634['h03c5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e2e] =  I0310077d53ae4ed9904df42e3f81c634['h03c5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e2f] =  I0310077d53ae4ed9904df42e3f81c634['h03c5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e30] =  I0310077d53ae4ed9904df42e3f81c634['h03c60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e31] =  I0310077d53ae4ed9904df42e3f81c634['h03c62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e32] =  I0310077d53ae4ed9904df42e3f81c634['h03c64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e33] =  I0310077d53ae4ed9904df42e3f81c634['h03c66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e34] =  I0310077d53ae4ed9904df42e3f81c634['h03c68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e35] =  I0310077d53ae4ed9904df42e3f81c634['h03c6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e36] =  I0310077d53ae4ed9904df42e3f81c634['h03c6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e37] =  I0310077d53ae4ed9904df42e3f81c634['h03c6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e38] =  I0310077d53ae4ed9904df42e3f81c634['h03c70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e39] =  I0310077d53ae4ed9904df42e3f81c634['h03c72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e3a] =  I0310077d53ae4ed9904df42e3f81c634['h03c74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e3b] =  I0310077d53ae4ed9904df42e3f81c634['h03c76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e3c] =  I0310077d53ae4ed9904df42e3f81c634['h03c78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e3d] =  I0310077d53ae4ed9904df42e3f81c634['h03c7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e3e] =  I0310077d53ae4ed9904df42e3f81c634['h03c7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e3f] =  I0310077d53ae4ed9904df42e3f81c634['h03c7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e40] =  I0310077d53ae4ed9904df42e3f81c634['h03c80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e41] =  I0310077d53ae4ed9904df42e3f81c634['h03c82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e42] =  I0310077d53ae4ed9904df42e3f81c634['h03c84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e43] =  I0310077d53ae4ed9904df42e3f81c634['h03c86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e44] =  I0310077d53ae4ed9904df42e3f81c634['h03c88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e45] =  I0310077d53ae4ed9904df42e3f81c634['h03c8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e46] =  I0310077d53ae4ed9904df42e3f81c634['h03c8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e47] =  I0310077d53ae4ed9904df42e3f81c634['h03c8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e48] =  I0310077d53ae4ed9904df42e3f81c634['h03c90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e49] =  I0310077d53ae4ed9904df42e3f81c634['h03c92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e4a] =  I0310077d53ae4ed9904df42e3f81c634['h03c94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e4b] =  I0310077d53ae4ed9904df42e3f81c634['h03c96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e4c] =  I0310077d53ae4ed9904df42e3f81c634['h03c98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e4d] =  I0310077d53ae4ed9904df42e3f81c634['h03c9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e4e] =  I0310077d53ae4ed9904df42e3f81c634['h03c9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e4f] =  I0310077d53ae4ed9904df42e3f81c634['h03c9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e50] =  I0310077d53ae4ed9904df42e3f81c634['h03ca0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e51] =  I0310077d53ae4ed9904df42e3f81c634['h03ca2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e52] =  I0310077d53ae4ed9904df42e3f81c634['h03ca4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e53] =  I0310077d53ae4ed9904df42e3f81c634['h03ca6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e54] =  I0310077d53ae4ed9904df42e3f81c634['h03ca8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e55] =  I0310077d53ae4ed9904df42e3f81c634['h03caa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e56] =  I0310077d53ae4ed9904df42e3f81c634['h03cac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e57] =  I0310077d53ae4ed9904df42e3f81c634['h03cae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e58] =  I0310077d53ae4ed9904df42e3f81c634['h03cb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e59] =  I0310077d53ae4ed9904df42e3f81c634['h03cb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e5a] =  I0310077d53ae4ed9904df42e3f81c634['h03cb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e5b] =  I0310077d53ae4ed9904df42e3f81c634['h03cb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e5c] =  I0310077d53ae4ed9904df42e3f81c634['h03cb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e5d] =  I0310077d53ae4ed9904df42e3f81c634['h03cba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e5e] =  I0310077d53ae4ed9904df42e3f81c634['h03cbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e5f] =  I0310077d53ae4ed9904df42e3f81c634['h03cbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e60] =  I0310077d53ae4ed9904df42e3f81c634['h03cc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e61] =  I0310077d53ae4ed9904df42e3f81c634['h03cc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e62] =  I0310077d53ae4ed9904df42e3f81c634['h03cc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e63] =  I0310077d53ae4ed9904df42e3f81c634['h03cc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e64] =  I0310077d53ae4ed9904df42e3f81c634['h03cc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e65] =  I0310077d53ae4ed9904df42e3f81c634['h03cca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e66] =  I0310077d53ae4ed9904df42e3f81c634['h03ccc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e67] =  I0310077d53ae4ed9904df42e3f81c634['h03cce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e68] =  I0310077d53ae4ed9904df42e3f81c634['h03cd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e69] =  I0310077d53ae4ed9904df42e3f81c634['h03cd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e6a] =  I0310077d53ae4ed9904df42e3f81c634['h03cd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e6b] =  I0310077d53ae4ed9904df42e3f81c634['h03cd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e6c] =  I0310077d53ae4ed9904df42e3f81c634['h03cd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e6d] =  I0310077d53ae4ed9904df42e3f81c634['h03cda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e6e] =  I0310077d53ae4ed9904df42e3f81c634['h03cdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e6f] =  I0310077d53ae4ed9904df42e3f81c634['h03cde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e70] =  I0310077d53ae4ed9904df42e3f81c634['h03ce0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e71] =  I0310077d53ae4ed9904df42e3f81c634['h03ce2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e72] =  I0310077d53ae4ed9904df42e3f81c634['h03ce4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e73] =  I0310077d53ae4ed9904df42e3f81c634['h03ce6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e74] =  I0310077d53ae4ed9904df42e3f81c634['h03ce8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e75] =  I0310077d53ae4ed9904df42e3f81c634['h03cea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e76] =  I0310077d53ae4ed9904df42e3f81c634['h03cec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e77] =  I0310077d53ae4ed9904df42e3f81c634['h03cee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e78] =  I0310077d53ae4ed9904df42e3f81c634['h03cf0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e79] =  I0310077d53ae4ed9904df42e3f81c634['h03cf2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e7a] =  I0310077d53ae4ed9904df42e3f81c634['h03cf4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e7b] =  I0310077d53ae4ed9904df42e3f81c634['h03cf6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e7c] =  I0310077d53ae4ed9904df42e3f81c634['h03cf8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e7d] =  I0310077d53ae4ed9904df42e3f81c634['h03cfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e7e] =  I0310077d53ae4ed9904df42e3f81c634['h03cfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e7f] =  I0310077d53ae4ed9904df42e3f81c634['h03cfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e80] =  I0310077d53ae4ed9904df42e3f81c634['h03d00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e81] =  I0310077d53ae4ed9904df42e3f81c634['h03d02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e82] =  I0310077d53ae4ed9904df42e3f81c634['h03d04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e83] =  I0310077d53ae4ed9904df42e3f81c634['h03d06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e84] =  I0310077d53ae4ed9904df42e3f81c634['h03d08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e85] =  I0310077d53ae4ed9904df42e3f81c634['h03d0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e86] =  I0310077d53ae4ed9904df42e3f81c634['h03d0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e87] =  I0310077d53ae4ed9904df42e3f81c634['h03d0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e88] =  I0310077d53ae4ed9904df42e3f81c634['h03d10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e89] =  I0310077d53ae4ed9904df42e3f81c634['h03d12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e8a] =  I0310077d53ae4ed9904df42e3f81c634['h03d14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e8b] =  I0310077d53ae4ed9904df42e3f81c634['h03d16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e8c] =  I0310077d53ae4ed9904df42e3f81c634['h03d18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e8d] =  I0310077d53ae4ed9904df42e3f81c634['h03d1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e8e] =  I0310077d53ae4ed9904df42e3f81c634['h03d1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e8f] =  I0310077d53ae4ed9904df42e3f81c634['h03d1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e90] =  I0310077d53ae4ed9904df42e3f81c634['h03d20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e91] =  I0310077d53ae4ed9904df42e3f81c634['h03d22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e92] =  I0310077d53ae4ed9904df42e3f81c634['h03d24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e93] =  I0310077d53ae4ed9904df42e3f81c634['h03d26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e94] =  I0310077d53ae4ed9904df42e3f81c634['h03d28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e95] =  I0310077d53ae4ed9904df42e3f81c634['h03d2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e96] =  I0310077d53ae4ed9904df42e3f81c634['h03d2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e97] =  I0310077d53ae4ed9904df42e3f81c634['h03d2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e98] =  I0310077d53ae4ed9904df42e3f81c634['h03d30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e99] =  I0310077d53ae4ed9904df42e3f81c634['h03d32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e9a] =  I0310077d53ae4ed9904df42e3f81c634['h03d34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e9b] =  I0310077d53ae4ed9904df42e3f81c634['h03d36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e9c] =  I0310077d53ae4ed9904df42e3f81c634['h03d38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e9d] =  I0310077d53ae4ed9904df42e3f81c634['h03d3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e9e] =  I0310077d53ae4ed9904df42e3f81c634['h03d3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01e9f] =  I0310077d53ae4ed9904df42e3f81c634['h03d3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea0] =  I0310077d53ae4ed9904df42e3f81c634['h03d40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea1] =  I0310077d53ae4ed9904df42e3f81c634['h03d42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea2] =  I0310077d53ae4ed9904df42e3f81c634['h03d44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea3] =  I0310077d53ae4ed9904df42e3f81c634['h03d46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea4] =  I0310077d53ae4ed9904df42e3f81c634['h03d48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea5] =  I0310077d53ae4ed9904df42e3f81c634['h03d4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea6] =  I0310077d53ae4ed9904df42e3f81c634['h03d4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea7] =  I0310077d53ae4ed9904df42e3f81c634['h03d4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea8] =  I0310077d53ae4ed9904df42e3f81c634['h03d50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ea9] =  I0310077d53ae4ed9904df42e3f81c634['h03d52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eaa] =  I0310077d53ae4ed9904df42e3f81c634['h03d54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eab] =  I0310077d53ae4ed9904df42e3f81c634['h03d56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eac] =  I0310077d53ae4ed9904df42e3f81c634['h03d58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ead] =  I0310077d53ae4ed9904df42e3f81c634['h03d5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eae] =  I0310077d53ae4ed9904df42e3f81c634['h03d5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eaf] =  I0310077d53ae4ed9904df42e3f81c634['h03d5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb0] =  I0310077d53ae4ed9904df42e3f81c634['h03d60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb1] =  I0310077d53ae4ed9904df42e3f81c634['h03d62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb2] =  I0310077d53ae4ed9904df42e3f81c634['h03d64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb3] =  I0310077d53ae4ed9904df42e3f81c634['h03d66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb4] =  I0310077d53ae4ed9904df42e3f81c634['h03d68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb5] =  I0310077d53ae4ed9904df42e3f81c634['h03d6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb6] =  I0310077d53ae4ed9904df42e3f81c634['h03d6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb7] =  I0310077d53ae4ed9904df42e3f81c634['h03d6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb8] =  I0310077d53ae4ed9904df42e3f81c634['h03d70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eb9] =  I0310077d53ae4ed9904df42e3f81c634['h03d72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eba] =  I0310077d53ae4ed9904df42e3f81c634['h03d74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ebb] =  I0310077d53ae4ed9904df42e3f81c634['h03d76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ebc] =  I0310077d53ae4ed9904df42e3f81c634['h03d78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ebd] =  I0310077d53ae4ed9904df42e3f81c634['h03d7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ebe] =  I0310077d53ae4ed9904df42e3f81c634['h03d7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ebf] =  I0310077d53ae4ed9904df42e3f81c634['h03d7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec0] =  I0310077d53ae4ed9904df42e3f81c634['h03d80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec1] =  I0310077d53ae4ed9904df42e3f81c634['h03d82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec2] =  I0310077d53ae4ed9904df42e3f81c634['h03d84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec3] =  I0310077d53ae4ed9904df42e3f81c634['h03d86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec4] =  I0310077d53ae4ed9904df42e3f81c634['h03d88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec5] =  I0310077d53ae4ed9904df42e3f81c634['h03d8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec6] =  I0310077d53ae4ed9904df42e3f81c634['h03d8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec7] =  I0310077d53ae4ed9904df42e3f81c634['h03d8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec8] =  I0310077d53ae4ed9904df42e3f81c634['h03d90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ec9] =  I0310077d53ae4ed9904df42e3f81c634['h03d92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eca] =  I0310077d53ae4ed9904df42e3f81c634['h03d94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ecb] =  I0310077d53ae4ed9904df42e3f81c634['h03d96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ecc] =  I0310077d53ae4ed9904df42e3f81c634['h03d98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ecd] =  I0310077d53ae4ed9904df42e3f81c634['h03d9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ece] =  I0310077d53ae4ed9904df42e3f81c634['h03d9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ecf] =  I0310077d53ae4ed9904df42e3f81c634['h03d9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed0] =  I0310077d53ae4ed9904df42e3f81c634['h03da0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed1] =  I0310077d53ae4ed9904df42e3f81c634['h03da2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed2] =  I0310077d53ae4ed9904df42e3f81c634['h03da4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed3] =  I0310077d53ae4ed9904df42e3f81c634['h03da6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed4] =  I0310077d53ae4ed9904df42e3f81c634['h03da8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed5] =  I0310077d53ae4ed9904df42e3f81c634['h03daa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed6] =  I0310077d53ae4ed9904df42e3f81c634['h03dac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed7] =  I0310077d53ae4ed9904df42e3f81c634['h03dae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed8] =  I0310077d53ae4ed9904df42e3f81c634['h03db0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ed9] =  I0310077d53ae4ed9904df42e3f81c634['h03db2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eda] =  I0310077d53ae4ed9904df42e3f81c634['h03db4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01edb] =  I0310077d53ae4ed9904df42e3f81c634['h03db6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01edc] =  I0310077d53ae4ed9904df42e3f81c634['h03db8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01edd] =  I0310077d53ae4ed9904df42e3f81c634['h03dba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ede] =  I0310077d53ae4ed9904df42e3f81c634['h03dbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01edf] =  I0310077d53ae4ed9904df42e3f81c634['h03dbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee0] =  I0310077d53ae4ed9904df42e3f81c634['h03dc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee1] =  I0310077d53ae4ed9904df42e3f81c634['h03dc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee2] =  I0310077d53ae4ed9904df42e3f81c634['h03dc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee3] =  I0310077d53ae4ed9904df42e3f81c634['h03dc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee4] =  I0310077d53ae4ed9904df42e3f81c634['h03dc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee5] =  I0310077d53ae4ed9904df42e3f81c634['h03dca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee6] =  I0310077d53ae4ed9904df42e3f81c634['h03dcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee7] =  I0310077d53ae4ed9904df42e3f81c634['h03dce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee8] =  I0310077d53ae4ed9904df42e3f81c634['h03dd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ee9] =  I0310077d53ae4ed9904df42e3f81c634['h03dd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eea] =  I0310077d53ae4ed9904df42e3f81c634['h03dd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eeb] =  I0310077d53ae4ed9904df42e3f81c634['h03dd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eec] =  I0310077d53ae4ed9904df42e3f81c634['h03dd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eed] =  I0310077d53ae4ed9904df42e3f81c634['h03dda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eee] =  I0310077d53ae4ed9904df42e3f81c634['h03ddc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eef] =  I0310077d53ae4ed9904df42e3f81c634['h03dde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef0] =  I0310077d53ae4ed9904df42e3f81c634['h03de0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef1] =  I0310077d53ae4ed9904df42e3f81c634['h03de2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef2] =  I0310077d53ae4ed9904df42e3f81c634['h03de4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef3] =  I0310077d53ae4ed9904df42e3f81c634['h03de6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef4] =  I0310077d53ae4ed9904df42e3f81c634['h03de8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef5] =  I0310077d53ae4ed9904df42e3f81c634['h03dea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef6] =  I0310077d53ae4ed9904df42e3f81c634['h03dec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef7] =  I0310077d53ae4ed9904df42e3f81c634['h03dee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef8] =  I0310077d53ae4ed9904df42e3f81c634['h03df0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ef9] =  I0310077d53ae4ed9904df42e3f81c634['h03df2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01efa] =  I0310077d53ae4ed9904df42e3f81c634['h03df4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01efb] =  I0310077d53ae4ed9904df42e3f81c634['h03df6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01efc] =  I0310077d53ae4ed9904df42e3f81c634['h03df8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01efd] =  I0310077d53ae4ed9904df42e3f81c634['h03dfa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01efe] =  I0310077d53ae4ed9904df42e3f81c634['h03dfc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01eff] =  I0310077d53ae4ed9904df42e3f81c634['h03dfe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f00] =  I0310077d53ae4ed9904df42e3f81c634['h03e00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f01] =  I0310077d53ae4ed9904df42e3f81c634['h03e02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f02] =  I0310077d53ae4ed9904df42e3f81c634['h03e04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f03] =  I0310077d53ae4ed9904df42e3f81c634['h03e06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f04] =  I0310077d53ae4ed9904df42e3f81c634['h03e08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f05] =  I0310077d53ae4ed9904df42e3f81c634['h03e0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f06] =  I0310077d53ae4ed9904df42e3f81c634['h03e0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f07] =  I0310077d53ae4ed9904df42e3f81c634['h03e0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f08] =  I0310077d53ae4ed9904df42e3f81c634['h03e10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f09] =  I0310077d53ae4ed9904df42e3f81c634['h03e12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f0a] =  I0310077d53ae4ed9904df42e3f81c634['h03e14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f0b] =  I0310077d53ae4ed9904df42e3f81c634['h03e16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f0c] =  I0310077d53ae4ed9904df42e3f81c634['h03e18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f0d] =  I0310077d53ae4ed9904df42e3f81c634['h03e1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f0e] =  I0310077d53ae4ed9904df42e3f81c634['h03e1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f0f] =  I0310077d53ae4ed9904df42e3f81c634['h03e1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f10] =  I0310077d53ae4ed9904df42e3f81c634['h03e20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f11] =  I0310077d53ae4ed9904df42e3f81c634['h03e22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f12] =  I0310077d53ae4ed9904df42e3f81c634['h03e24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f13] =  I0310077d53ae4ed9904df42e3f81c634['h03e26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f14] =  I0310077d53ae4ed9904df42e3f81c634['h03e28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f15] =  I0310077d53ae4ed9904df42e3f81c634['h03e2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f16] =  I0310077d53ae4ed9904df42e3f81c634['h03e2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f17] =  I0310077d53ae4ed9904df42e3f81c634['h03e2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f18] =  I0310077d53ae4ed9904df42e3f81c634['h03e30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f19] =  I0310077d53ae4ed9904df42e3f81c634['h03e32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f1a] =  I0310077d53ae4ed9904df42e3f81c634['h03e34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f1b] =  I0310077d53ae4ed9904df42e3f81c634['h03e36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f1c] =  I0310077d53ae4ed9904df42e3f81c634['h03e38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f1d] =  I0310077d53ae4ed9904df42e3f81c634['h03e3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f1e] =  I0310077d53ae4ed9904df42e3f81c634['h03e3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f1f] =  I0310077d53ae4ed9904df42e3f81c634['h03e3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f20] =  I0310077d53ae4ed9904df42e3f81c634['h03e40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f21] =  I0310077d53ae4ed9904df42e3f81c634['h03e42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f22] =  I0310077d53ae4ed9904df42e3f81c634['h03e44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f23] =  I0310077d53ae4ed9904df42e3f81c634['h03e46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f24] =  I0310077d53ae4ed9904df42e3f81c634['h03e48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f25] =  I0310077d53ae4ed9904df42e3f81c634['h03e4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f26] =  I0310077d53ae4ed9904df42e3f81c634['h03e4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f27] =  I0310077d53ae4ed9904df42e3f81c634['h03e4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f28] =  I0310077d53ae4ed9904df42e3f81c634['h03e50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f29] =  I0310077d53ae4ed9904df42e3f81c634['h03e52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f2a] =  I0310077d53ae4ed9904df42e3f81c634['h03e54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f2b] =  I0310077d53ae4ed9904df42e3f81c634['h03e56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f2c] =  I0310077d53ae4ed9904df42e3f81c634['h03e58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f2d] =  I0310077d53ae4ed9904df42e3f81c634['h03e5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f2e] =  I0310077d53ae4ed9904df42e3f81c634['h03e5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f2f] =  I0310077d53ae4ed9904df42e3f81c634['h03e5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f30] =  I0310077d53ae4ed9904df42e3f81c634['h03e60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f31] =  I0310077d53ae4ed9904df42e3f81c634['h03e62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f32] =  I0310077d53ae4ed9904df42e3f81c634['h03e64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f33] =  I0310077d53ae4ed9904df42e3f81c634['h03e66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f34] =  I0310077d53ae4ed9904df42e3f81c634['h03e68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f35] =  I0310077d53ae4ed9904df42e3f81c634['h03e6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f36] =  I0310077d53ae4ed9904df42e3f81c634['h03e6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f37] =  I0310077d53ae4ed9904df42e3f81c634['h03e6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f38] =  I0310077d53ae4ed9904df42e3f81c634['h03e70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f39] =  I0310077d53ae4ed9904df42e3f81c634['h03e72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f3a] =  I0310077d53ae4ed9904df42e3f81c634['h03e74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f3b] =  I0310077d53ae4ed9904df42e3f81c634['h03e76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f3c] =  I0310077d53ae4ed9904df42e3f81c634['h03e78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f3d] =  I0310077d53ae4ed9904df42e3f81c634['h03e7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f3e] =  I0310077d53ae4ed9904df42e3f81c634['h03e7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f3f] =  I0310077d53ae4ed9904df42e3f81c634['h03e7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f40] =  I0310077d53ae4ed9904df42e3f81c634['h03e80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f41] =  I0310077d53ae4ed9904df42e3f81c634['h03e82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f42] =  I0310077d53ae4ed9904df42e3f81c634['h03e84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f43] =  I0310077d53ae4ed9904df42e3f81c634['h03e86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f44] =  I0310077d53ae4ed9904df42e3f81c634['h03e88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f45] =  I0310077d53ae4ed9904df42e3f81c634['h03e8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f46] =  I0310077d53ae4ed9904df42e3f81c634['h03e8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f47] =  I0310077d53ae4ed9904df42e3f81c634['h03e8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f48] =  I0310077d53ae4ed9904df42e3f81c634['h03e90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f49] =  I0310077d53ae4ed9904df42e3f81c634['h03e92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f4a] =  I0310077d53ae4ed9904df42e3f81c634['h03e94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f4b] =  I0310077d53ae4ed9904df42e3f81c634['h03e96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f4c] =  I0310077d53ae4ed9904df42e3f81c634['h03e98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f4d] =  I0310077d53ae4ed9904df42e3f81c634['h03e9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f4e] =  I0310077d53ae4ed9904df42e3f81c634['h03e9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f4f] =  I0310077d53ae4ed9904df42e3f81c634['h03e9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f50] =  I0310077d53ae4ed9904df42e3f81c634['h03ea0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f51] =  I0310077d53ae4ed9904df42e3f81c634['h03ea2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f52] =  I0310077d53ae4ed9904df42e3f81c634['h03ea4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f53] =  I0310077d53ae4ed9904df42e3f81c634['h03ea6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f54] =  I0310077d53ae4ed9904df42e3f81c634['h03ea8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f55] =  I0310077d53ae4ed9904df42e3f81c634['h03eaa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f56] =  I0310077d53ae4ed9904df42e3f81c634['h03eac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f57] =  I0310077d53ae4ed9904df42e3f81c634['h03eae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f58] =  I0310077d53ae4ed9904df42e3f81c634['h03eb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f59] =  I0310077d53ae4ed9904df42e3f81c634['h03eb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f5a] =  I0310077d53ae4ed9904df42e3f81c634['h03eb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f5b] =  I0310077d53ae4ed9904df42e3f81c634['h03eb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f5c] =  I0310077d53ae4ed9904df42e3f81c634['h03eb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f5d] =  I0310077d53ae4ed9904df42e3f81c634['h03eba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f5e] =  I0310077d53ae4ed9904df42e3f81c634['h03ebc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f5f] =  I0310077d53ae4ed9904df42e3f81c634['h03ebe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f60] =  I0310077d53ae4ed9904df42e3f81c634['h03ec0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f61] =  I0310077d53ae4ed9904df42e3f81c634['h03ec2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f62] =  I0310077d53ae4ed9904df42e3f81c634['h03ec4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f63] =  I0310077d53ae4ed9904df42e3f81c634['h03ec6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f64] =  I0310077d53ae4ed9904df42e3f81c634['h03ec8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f65] =  I0310077d53ae4ed9904df42e3f81c634['h03eca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f66] =  I0310077d53ae4ed9904df42e3f81c634['h03ecc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f67] =  I0310077d53ae4ed9904df42e3f81c634['h03ece] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f68] =  I0310077d53ae4ed9904df42e3f81c634['h03ed0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f69] =  I0310077d53ae4ed9904df42e3f81c634['h03ed2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f6a] =  I0310077d53ae4ed9904df42e3f81c634['h03ed4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f6b] =  I0310077d53ae4ed9904df42e3f81c634['h03ed6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f6c] =  I0310077d53ae4ed9904df42e3f81c634['h03ed8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f6d] =  I0310077d53ae4ed9904df42e3f81c634['h03eda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f6e] =  I0310077d53ae4ed9904df42e3f81c634['h03edc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f6f] =  I0310077d53ae4ed9904df42e3f81c634['h03ede] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f70] =  I0310077d53ae4ed9904df42e3f81c634['h03ee0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f71] =  I0310077d53ae4ed9904df42e3f81c634['h03ee2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f72] =  I0310077d53ae4ed9904df42e3f81c634['h03ee4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f73] =  I0310077d53ae4ed9904df42e3f81c634['h03ee6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f74] =  I0310077d53ae4ed9904df42e3f81c634['h03ee8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f75] =  I0310077d53ae4ed9904df42e3f81c634['h03eea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f76] =  I0310077d53ae4ed9904df42e3f81c634['h03eec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f77] =  I0310077d53ae4ed9904df42e3f81c634['h03eee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f78] =  I0310077d53ae4ed9904df42e3f81c634['h03ef0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f79] =  I0310077d53ae4ed9904df42e3f81c634['h03ef2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f7a] =  I0310077d53ae4ed9904df42e3f81c634['h03ef4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f7b] =  I0310077d53ae4ed9904df42e3f81c634['h03ef6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f7c] =  I0310077d53ae4ed9904df42e3f81c634['h03ef8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f7d] =  I0310077d53ae4ed9904df42e3f81c634['h03efa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f7e] =  I0310077d53ae4ed9904df42e3f81c634['h03efc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f7f] =  I0310077d53ae4ed9904df42e3f81c634['h03efe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f80] =  I0310077d53ae4ed9904df42e3f81c634['h03f00] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f81] =  I0310077d53ae4ed9904df42e3f81c634['h03f02] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f82] =  I0310077d53ae4ed9904df42e3f81c634['h03f04] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f83] =  I0310077d53ae4ed9904df42e3f81c634['h03f06] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f84] =  I0310077d53ae4ed9904df42e3f81c634['h03f08] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f85] =  I0310077d53ae4ed9904df42e3f81c634['h03f0a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f86] =  I0310077d53ae4ed9904df42e3f81c634['h03f0c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f87] =  I0310077d53ae4ed9904df42e3f81c634['h03f0e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f88] =  I0310077d53ae4ed9904df42e3f81c634['h03f10] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f89] =  I0310077d53ae4ed9904df42e3f81c634['h03f12] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f8a] =  I0310077d53ae4ed9904df42e3f81c634['h03f14] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f8b] =  I0310077d53ae4ed9904df42e3f81c634['h03f16] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f8c] =  I0310077d53ae4ed9904df42e3f81c634['h03f18] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f8d] =  I0310077d53ae4ed9904df42e3f81c634['h03f1a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f8e] =  I0310077d53ae4ed9904df42e3f81c634['h03f1c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f8f] =  I0310077d53ae4ed9904df42e3f81c634['h03f1e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f90] =  I0310077d53ae4ed9904df42e3f81c634['h03f20] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f91] =  I0310077d53ae4ed9904df42e3f81c634['h03f22] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f92] =  I0310077d53ae4ed9904df42e3f81c634['h03f24] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f93] =  I0310077d53ae4ed9904df42e3f81c634['h03f26] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f94] =  I0310077d53ae4ed9904df42e3f81c634['h03f28] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f95] =  I0310077d53ae4ed9904df42e3f81c634['h03f2a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f96] =  I0310077d53ae4ed9904df42e3f81c634['h03f2c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f97] =  I0310077d53ae4ed9904df42e3f81c634['h03f2e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f98] =  I0310077d53ae4ed9904df42e3f81c634['h03f30] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f99] =  I0310077d53ae4ed9904df42e3f81c634['h03f32] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f9a] =  I0310077d53ae4ed9904df42e3f81c634['h03f34] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f9b] =  I0310077d53ae4ed9904df42e3f81c634['h03f36] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f9c] =  I0310077d53ae4ed9904df42e3f81c634['h03f38] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f9d] =  I0310077d53ae4ed9904df42e3f81c634['h03f3a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f9e] =  I0310077d53ae4ed9904df42e3f81c634['h03f3c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01f9f] =  I0310077d53ae4ed9904df42e3f81c634['h03f3e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa0] =  I0310077d53ae4ed9904df42e3f81c634['h03f40] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa1] =  I0310077d53ae4ed9904df42e3f81c634['h03f42] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa2] =  I0310077d53ae4ed9904df42e3f81c634['h03f44] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa3] =  I0310077d53ae4ed9904df42e3f81c634['h03f46] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa4] =  I0310077d53ae4ed9904df42e3f81c634['h03f48] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa5] =  I0310077d53ae4ed9904df42e3f81c634['h03f4a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa6] =  I0310077d53ae4ed9904df42e3f81c634['h03f4c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa7] =  I0310077d53ae4ed9904df42e3f81c634['h03f4e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa8] =  I0310077d53ae4ed9904df42e3f81c634['h03f50] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fa9] =  I0310077d53ae4ed9904df42e3f81c634['h03f52] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01faa] =  I0310077d53ae4ed9904df42e3f81c634['h03f54] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fab] =  I0310077d53ae4ed9904df42e3f81c634['h03f56] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fac] =  I0310077d53ae4ed9904df42e3f81c634['h03f58] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fad] =  I0310077d53ae4ed9904df42e3f81c634['h03f5a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fae] =  I0310077d53ae4ed9904df42e3f81c634['h03f5c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01faf] =  I0310077d53ae4ed9904df42e3f81c634['h03f5e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb0] =  I0310077d53ae4ed9904df42e3f81c634['h03f60] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb1] =  I0310077d53ae4ed9904df42e3f81c634['h03f62] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb2] =  I0310077d53ae4ed9904df42e3f81c634['h03f64] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb3] =  I0310077d53ae4ed9904df42e3f81c634['h03f66] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb4] =  I0310077d53ae4ed9904df42e3f81c634['h03f68] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb5] =  I0310077d53ae4ed9904df42e3f81c634['h03f6a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb6] =  I0310077d53ae4ed9904df42e3f81c634['h03f6c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb7] =  I0310077d53ae4ed9904df42e3f81c634['h03f6e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb8] =  I0310077d53ae4ed9904df42e3f81c634['h03f70] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fb9] =  I0310077d53ae4ed9904df42e3f81c634['h03f72] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fba] =  I0310077d53ae4ed9904df42e3f81c634['h03f74] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fbb] =  I0310077d53ae4ed9904df42e3f81c634['h03f76] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fbc] =  I0310077d53ae4ed9904df42e3f81c634['h03f78] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fbd] =  I0310077d53ae4ed9904df42e3f81c634['h03f7a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fbe] =  I0310077d53ae4ed9904df42e3f81c634['h03f7c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fbf] =  I0310077d53ae4ed9904df42e3f81c634['h03f7e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc0] =  I0310077d53ae4ed9904df42e3f81c634['h03f80] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc1] =  I0310077d53ae4ed9904df42e3f81c634['h03f82] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc2] =  I0310077d53ae4ed9904df42e3f81c634['h03f84] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc3] =  I0310077d53ae4ed9904df42e3f81c634['h03f86] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc4] =  I0310077d53ae4ed9904df42e3f81c634['h03f88] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc5] =  I0310077d53ae4ed9904df42e3f81c634['h03f8a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc6] =  I0310077d53ae4ed9904df42e3f81c634['h03f8c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc7] =  I0310077d53ae4ed9904df42e3f81c634['h03f8e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc8] =  I0310077d53ae4ed9904df42e3f81c634['h03f90] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fc9] =  I0310077d53ae4ed9904df42e3f81c634['h03f92] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fca] =  I0310077d53ae4ed9904df42e3f81c634['h03f94] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fcb] =  I0310077d53ae4ed9904df42e3f81c634['h03f96] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fcc] =  I0310077d53ae4ed9904df42e3f81c634['h03f98] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fcd] =  I0310077d53ae4ed9904df42e3f81c634['h03f9a] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fce] =  I0310077d53ae4ed9904df42e3f81c634['h03f9c] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fcf] =  I0310077d53ae4ed9904df42e3f81c634['h03f9e] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd0] =  I0310077d53ae4ed9904df42e3f81c634['h03fa0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd1] =  I0310077d53ae4ed9904df42e3f81c634['h03fa2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd2] =  I0310077d53ae4ed9904df42e3f81c634['h03fa4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd3] =  I0310077d53ae4ed9904df42e3f81c634['h03fa6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd4] =  I0310077d53ae4ed9904df42e3f81c634['h03fa8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd5] =  I0310077d53ae4ed9904df42e3f81c634['h03faa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd6] =  I0310077d53ae4ed9904df42e3f81c634['h03fac] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd7] =  I0310077d53ae4ed9904df42e3f81c634['h03fae] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd8] =  I0310077d53ae4ed9904df42e3f81c634['h03fb0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fd9] =  I0310077d53ae4ed9904df42e3f81c634['h03fb2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fda] =  I0310077d53ae4ed9904df42e3f81c634['h03fb4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fdb] =  I0310077d53ae4ed9904df42e3f81c634['h03fb6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fdc] =  I0310077d53ae4ed9904df42e3f81c634['h03fb8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fdd] =  I0310077d53ae4ed9904df42e3f81c634['h03fba] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fde] =  I0310077d53ae4ed9904df42e3f81c634['h03fbc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fdf] =  I0310077d53ae4ed9904df42e3f81c634['h03fbe] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe0] =  I0310077d53ae4ed9904df42e3f81c634['h03fc0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe1] =  I0310077d53ae4ed9904df42e3f81c634['h03fc2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe2] =  I0310077d53ae4ed9904df42e3f81c634['h03fc4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe3] =  I0310077d53ae4ed9904df42e3f81c634['h03fc6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe4] =  I0310077d53ae4ed9904df42e3f81c634['h03fc8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe5] =  I0310077d53ae4ed9904df42e3f81c634['h03fca] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe6] =  I0310077d53ae4ed9904df42e3f81c634['h03fcc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe7] =  I0310077d53ae4ed9904df42e3f81c634['h03fce] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe8] =  I0310077d53ae4ed9904df42e3f81c634['h03fd0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fe9] =  I0310077d53ae4ed9904df42e3f81c634['h03fd2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fea] =  I0310077d53ae4ed9904df42e3f81c634['h03fd4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01feb] =  I0310077d53ae4ed9904df42e3f81c634['h03fd6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fec] =  I0310077d53ae4ed9904df42e3f81c634['h03fd8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fed] =  I0310077d53ae4ed9904df42e3f81c634['h03fda] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fee] =  I0310077d53ae4ed9904df42e3f81c634['h03fdc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fef] =  I0310077d53ae4ed9904df42e3f81c634['h03fde] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff0] =  I0310077d53ae4ed9904df42e3f81c634['h03fe0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff1] =  I0310077d53ae4ed9904df42e3f81c634['h03fe2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff2] =  I0310077d53ae4ed9904df42e3f81c634['h03fe4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff3] =  I0310077d53ae4ed9904df42e3f81c634['h03fe6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff4] =  I0310077d53ae4ed9904df42e3f81c634['h03fe8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff5] =  I0310077d53ae4ed9904df42e3f81c634['h03fea] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff6] =  I0310077d53ae4ed9904df42e3f81c634['h03fec] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff7] =  I0310077d53ae4ed9904df42e3f81c634['h03fee] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff8] =  I0310077d53ae4ed9904df42e3f81c634['h03ff0] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ff9] =  I0310077d53ae4ed9904df42e3f81c634['h03ff2] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ffa] =  I0310077d53ae4ed9904df42e3f81c634['h03ff4] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ffb] =  I0310077d53ae4ed9904df42e3f81c634['h03ff6] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ffc] =  I0310077d53ae4ed9904df42e3f81c634['h03ff8] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ffd] =  I0310077d53ae4ed9904df42e3f81c634['h03ffa] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01ffe] =  I0310077d53ae4ed9904df42e3f81c634['h03ffc] ;
//end
//always_comb begin // 
               Ifcca41d795dde8a35d1654b9520c92e7['h01fff] =  I0310077d53ae4ed9904df42e3f81c634['h03ffe] ;
//end
