parameter flogtanh_WDTH = 10 ,
parameter flogtanh_MAX = 'h380 ,
parameter flogtanh_LIMIT_MAX = 'h800 ,
parameter flogtanh_LEN = 'h164 ,
parameter flogtanh_SEL = 9
