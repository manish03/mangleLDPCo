//`include "GF2_LDPC_fgallag_0x0000c_assign_inc.sv"
//always_comb begin
              Ia2f891646e6ab8d9fb9ea77d93148790['h00000] = 
          (!fgallag_sel['h0000c]) ? 
                       Ibbc4b022828a232d4b3d3eccc478fd3f['h00000] : //%
                       Ibbc4b022828a232d4b3d3eccc478fd3f['h00001] ;
//end
//always_comb begin
              Ia2f891646e6ab8d9fb9ea77d93148790['h00001] = 
          (!fgallag_sel['h0000c]) ? 
                       Ibbc4b022828a232d4b3d3eccc478fd3f['h00002] : //%
                       Ibbc4b022828a232d4b3d3eccc478fd3f['h00003] ;
//end
//always_comb begin
              Ia2f891646e6ab8d9fb9ea77d93148790['h00002] = 
          (!fgallag_sel['h0000c]) ? 
                       Ibbc4b022828a232d4b3d3eccc478fd3f['h00004] : //%
                       Ibbc4b022828a232d4b3d3eccc478fd3f['h00005] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00003] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00006] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00004] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00008] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00005] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0000a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00006] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0000c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00007] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0000e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00008] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00010] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00009] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00012] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0000a] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00014] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0000b] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00016] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0000c] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00018] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0000d] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0001a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0000e] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0001c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0000f] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0001e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00010] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00020] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00011] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00022] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00012] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00024] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00013] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00026] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00014] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00028] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00015] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0002a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00016] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0002c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00017] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0002e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00018] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00030] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00019] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00032] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0001a] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00034] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0001b] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00036] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0001c] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00038] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0001d] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0003a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0001e] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0003c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0001f] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0003e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00020] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00040] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00021] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00042] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00022] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00044] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00023] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00046] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00024] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00048] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00025] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0004a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00026] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0004c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00027] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0004e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00028] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00050] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00029] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00052] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0002a] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00054] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0002b] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00056] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0002c] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00058] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0002d] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0005a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0002e] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0005c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0002f] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0005e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00030] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00060] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00031] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00062] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00032] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00064] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00033] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00066] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00034] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00068] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00035] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0006a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00036] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0006c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00037] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0006e] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00038] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00070] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h00039] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00072] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0003a] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00074] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0003b] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00076] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0003c] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h00078] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0003d] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0007a] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0003e] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0007c] ;
//end
//always_comb begin // 
               Ia2f891646e6ab8d9fb9ea77d93148790['h0003f] =  Ibbc4b022828a232d4b3d3eccc478fd3f['h0007e] ;
//end
