 reg  ['hff:0] [$clog2('h7000+1)-1:0] I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd ;
