//#;; Ic23fa9996925b610710d93e28c59a3e2 I10df3d67626099df882920ba6552f16d I93762d802eed04b3e1c59d1d46b35248 Ic9f869114804f0a61ce9b03def9d71f5 I9fc5887c030f7a3e19821ebec457e719
/*I816842ff6f8526885b6ad2d49236bc84*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /Ic1111bd512b29e821b120b86446026b8/Id67f249b90615ca158b1258712c3a9fc -Ibea2f3fe6ec7414cdf0bf233abba7ef0 *I66986ae1d2ec0253762b97e22f881595* *If4ed727b4ff4652b44f0b32f7198402e* ; If83a0aa1f9ca0f7dd5994445ba7d9e80 I21f66e7dd81ae29064c26b66d9b3e967.I288404204e3d452229308317344a285d -If83a0aa1f9ca0f7dd5994445ba7d9e80 Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.sv > Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv ; Id6bfe3ce1bf5714887f4ffbb7b94feab -I958fb7ed1fb6d4960d15ffd3254be634 -Ie1e1d3d40573127e9ee0480caf1283d6 -Ia823f97963868b5794f5a36e4dbe5dec Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv -I2db95e8e1a9267b7a1188556b2013b33 Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv.Idc1d71bbb5c4d2a5e936db79ef10c19f

 /*I816842ff6f8526885b6ad2d49236bc84*/

/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I54a78636e8c6bd0efb73150b779d5eb5 */
//`default_nettype I334c4a4c42fdb79d7ebc3e73b517e6f8
//`timescale 1 ns / 1 ps

module  sntc_ldpc_syndrome_tb #(
// NR_2_0_4/I58d53a433022417c56e36facb426c2b8.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 
// 208
// 168
parameter SUM_NN         = $clog2(NN+1), // 8 : I307afb7f348272492f3cca58ef2f95d8
parameter SUM_MM         = $clog2(MM+1), // 8 : If78618843e4df2223e60ec190987c019
parameter LEN            = MM,
parameter SUM_NN_WDTH    = $clog2(SUM_NN+2),
parameter SUM_MM_WDTH    = $clog2(SUM_MM+2),
`include  "NR_2_0_4/sntc_LDPC_dec_param.sv"
parameter MAX_SUM_WDTH_LONG = MAX_SUM_WDTH +1,
parameter SUM_LEN= $clog2(NN+1)

) (

input wire clk_tb,
input wire rstn_tb
);

`ifdef ENCRYPT
`endif


bit I9849f97a8c5546c9906a059d1dd3ec64 =0;
bit [31:0] [150/*int*/:0]  I1bd3a0484883ca6deaada8395a8f6e85;
bit [31:0] [150/*int*/:0]  I461b1990fe86af962cd15a16a26dceb8;
bit [31:0] [150/*int*/:0]  I7e9293e90055a83d4943872232ff638f;
bit [31:0] [150/*int*/:0]    A;
bit [31:0] [150/*int*/:0]    I21c2e59531c8710156d34a3c30ac81d5;
int I680d7a67cf333b19f87ab59686c7b332     ;
int Ia8faf93382d2e794cad57d11e102656e    ;
real I041d491d3db37dd3d487a281d85f883d ;
string I66728d981980ea61d5c4e78a5192f5ed;
real Ice82750cacab30e6be8da3bb371f8441 ;
string I0cd3056ebfd4015fc53f149b8821d540;
real I008042664f7e640b5003f73aca5840cc ;
string Id77537bd9ea00a288f68886c448a9839;
real I063199a0348003d635c167af585e43d9 ;
string I8373077ab53f3c51daa3d544264ea7e5;
real I6bdb288f8bcad3a49a602451074bce26 ;
string I392cc984ed7cbdda0c0e1a0ad019faee;
real Id3f8037c35dfff19c21fcfbc7c26f09b ;
string I62b53a8231278f8228979bb7cbfa785d;
real I4d10c3daef7f20ac1f4d385c1bda95a3 ;
string I8c6f6a125c7be2a3803d128b5e8ed1e9;
real Id9f27d2391a03bc98a5bb6bc5925774d ;
string I26a2e345d1b41b3c45264040deccd7b1;
real I4861b5aec231ac5130ba30f990bbc161 ;
string Ib2d46624331c36e2c37e3b075d9e100e;
real I1814ce52608d992a2342fb439230eed0 ;
string I0d4e7dd3191e0053c4c1fa78f8a88f0b;
real I13164a39f30c204521076cfc674a22b5 ;
string I554a89331063a22c45fbfb822c5daf56;
real I04665defb04781dc87dd97e01f9c97bf ;
string I5c3639d7864bb49306fd6e52d5f5b53d;
real Ie4a8bc7b5eba426f1f22ed4237c1e395 ;
string I330e65820422fd85f34528f60f4deb31;
real I4ca566c9b7a8dafe56cce925952bb54a ;
string I0e6d5034ebd18f0c9e0d43a0e5067e48;
real Ie85ec7f87458e4cc2e0381661e23dc68 ;
string I124e3f4de0cc7a197b7b5060a18a2936;
real I32ccc376bc67772962ac3b55bc4db12d ;
string Ib752169206b316257c2e892cedd9d7b3;
real I9ab10bf13c49cd9bd351b10e1bbe02c4 ;
string I0a87abcd902686ade01f17f11b30141d;
real I1bd52652d791448ba8b2e988ed0f4c45 ;
string I1eb90eef09fc3762def8acaad9e815de;
real I3c44027069b2d0a279d21977b15159c6 ;
string I6359a292a3e344d6fc65567ce911292f;
real I8e234521cc7c01a8d46ea6e32a0790f2 ;
string Id455fea6020d386c588f4b7685cc7c94;
real I60a4ef194097807f60d55a344f272ee8 ;
string Ica491b503c88cb6f0090347e25ec9194;
real I78c7b8c2f6c08e06dd3fe94b1780df36 ;
string Ibc47d9c1b66633cfe9b8c840e9ca4a94;
real I13ac75f3d74c5d40d59f2ef13825e967 ;
string I4ae3f1e57e01a982c6753ce998871490;
real I3abeb1cddd05f3ed3cf351e185ec8b9a ;
string I1613b4ca977ab0484f7287417b03445d;
real I0fb8fd5b10a560d9e4b34f89bfb6ebe6 ;
string I8d462af6fa9413b64b364d1d4dc06530;
real I4c84184b303150deecb16c311fc3d2e7 ;
string Ie462f3ff20c9eae160e60cd32befa082;
real I35f34a1fbc2316b056ac8f3e054768aa ;
string Ibda3c321a1d7c69ad194e3e96338ae85;
real Iaf193bf234240fda68149737220f26f7 ;
string I76d01d348b392373da3e5ba3226426ea;
real I066bd0bc1075b584aace9a70ce458100 ;
string Id4d43c17828a34dc74c91bd196b5fa15;
real Iab501fd728018643547393afe617dbb5 ;
string I24743cc72845877cbeee57b56cc1e311;
real I9531876b777a57bc770c69bffbd75d7d ;
string I129c2799cd95848db9acbef09b9fc833;
real Ia9b3ded8c4b4df0f340976360a8ae120 ;
string I2aba999392b7a9c3be1a485b9996bb6c;
real Ib7d5d99937157987bb421cf5d676207b ;
string Ie936cb5058108147f9310e05ea046e39;
real I068bdaa8253aedc29eebb5023dd83903 ;
string I022ee38d1d2bbd7e704773aef3f234a4;
real I310aae59087e8b02e297483a7fc0b3c2 ;
string I43d5e4240d17f6385a6b3a70da4490b4;
real I656b7e9c8184a1be3462dd391dbac80b ;
string I809e11476ee6548c42fa12b46f5162e6;
real Ib13bffc02fcbb12de67957ba695dbe11 ;
string I755d866626f4f976d4f3b1be75b32cbf;
real Iaebbaf7858e6d1d0cf44801448b6a588 ;
string Ida9094a1a1190bf89a5ecfa778d06c07;
real I07bb3693c696eea928ba3839afa10398 ;
string Icaf4d656643680116d687d1ea2135359;
real If1e9ad94e37fd7ef189ed150fc2bc4ec ;
string I6588d1f52a799c597ebfcfebe7916dbe;
real Ie5e178b74c6eb4554b0fa6e4c4d3ed78 ;
string I77a58fdba96cd4b7cb84eeb3065f5490;
real I41a1b293c4b61920f6e0504f51d199f7 ;
string Ia673c74384dba43d639347c5bcc7a587;
real I2a4e9185fb4387e03992ef825d9a64dd ;
string If8aba14cfa5bdef2e3c74b7a0c560723;
real I27ce163b3e8fb3b08a120bb78ca3883c ;
string Ia0bbff612d39d36ff506a0f61649ef8f;
real I0a5c2bf1d14366e9bdf63a95c9f1dd08 ;
string Ieb90619950c09bffc6192a49cc88e961;
real Ie8327512d3df7102e73595b046d78f90 ;
string I3db1cbad580dda99490bc1d0e074ff2e;
real I091196adb9bd28ac06b0d8b6c9a60909 ;
string I561269286fae11c600f849eeae0e1b46;
real Ie4a70a6e05e18f1a8541c0d4d1a37c37 ;
string I15873980a25f1e4156dce47a6373b601;
real I6562b0db0d66d401ea4e45bda429cd53 ;
string I881c2dfcd7181dd754f6e9452ca36c26;
real Ib32a2ef64966dd61fc49559994111d66 ;
string I93744d7253e201beac98054c8edb3a4b;
real I81d7c343f6311a7274e96066b259038e ;
string I31ee8dcc5cc4a1fcdfd80486c06fa76b;
real I108f200e4b9a869ee151b560fb82b2d1 ;
string I773aefae4577fb5ba1abd0dc8480c355;
real Ia82c634bf043c61daf94f71025052af7 ;
string I5f55c4b0ca264cd374a95711d8cea6dd;
real I9f9c8417258c5b21c37f921bcca955cc ;
string I8a1aaba08d5fbff7da33d6c150c648b1;
real I7116bd6af04920ff7eb964f88570020e ;
string I06091fccb3c6f2af1053ce83342ed71a;
real I3fefc853340d936b45283ea808e17b9e ;
string Icdd5f27fd0f7c8b85c633caaee59c2b6;
real Ie573808e06c1896c1981bac6d6d777df ;
string If1c1e1e48d3f6fe43431ef5b93151f61;
real I09d4ddac066a0ac6ff6aac51709347c1 ;
string I615147a0262ea201531dc8172141ec28;
real Id57dc980e439baadfd865dbe749c87d7 ;
string Iefcb8381273e0f1929e4acc1301393b9;
real Idc16547311e95f3b4e24a2488d6dcc61 ;
string I82008685277ca9c199c3a2d790f210c3;
real I8f52f481d4f0de58819e2685651ca17a ;
string I1a6a2c2ee2945c3eb67847f11c2af931;
real Iea89d6322a76ad368385ef97dc4f9eef ;
string I1f5101292324bafcc87f333d2c941b7b;
real I1d1f6dc8396366c974c1526e1a639468 ;
string I161ecc1c467dfbaa7160f51c2cbde8cf;
real I0c76adcfb28bfd3ababde368f878c47a ;
string Id45c2931318e51f29760afe71e869c29;
real I5c0f2d32067dd55b33f715f05b529cd3 ;
string I9a94a17450c0d37dce6fc481aac687d6;
real Ia9fd736f9384262688f43108e6f0f512 ;
string Ica8e3000994dcb8c743e4bbee5f02e01;
real I743c59645aa659f7d3a013cdfbd46620 ;
string Ib79be162ecead96363f46f6f8a6bef7b;
real I76f5ef93e6cbfeeafec0c076ee2401f9 ;
string I3ed1a2aa3d57e5939bc936e4db08b218;
real I33f1ff2c21f954fcba24cc9404e0420a ;
string Ia52604e308b534f02c9626d65a4e4772;
real I171ebffcc1b7a4782f350ecb33a368a8 ;
string I174b39d9bd5c7c1c3314eff3bd45deea;
real Ic01c6dad4081aa8cbf8d1b690333dbfc ;
string Ie1499d5b68e178b2b6d922f8666fbd20;
real I99009951f130f09a85b61ee7847b138d ;
string Ib73f2379e9f8e5f964b55bb82c339d15;
real Ibe1ed5c23d4f3deacc8a17e010a19e6d ;
string I91e2b00feb733024632ad2390799ebb5;
real Ic739a419f112ec796e4e6d1f16dfac5f ;
string I213d7f04f870f9be53686e07da0eecf1;
real Ib6100b0fecb09bf81a1d496a74bd68bc ;
string I5db98931b33031bf3a895b09ce00da30;
real Ie11211db877ae7931b2212828767e077 ;
string I8b78afe0d27c51c64bd77bb6f0394bba;
real I5146a988cb19b206d3b77a71f17680c3 ;
string I522a698492d6c5bc41add99134f6aa57;
real I9f2575295a210e3b2d2f4f76a09b3e2f ;
string I0e0f3f1c743528a1b11232a445c87807;
real I7dac8ad08c2bbcbb424738b5c24c7468 ;
string I69a9811dbaf4e3c974039c21310f86a4;
real I35b723ce016238903d276496dc65476a ;
string Ie9b5edd2cfbfcfab73b3489e0783571d;
real Ied751b3d3e14d5a29e0d7e50a0f71070 ;
string Icdb612e518fee711afd0b4666212a96a;
real I9df88da58c6c6520e9b44fa10d062f8f ;
string Ibcc6bb0948604a9fbe763162ed5ff08d;
real Ieb3883a9dc81b97abb5111b806a20210 ;
string Id35867526784204032082c8f9bce8e89;
real If9a817ef2cfbcb526a80ae94c20fd24d ;
string Iac98b08dca97cc20db7d8478bbffee1f;
real I9857f502c20529706d320c258863b1c8 ;
string I3cbea822a06bc7de47bfc893549f1009;
real Ida567e4e8b2a7b2abbc304b5d5d8a817 ;
string Iab03b367005c2a285ac2e12ea67ba587;
real I94ac4090b1bae29fa174cc017ccd7264 ;
string Ie2e582fd36b101c8c695472e28687414;
real I208eb0ab24696d9faa69c276606b5467 ;
string I65d195472be43c160475f7a7daaaee87;
real I52bedb38090c611edaa00fd6102f2a8d ;
string Idbe6259e292d1a3d8784f5c8695b9a06;
real I4af91415fc0408b64bb4be0fe66b270b ;
string I11a30b96d26b358acd1ec10875b44c70;
real I31472bac41773613648ff29fdc5ed119 ;
string I632789bf1e28a9d9e156ef49bf25c93a;
real I566bd7f2a2b77a0a6a371d140395508d ;
string I12a7cf28ef0aed9680955631f89fb6b5;
real I8679ec448b6c689fa27b82393e05d116 ;
string I36979f9dd020af47874e3c4d1d83a492;
real Ia8780ff6e2b75f06913b5ed3d131d2aa ;
string I2997b11c880fd30fde0d30ec20009f50;
real I3f49e9fc58809b8d7286437f164eef4b ;
string I6fa422edfa1fa5129a78468f9d3e2289;
real Ic3704d821df6c5ee9a3f4c52860b8ef4 ;
string Ibf0a8a6654a6b93ed000f217e6a93972;
real I6e13b1bb5582c7ab55d08d9c3e6a8a8d ;
string I6b85238e2a7f79b63af4e812bba3e71c;
real Iba0667763a0df496bf0df27c261109f6 ;
string Id213b0550c89d4a0557ea8a46b817222;
real I88acd1105daddfc526e2f72e1bbe4370 ;
string I5aebc60ecfa7112d99ff2abcb2e8f7be;
real I417e21779c134ca6cb5696c9ea126e7b ;
string Ib4d268d5d7da92b1c9706a573e4a7053;
real I7a3a6c74f11d67bea8d0a3411f4c19de ;
string Ibb0b846893f2dcacae3989e01ea81db4;
real I68fad9d0dc23e65d35492ae6ce7ede43 ;
string I5b7849b5198e5f06b7d170528f72433d;
real I016bd64256942460cafa870fa9767f29 ;
string I6cb00ad8c59156406d2c54d12d958943;
real I69175952533ce230691b0d41185f73ed ;
string I02191f115223e5d16a7aa846c916ed50;
real I006d3763207bec11f72fe478fb7059f8 ;
string I2a4e7eb3e181e16217ecc212c6564a37;
real Ieb127e866e30c8000d046d152182f718 ;
string Iaa5a13030697a4b11cd99437b9c200cc;
real Idcd6887fc060a9862c0c539cdcce80cf ;
string I3573e9457f4107cf46802535a9c9dac1;
real I0d637be1e321aa1689e428a47afe9a1d ;
string I4de741ee35eb3ad7b1f365b2e31a272f;
real I8d168f2f3c4afe033658c3d411cde850 ;
string Ibcba6fcb883796c52a482f327c467d9c;
real I1790e02762e0adfdac36c6e3429afada ;
string Ibdde55097b6214929866994501913d2d;
real I7fb4bdc82336c690c3037724c8ff433d ;
string I1ff6754a6dfb612192e4702ff6b28c00;
real I20c28f0cc20cd997bcbc2e7703330402 ;
string I4adb4aae5bb881423b21b82e1923d0f1;
real I41390b9833367be94eae4cc1a1ca377c ;
string I593a607afa403f5942fdfc2de0f444ac;
real I1f6f25f1e784fc3f7ab800e715cd8158 ;
string I66057ab775253511c93d0aaa181523af;
real I84be8553fb5d8418b22b0e96753014b9 ;
string Ia98f52f37f95b9ba8c49875a384b2de5;
real I861e8b0d0ae393a89e5ce7093bbb3b06 ;
string I9f4263e11444b59093efb75304ed5b78;
real I88fa892c4a6e6a789503fb4f719b3634 ;
string If3d9f9527196c1eee46e34ed8b1ca20f;
real I112e771ffd1147507331c3f407d0fe5f ;
string Ibfad8563c458f63154c6cbd86cc7d97c;
real I3bc80849aa22396280553cccdc2345a3 ;
string I52fe04ff3fa957f55f386e357d7fe260;
real Iae254415a32ebbe3d7e166d08a4d093f ;
string I3d05f05876ed3434a983340fea38491d;
real I9e8d5ba657ebad083c6a5b12b6ac72c5 ;
string I92de9ad4dd3c4da78726f7161bae2087;
real I1cd574808e24f3b7ffde2547ad58548f ;
string I298fb7b4a1196668dbed710a01ea5f9c;
real Ic8c428f6169f8b91c686a9fb94615e9c ;
string I9cfad560131bdb24ad2ae33b2ea15300;
real I4d0af269b285c85593ab2ad93b6192ca ;
string I43f6aac9c0bb10e9d79636e15a0e049b;
real I561564e9f78c9e35ad742a704258084b ;
string I7835cfd4a0de695bcf1fddfb49e82242;
real I1d51669925bdf956ef1cecba7deba70a ;
string Ie2ec46b365bf63516903b03cef0521a9;
real I9c2a96246fbd4376fa7736a83fc0e9fb ;
string I730b21a917c2c56cf4313fb4e728d040;
real I16ffe5da86128750d03105acf9b162da ;
string Id158da98fcadcc931d69f7642e46e08a;
real I286203337d5c5e036453c252f347a63a ;
string Id989b3d79501498a3db58048a0b2e2e9;
real I1bf77e202622f9067f475bd8f2b4e4c9 ;
string I5dfff598c558eb9ff8f2002e4ab13e88;
real I529eaf19e7234ee8dd594b2104bd1c26 ;
string I5d2fa444646c4074d9c243be6b59f61f;
real I94d8fb8446d827c19d48b424cbe1b025 ;
string I6e54873fccd867eee40c355ae915b7a1;
real Id31e57ffd7f012b7e2ef207e61a5de59 ;
string Ifffa8c78712a8a2ca3a881cf3f390725;
real I7d91ea5d5bda466296344bc728c77089 ;
string I7c85a36febe45f21b8fda8a0ae143f44;
real Iaa08501162ec50e4ddc9ebf88d7593e4 ;
string I361d2071e439cc8a1ea223aa13fe1b08;
real I0e9ff8e0b3fb7ffe35922a4daeebd3df ;
string Iab4fd20360fdc46a4bfb9d97677aa531;
real Iad1e9049c550c2994b7eff96094199b6 ;
string I5588d9ef2dcf58df8090b4452a18ba51;
real I32dac8554f5ce05d74f1d0ca449237e7 ;
string Ic090d1e475405407995d2784d2e6df5d;
real Id1797d69f67972dc35de74f028bf3374 ;
string Ieaeef2f90dadf2e75c7e7e1e417bc5a1;
real I1c565efc669880d59741b637cf60883a ;
string Ia6d28169bb945021a239794f458634fd;
real Ie93b565ae5611ffe367eb4e5c83f4149 ;
string I5b0545f33f97d4fbf571ae637c7af810;
real I7f54926b9d6692ac20f8e9c27e6fcdf6 ;
string I25ccf3347306971223fa06b7665616e6;
real I6e7c12d81076a8cff47daed26c020dfd ;
string I42b4f206dfb56e9e88d0b67108b1767d;
real I037ce03738340baf17eaab9598122faa ;
string I06308bd8357c99fd486b9eb2c9324e0b;
real I3ac9b34c65e3c564e334281261c90abf ;
string Id90e9a7166cfcca424f45d7a3ff8055a;
real I1b9924e4d0d0cbe29c9ff1a0b5f5917b ;
string I93c0aa630ce2748f1edbc787ee0cdabf;
real Ie2c08f886a5b81db14d1fb5d784d16af ;
string Iaebf4876732c2244bb8b59d8eb127a5e;
real I126ab1bc306a37834ebf2f24f34a5fde ;
string I3c6a1299ee32cec3072beee04a62ad99;
real Iaa72597813cc3921f17977ad505ba2cc ;
string I1cc6bdbc8b277fa8394f82725b14976c;
real Ifa402fc88dbd79eb79c809e27f27a36c ;
string Ic2c9f984d9bc815d646e9d699316363c;






// -1 : I8560273e5cfe310f2c9d5ab5defa48f3
// NR_2_0_4.I46d9a76ee9f25d6fe22e820d7ccc99b3 : I7398678ae6fe7c505be08e7bebdcfca3 Ib068931cc450442b63f5b3d276ea4297


// Id17d8f0661f8f44dd7dc5110c8825246 : Ic3938dd81fe1366e93d2e29a6ffe2005 2 0 4.I46d9a76ee9f25d6fe22e820d7ccc99b3
// I794f7c3f9d2c2287034081a9c64f4073: 2

// I6a0ad5eaf9d47f99b7f194646dacab10: $NR_Z





reg  [NN-1:0]                 tmp_bit;
reg  [NN-1:0] [1:0]           I61e23fc401e882840b471b3b125a68a9;
wire [MM-1:0]                 syndrome;
reg  [MM-1:0]                 exp_syn;
wire [SUM_LEN-1:0]            HamDist_sum_mm;
reg  [SUM_LEN-1:0]            HamDist_loop;
reg  [SUM_LEN-1:0]            HamDist_cntr;
reg  [SUM_LEN-1:0]            HamDist_loop_max;
reg  [SUM_LEN-1:0]            HamDist_loop_percentage;
wire [1:0]                    I7de33615d7fbc1cb7bc608d12f1993d2;
wire                          I988ac9ae2dc175e23b845ba27cb36625;
reg                           I06e0a59e15a77350b25fe9ca79a311b3;
wire                          I53efd0678e8d3a37c9fc26da5613b3c2;
reg                           clk;
reg                           rstn;
int                           I3240712af92cc8a4d47f14e9b94ec0e6;
reg                           clr;
reg                           Iea2b2676c28c0db26d39331a336c6b92;
wire                          valid;
wire [31:0]                   percent_probability_int;

reg  [SUM_LEN-1:0]            HamDist_iir1;
reg  [SUM_LEN-1:0]            HamDist_iir2;
reg  [SUM_LEN-1:0]            HamDist_iir3;
reg                           Iadfe5fe147b14daeca7d68a0b2f6579e =0;

always_comb begin
          HamDist_iir1 = 85;
          HamDist_iir2 = 15;
          HamDist_iir3 = 5;

end

wire valid_cword;
wire valid_cword_dec;
wire [NN-1:0] I8d1e6fa299262b2bef3b696c48864ad9;
reg [NN-MM-1:0] y_nr_in;
reg [NN-1:0] I81dab9b4f78627240b44ac785b16acf9;

sntc_ldpc_syndrome_wrapper i_sntc_ldpc_syndrome_wrapper
(


                                  .y_nr_in                (tmp_bit),
                                  .syn_nr                 (syndrome),
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I3bc180bd00be2c60a3a5a68e0dd49503 */
                                  .clr                    (clr),
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 I18c0d99dcef0c6b3cc1cadd623fdbf9f I3bc180bd00be2c60a3a5a68e0dd49503 */
                                  .valid_cword            (valid_cword),
                                  .rstn                   (rstn),
                                  .clk                    (clk)
);





`ifdef SIMULATION
 int I9e5210b8cd60e37903cfe362297f07aa =1;
initial
begin
  clk = 0;
  I3240712af92cc8a4d47f14e9b94ec0e6 = 1;
  forever
  begin
    clk = ~clk;
    if (clk) I3240712af92cc8a4d47f14e9b94ec0e6 = I3240712af92cc8a4d47f14e9b94ec0e6 + 1;
    //if (clk) if ((I3240712af92cc8a4d47f14e9b94ec0e6 % 1000) === 0) $display("I4f62dc0a0e700849a9987d10e9dc369b:I3240712af92cc8a4d47f14e9b94ec0e6:%05d %t", I3240712af92cc8a4d47f14e9b94ec0e6, $time);
    if (clk) $display("I4f62dc0a0e700849a9987d10e9dc369b:I3240712af92cc8a4d47f14e9b94ec0e6:%05d %t", I3240712af92cc8a4d47f14e9b94ec0e6, $time);
    #5;
  end
end
initial
begin
  rstn = 0;
  clr = 0;
  repeat (10) @ (posedge clk);
  rstn = 1;
end


always_comb HamDist_loop_max        =  10;
always_comb HamDist_loop_percentage =  110;

initial
begin
I7e9293e90055a83d4943872232ff638f[00]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 0]= 9396;A[ 0]=8832;I66728d981980ea61d5c4e78a5192f5ed="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[01]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 1]=10566;A[ 1]=8832;I0cd3056ebfd4015fc53f149b8821d540="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[02]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 2]= 9392;A[ 2]=8832;Id77537bd9ea00a288f68886c448a9839="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[03]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 3]=12368;A[ 3]=8832;I8373077ab53f3c51daa3d544264ea7e5="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[04]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 4]=14460;A[ 4]=8832;I392cc984ed7cbdda0c0e1a0ad019faee="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[05]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 5]=20768;A[ 5]=8832;I62b53a8231278f8228979bb7cbfa785d="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[06]=3840;I1bd3a0484883ca6deaada8395a8f6e85[ 6]=19200;A[ 6]=4032;I8c6f6a125c7be2a3803d128b5e8ed1e9="I8930f12f516428fc23bc164621b19d4f" ;
I7e9293e90055a83d4943872232ff638f[07]=3840;I1bd3a0484883ca6deaada8395a8f6e85[ 7]=19200;A[ 7]=4032;I26a2e345d1b41b3c45264040deccd7b1="I8930f12f516428fc23bc164621b19d4f" ;

I7e9293e90055a83d4943872232ff638f[ 8]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 8]=14556;A[ 8]=8832;Ib2d46624331c36e2c37e3b075d9e100e="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[ 9]=8448;I1bd3a0484883ca6deaada8395a8f6e85[ 9]=21048;A[ 9]=8832;I0d4e7dd3191e0053c4c1fa78f8a88f0b="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[10]=8448;I1bd3a0484883ca6deaada8395a8f6e85[10]=25344;A[10]=8832;I554a89331063a22c45fbfb822c5daf56="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[11]=3840;I1bd3a0484883ca6deaada8395a8f6e85[11]=19200;A[11]=4032;I5c3639d7864bb49306fd6e52d5f5b53d="I8930f12f516428fc23bc164621b19d4f" ;


I7e9293e90055a83d4943872232ff638f[12]= 501;I1bd3a0484883ca6deaada8395a8f6e85[12]= 864 ;A[12]= 546;I330e65820422fd85f34528f60f4deb31="I8231507cfb68527311772d51ac55cb18" ;
I7e9293e90055a83d4943872232ff638f[13]= 231;I1bd3a0484883ca6deaada8395a8f6e85[13]= 576 ;A[13]= 252;I0e6d5034ebd18f0c9e0d43a0e5067e48="If815a5240829d01419117bb9e280812c"  ;
I7e9293e90055a83d4943872232ff638f[14]=  57;I1bd3a0484883ca6deaada8395a8f6e85[14]= 288 ;A[14]=  84;I124e3f4de0cc7a197b7b5060a18a2936="Icea89eb072364858f820071032afb467"  ;
I7e9293e90055a83d4943872232ff638f[15]=  28;I1bd3a0484883ca6deaada8395a8f6e85[15]= 140 ;A[15]=  84;Ib752169206b316257c2e892cedd9d7b3="Icea89eb072364858f820071032afb467"  ;
I7e9293e90055a83d4943872232ff638f[16]=1003;I1bd3a0484883ca6deaada8395a8f6e85[16]=1728 ;A[16]=1096;I0a87abcd902686ade01f17f11b30141d="I71aae66d47b808b53a20d58a74902074" ;
I7e9293e90055a83d4943872232ff638f[17]= 462;I1bd3a0484883ca6deaada8395a8f6e85[17]=1152 ;A[17]= 504;I1eb90eef09fc3762def8acaad9e815de="Iafbc30d0bdee0217a07538df70f416cc" ;
I7e9293e90055a83d4943872232ff638f[18]= 115;I1bd3a0484883ca6deaada8395a8f6e85[18]= 576 ;A[18]= 126;I6359a292a3e344d6fc65567ce911292f="If27d61c6ed0b84b26da1e70364750452"  ;
I7e9293e90055a83d4943872232ff638f[19]=  57;I1bd3a0484883ca6deaada8395a8f6e85[19]= 286 ;A[19]=  84;Id455fea6020d386c588f4b7685cc7c94="Icea89eb072364858f820071032afb467"  ;


I7e9293e90055a83d4943872232ff638f[20]=8448;I1bd3a0484883ca6deaada8395a8f6e85[20]=25344;A[20]=8832;Ica491b503c88cb6f0090347e25ec9194="I50f595021a9bf9cb7f3cc62e720730eb";

I7e9293e90055a83d4943872232ff638f[21]=8448;I1bd3a0484883ca6deaada8395a8f6e85[21]=14556;A[21]=8832;Ibc47d9c1b66633cfe9b8c840e9ca4a94="I50f595021a9bf9cb7f3cc62e720730eb";
I7e9293e90055a83d4943872232ff638f[22]=4162;I1bd3a0484883ca6deaada8395a8f6e85[22]=10368;A[22]=4416;I4ae3f1e57e01a982c6753ce998871490="I91962bb5d2be35247a651d8174c89d1a" ;
I7e9293e90055a83d4943872232ff638f[23]=1036;I1bd3a0484883ca6deaada8395a8f6e85[23]= 5180;A[23]=1096;I1613b4ca977ab0484f7287417b03445d="I71aae66d47b808b53a20d58a74902074" ;
I7e9293e90055a83d4943872232ff638f[24]= 518;I1bd3a0484883ca6deaada8395a8f6e85[24]= 2590;A[24]= 546;I8d462af6fa9413b64b364d1d4dc06530="I8231507cfb68527311772d51ac55cb18" ;

I7e9293e90055a83d4943872232ff638f[25]=4326;I1bd3a0484883ca6deaada8395a8f6e85[25]=4162 ;A[25]=4784;Ie462f3ff20c9eae160e60cd32befa082="Ia4dcc6cd7be7fc538df90fabd97996d2";

I7e9293e90055a83d4943872232ff638f[26]=1036;I1bd3a0484883ca6deaada8395a8f6e85[26]=5180 ;A[26]=1092;Ibda3c321a1d7c69ad194e3e96338ae85="I71aae66d47b808b53a20d58a74902074" ;
I7e9293e90055a83d4943872232ff638f[27]=518 ;I1bd3a0484883ca6deaada8395a8f6e85[27]=2590 ;A[27]= 546;I76d01d348b392373da3e5ba3226426ea="I8231507cfb68527311772d51ac55cb18" ;

end
initial
begin

  static int Ifb48ed869c44bdc930da7ccc778d5014;
  static int I2cb9df9898e55fd0ad829dc202ddbd1c;
  static int I7a1d27b4c6e920486ea97597d7e919ee;
  static int I3dc53e26c8e2ca3d2b6896df6f30eca4;
  static int Ie18a4d4830028f90f158755e5e80fec5 = 0;

  Iea2b2676c28c0db26d39331a336c6b92                          <= 1'b0;
  I7a1d27b4c6e920486ea97597d7e919ee = 0;

  repeat (1) @ (posedge rstn);
  repeat (10) @ (posedge clk);

  if (Iadfe5fe147b14daeca7d68a0b2f6579e) begin


              I61e23fc401e882840b471b3b125a68a9  [0] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [1] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [2] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [3] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [4] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [5] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [6] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [7] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [8] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [9] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [10] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [11] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [12] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [13] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [14] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [15] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [16] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [17] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [18] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [19] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [20] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [21] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [22] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [23] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [24] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [25] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [26] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [27] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [28] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [29] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [30] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [31] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [32] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [33] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [34] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [35] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [36] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [37] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [38] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [39] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [40] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [41] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [42] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [43] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [44] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [45] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [46] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [47] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [48] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [49] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [50] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [51] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [52] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [53] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [54] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [55] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [56] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [57] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [58] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [59] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [60] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [61] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [62] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [63] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [64] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [65] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [66] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [67] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [68] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [69] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [70] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [71] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [72] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [73] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [74] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [75] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [76] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [77] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [78] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [79] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [80] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [81] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [82] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [83] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [84] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [85] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [86] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [87] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [88] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [89] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [90] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [91] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [92] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [93] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [94] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [95] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [96] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [97] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [98] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [99] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [100] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [101] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [102] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [103] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [104] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [105] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [106] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [107] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [108] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [109] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [110] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [111] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [112] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [113] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [114] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [115] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [116] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [117] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [118] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [119] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [120] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [121] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [122] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [123] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [124] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [125] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [126] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [127] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [128] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [129] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [130] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [131] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [132] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [133] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [134] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [135] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [136] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [137] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [138] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [139] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [140] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [141] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [142] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [143] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [144] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [145] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [146] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [147] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [148] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [149] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [150] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [151] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [152] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [153] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [154] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [155] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [156] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [157] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [158] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [159] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [160] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [161] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [162] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [163] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [164] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [165] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [166] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [167] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [168] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [169] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [170] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [171] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [172] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [173] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [174] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [175] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [176] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [177] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [178] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [179] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [180] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [181] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [182] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [183] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [184] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [185] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [186] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [187] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [188] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [189] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [190] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [191] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [192] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [193] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [194] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [195] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [196] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [197] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [198] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [199] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [200] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [201] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [202] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [203] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [204] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [205] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
              I61e23fc401e882840b471b3b125a68a9  [206] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
              I61e23fc401e882840b471b3b125a68a9  [207] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                 // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01

         exp_syn [0] <= 1'b1;
         exp_syn [1] <= 1'b1;
         exp_syn [2] <= 1'b1;
         exp_syn [3] <= 1'b1;
         exp_syn [4] <= 1'b1;
         exp_syn [5] <= 1'b1;
         exp_syn [6] <= 1'b1;
         exp_syn [7] <= 1'b1;
         exp_syn [8] <= 1'b1;
         exp_syn [9] <= 1'b1;
         exp_syn [10] <= 1'b1;
         exp_syn [11] <= 1'b1;
         exp_syn [12] <= 1'b1;
         exp_syn [13] <= 1'b1;
         exp_syn [14] <= 1'b1;
         exp_syn [15] <= 1'b1;
         exp_syn [16] <= 1'b1;
         exp_syn [17] <= 1'b1;
         exp_syn [18] <= 1'b1;
         exp_syn [19] <= 1'b1;
         exp_syn [20] <= 1'b1;
         exp_syn [21] <= 1'b1;
         exp_syn [22] <= 1'b1;
         exp_syn [23] <= 1'b1;
         exp_syn [24] <= 1'b1;
         exp_syn [25] <= 1'b1;
         exp_syn [26] <= 1'b1;
         exp_syn [27] <= 1'b1;
         exp_syn [28] <= 1'b1;
         exp_syn [29] <= 1'b1;
         exp_syn [30] <= 1'b1;
         exp_syn [31] <= 1'b1;
         exp_syn [32] <= 1'b1;
         exp_syn [33] <= 1'b1;
         exp_syn [34] <= 1'b1;
         exp_syn [35] <= 1'b1;
         exp_syn [36] <= 1'b1;
         exp_syn [37] <= 1'b1;
         exp_syn [38] <= 1'b1;
         exp_syn [39] <= 1'b1;
         exp_syn [40] <= 1'b1;
         exp_syn [41] <= 1'b1;
         exp_syn [42] <= 1'b1;
         exp_syn [43] <= 1'b1;
         exp_syn [44] <= 1'b1;
         exp_syn [45] <= 1'b1;
         exp_syn [46] <= 1'b1;
         exp_syn [47] <= 1'b1;
         exp_syn [48] <= 1'b1;
         exp_syn [49] <= 1'b1;
         exp_syn [50] <= 1'b1;
         exp_syn [51] <= 1'b1;
         exp_syn [52] <= 1'b1;
         exp_syn [53] <= 1'b1;
         exp_syn [54] <= 1'b1;
         exp_syn [55] <= 1'b1;
         exp_syn [56] <= 1'b1;
         exp_syn [57] <= 1'b1;
         exp_syn [58] <= 1'b1;
         exp_syn [59] <= 1'b1;
         exp_syn [60] <= 1'b1;
         exp_syn [61] <= 1'b1;
         exp_syn [62] <= 1'b1;
         exp_syn [63] <= 1'b1;
         exp_syn [64] <= 1'b1;
         exp_syn [65] <= 1'b1;
         exp_syn [66] <= 1'b1;
         exp_syn [67] <= 1'b1;
         exp_syn [68] <= 1'b1;
         exp_syn [69] <= 1'b1;
         exp_syn [70] <= 1'b1;
         exp_syn [71] <= 1'b1;
         exp_syn [72] <= 1'b1;
         exp_syn [73] <= 1'b1;
         exp_syn [74] <= 1'b1;
         exp_syn [75] <= 1'b1;
         exp_syn [76] <= 1'b1;
         exp_syn [77] <= 1'b1;
         exp_syn [78] <= 1'b1;
         exp_syn [79] <= 1'b1;
         exp_syn [80] <= 1'b1;
         exp_syn [81] <= 1'b1;
         exp_syn [82] <= 1'b1;
         exp_syn [83] <= 1'b1;
         exp_syn [84] <= 1'b1;
         exp_syn [85] <= 1'b1;
         exp_syn [86] <= 1'b1;
         exp_syn [87] <= 1'b1;
         exp_syn [88] <= 1'b1;
         exp_syn [89] <= 1'b1;
         exp_syn [90] <= 1'b1;
         exp_syn [91] <= 1'b1;
         exp_syn [92] <= 1'b1;
         exp_syn [93] <= 1'b1;
         exp_syn [94] <= 1'b1;
         exp_syn [95] <= 1'b1;
         exp_syn [96] <= 1'b1;
         exp_syn [97] <= 1'b1;
         exp_syn [98] <= 1'b1;
         exp_syn [99] <= 1'b1;
         exp_syn [100] <= 1'b1;
         exp_syn [101] <= 1'b1;
         exp_syn [102] <= 1'b1;
         exp_syn [103] <= 1'b1;
         exp_syn [104] <= 1'b1;
         exp_syn [105] <= 1'b1;
         exp_syn [106] <= 1'b1;
         exp_syn [107] <= 1'b1;
         exp_syn [108] <= 1'b1;
         exp_syn [109] <= 1'b1;
         exp_syn [110] <= 1'b1;
         exp_syn [111] <= 1'b1;
         exp_syn [112] <= 1'b1;
         exp_syn [113] <= 1'b1;
         exp_syn [114] <= 1'b1;
         exp_syn [115] <= 1'b1;
         exp_syn [116] <= 1'b1;
         exp_syn [117] <= 1'b1;
         exp_syn [118] <= 1'b1;
         exp_syn [119] <= 1'b1;
         exp_syn [120] <= 1'b1;
         exp_syn [121] <= 1'b1;
         exp_syn [122] <= 1'b1;
         exp_syn [123] <= 1'b1;
         exp_syn [124] <= 1'b1;
         exp_syn [125] <= 1'b1;
         exp_syn [126] <= 1'b1;
         exp_syn [127] <= 1'b1;
         exp_syn [128] <= 1'b1;
         exp_syn [129] <= 1'b1;
         exp_syn [130] <= 1'b1;
         exp_syn [131] <= 1'b1;
         exp_syn [132] <= 1'b1;
         exp_syn [133] <= 1'b1;
         exp_syn [134] <= 1'b1;
         exp_syn [135] <= 1'b1;
         exp_syn [136] <= 1'b1;
         exp_syn [137] <= 1'b1;
         exp_syn [138] <= 1'b1;
         exp_syn [139] <= 1'b1;
         exp_syn [140] <= 1'b1;
         exp_syn [141] <= 1'b1;
         exp_syn [142] <= 1'b1;
         exp_syn [143] <= 1'b1;
         exp_syn [144] <= 1'b1;
         exp_syn [145] <= 1'b1;
         exp_syn [146] <= 1'b1;
         exp_syn [147] <= 1'b1;
         exp_syn [148] <= 1'b1;
         exp_syn [149] <= 1'b1;
         exp_syn [150] <= 1'b1;
         exp_syn [151] <= 1'b1;
         exp_syn [152] <= 1'b1;
         exp_syn [153] <= 1'b1;
         exp_syn [154] <= 1'b1;
         exp_syn [155] <= 1'b1;
         exp_syn [156] <= 1'b1;
         exp_syn [157] <= 1'b1;
         exp_syn [158] <= 1'b1;
         exp_syn [159] <= 1'b1;
         exp_syn [160] <= 1'b1;
         exp_syn [161] <= 1'b1;
         exp_syn [162] <= 1'b1;
         exp_syn [163] <= 1'b1;
         exp_syn [164] <= 1'b1;
         exp_syn [165] <= 1'b1;
         exp_syn [166] <= 1'b1;
         exp_syn [167] <= 1'b1;

  end else begin //Iadfe5fe147b14daeca7d68a0b2f6579e==0
     bit I798dd71209184f626a7f6bed517aa125;
         y_nr_in[0] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[1] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[2] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[3] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[4] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[5] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[6] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[7] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[8] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[9] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[10] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[11] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[12] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[13] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[14] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[15] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[16] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[17] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[18] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[19] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[20] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[21] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[22] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[23] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[24] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[25] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[26] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[27] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[28] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[29] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[30] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[31] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[32] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[33] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[34] = 1; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[35] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[36] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[37] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[38] = 0; //I8d777f385d3dfec8815d20f7496026dc
         y_nr_in[39] = 0; //I8d777f385d3dfec8815d20f7496026dc
     repeat (1) @ (posedge clk);
     for (int I865c0c0b4ab0e063e5caa3387c1a8741=0;I865c0c0b4ab0e063e5caa3387c1a8741<NN-MM;I865c0c0b4ab0e063e5caa3387c1a8741++) begin
         $display("I8d777f385d3dfec8815d20f7496026dc  y_nr_in [%0d]:%0d I8d1e6fa299262b2bef3b696c48864ad9[%0d]:%0d", I865c0c0b4ab0e063e5caa3387c1a8741,y_nr_in [I865c0c0b4ab0e063e5caa3387c1a8741],I865c0c0b4ab0e063e5caa3387c1a8741,I8d1e6fa299262b2bef3b696c48864ad9[I865c0c0b4ab0e063e5caa3387c1a8741]);
     end
     for (int I865c0c0b4ab0e063e5caa3387c1a8741=NN-MM;I865c0c0b4ab0e063e5caa3387c1a8741<NN;I865c0c0b4ab0e063e5caa3387c1a8741++) begin
         $display("Iaabadcf006405a774607e6b0bf567558  I8d1e6fa299262b2bef3b696c48864ad9 [%0d]:%0d", I865c0c0b4ab0e063e5caa3387c1a8741,I8d1e6fa299262b2bef3b696c48864ad9 [I865c0c0b4ab0e063e5caa3387c1a8741]);
     end
     //if (~valid_cword)
     //     $fatal (0,"Ideacadfc0571c0d4ce5104ae300edbaf I0ba4439ee9a46d9d9f14c60f88f45f87 I724a00e315992b82d662231ea0dcbe50 not a valid Ic13367945d5d4c91047b3b50234aa7ab Ic47d187067c6cf953245f128b5fde62a");
     //else
     //     $info ("Ia2a551a6458a8de22446cc76d639a9e9 a valid Ic13367945d5d4c91047b3b50234aa7ab Ic47d187067c6cf953245f128b5fde62a");

       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 0, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[0] = I8d1e6fa299262b2bef3b696c48864ad9[0] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 1, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[1] = I8d1e6fa299262b2bef3b696c48864ad9[1] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 2, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[2] = I8d1e6fa299262b2bef3b696c48864ad9[2] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 3, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[3] = I8d1e6fa299262b2bef3b696c48864ad9[3] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 4, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[4] = I8d1e6fa299262b2bef3b696c48864ad9[4] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 5, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[5] = I8d1e6fa299262b2bef3b696c48864ad9[5] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 6, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[6] = I8d1e6fa299262b2bef3b696c48864ad9[6] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 7, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[7] = I8d1e6fa299262b2bef3b696c48864ad9[7] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 8, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[8] = I8d1e6fa299262b2bef3b696c48864ad9[8] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 9, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[9] = I8d1e6fa299262b2bef3b696c48864ad9[9] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 10, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[10] = I8d1e6fa299262b2bef3b696c48864ad9[10] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 11, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[11] = I8d1e6fa299262b2bef3b696c48864ad9[11] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 12, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[12] = I8d1e6fa299262b2bef3b696c48864ad9[12] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 13, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[13] = I8d1e6fa299262b2bef3b696c48864ad9[13] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 14, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[14] = I8d1e6fa299262b2bef3b696c48864ad9[14] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 15, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[15] = I8d1e6fa299262b2bef3b696c48864ad9[15] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 16, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[16] = I8d1e6fa299262b2bef3b696c48864ad9[16] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 17, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[17] = I8d1e6fa299262b2bef3b696c48864ad9[17] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 18, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[18] = I8d1e6fa299262b2bef3b696c48864ad9[18] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 19, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[19] = I8d1e6fa299262b2bef3b696c48864ad9[19] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 20, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[20] = I8d1e6fa299262b2bef3b696c48864ad9[20] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 21, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[21] = I8d1e6fa299262b2bef3b696c48864ad9[21] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 22, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[22] = I8d1e6fa299262b2bef3b696c48864ad9[22] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 23, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[23] = I8d1e6fa299262b2bef3b696c48864ad9[23] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 24, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[24] = I8d1e6fa299262b2bef3b696c48864ad9[24] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 25, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[25] = I8d1e6fa299262b2bef3b696c48864ad9[25] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 26, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[26] = I8d1e6fa299262b2bef3b696c48864ad9[26] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 27, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[27] = I8d1e6fa299262b2bef3b696c48864ad9[27] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 28, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[28] = I8d1e6fa299262b2bef3b696c48864ad9[28] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 29, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[29] = I8d1e6fa299262b2bef3b696c48864ad9[29] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 30, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[30] = I8d1e6fa299262b2bef3b696c48864ad9[30] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 31, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[31] = I8d1e6fa299262b2bef3b696c48864ad9[31] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 32, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[32] = I8d1e6fa299262b2bef3b696c48864ad9[32] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 33, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[33] = I8d1e6fa299262b2bef3b696c48864ad9[33] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 34, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[34] = I8d1e6fa299262b2bef3b696c48864ad9[34] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 35, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[35] = I8d1e6fa299262b2bef3b696c48864ad9[35] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 36, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[36] = I8d1e6fa299262b2bef3b696c48864ad9[36] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 37, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[37] = I8d1e6fa299262b2bef3b696c48864ad9[37] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 38, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[38] = I8d1e6fa299262b2bef3b696c48864ad9[38] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 39, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[39] = I8d1e6fa299262b2bef3b696c48864ad9[39] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 40, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[40] = I8d1e6fa299262b2bef3b696c48864ad9[40] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 41, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[41] = I8d1e6fa299262b2bef3b696c48864ad9[41] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 42, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[42] = I8d1e6fa299262b2bef3b696c48864ad9[42] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 43, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[43] = I8d1e6fa299262b2bef3b696c48864ad9[43] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 44, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[44] = I8d1e6fa299262b2bef3b696c48864ad9[44] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 45, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[45] = I8d1e6fa299262b2bef3b696c48864ad9[45] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 46, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[46] = I8d1e6fa299262b2bef3b696c48864ad9[46] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 47, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[47] = I8d1e6fa299262b2bef3b696c48864ad9[47] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 48, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[48] = I8d1e6fa299262b2bef3b696c48864ad9[48] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 49, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[49] = I8d1e6fa299262b2bef3b696c48864ad9[49] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 50, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[50] = I8d1e6fa299262b2bef3b696c48864ad9[50] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 51, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[51] = I8d1e6fa299262b2bef3b696c48864ad9[51] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 52, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[52] = I8d1e6fa299262b2bef3b696c48864ad9[52] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 53, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[53] = I8d1e6fa299262b2bef3b696c48864ad9[53] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 54, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[54] = I8d1e6fa299262b2bef3b696c48864ad9[54] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 55, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[55] = I8d1e6fa299262b2bef3b696c48864ad9[55] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 56, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[56] = I8d1e6fa299262b2bef3b696c48864ad9[56] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 57, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[57] = I8d1e6fa299262b2bef3b696c48864ad9[57] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 58, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[58] = I8d1e6fa299262b2bef3b696c48864ad9[58] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 59, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[59] = I8d1e6fa299262b2bef3b696c48864ad9[59] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 60, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[60] = I8d1e6fa299262b2bef3b696c48864ad9[60] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 61, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[61] = I8d1e6fa299262b2bef3b696c48864ad9[61] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 62, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[62] = I8d1e6fa299262b2bef3b696c48864ad9[62] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 63, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[63] = I8d1e6fa299262b2bef3b696c48864ad9[63] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 64, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[64] = I8d1e6fa299262b2bef3b696c48864ad9[64] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 65, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[65] = I8d1e6fa299262b2bef3b696c48864ad9[65] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 66, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[66] = I8d1e6fa299262b2bef3b696c48864ad9[66] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 67, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[67] = I8d1e6fa299262b2bef3b696c48864ad9[67] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 68, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[68] = I8d1e6fa299262b2bef3b696c48864ad9[68] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 69, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[69] = I8d1e6fa299262b2bef3b696c48864ad9[69] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 70, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[70] = I8d1e6fa299262b2bef3b696c48864ad9[70] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 71, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[71] = I8d1e6fa299262b2bef3b696c48864ad9[71] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 72, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[72] = I8d1e6fa299262b2bef3b696c48864ad9[72] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 73, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[73] = I8d1e6fa299262b2bef3b696c48864ad9[73] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 74, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[74] = I8d1e6fa299262b2bef3b696c48864ad9[74] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 75, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[75] = I8d1e6fa299262b2bef3b696c48864ad9[75] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 76, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[76] = I8d1e6fa299262b2bef3b696c48864ad9[76] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 77, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[77] = I8d1e6fa299262b2bef3b696c48864ad9[77] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 78, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[78] = I8d1e6fa299262b2bef3b696c48864ad9[78] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 79, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[79] = I8d1e6fa299262b2bef3b696c48864ad9[79] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 80, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[80] = I8d1e6fa299262b2bef3b696c48864ad9[80] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 81, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[81] = I8d1e6fa299262b2bef3b696c48864ad9[81] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 82, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[82] = I8d1e6fa299262b2bef3b696c48864ad9[82] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 83, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[83] = I8d1e6fa299262b2bef3b696c48864ad9[83] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 84, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[84] = I8d1e6fa299262b2bef3b696c48864ad9[84] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 85, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[85] = I8d1e6fa299262b2bef3b696c48864ad9[85] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 86, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[86] = I8d1e6fa299262b2bef3b696c48864ad9[86] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 87, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[87] = I8d1e6fa299262b2bef3b696c48864ad9[87] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 88, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[88] = I8d1e6fa299262b2bef3b696c48864ad9[88] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 89, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[89] = I8d1e6fa299262b2bef3b696c48864ad9[89] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 90, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[90] = I8d1e6fa299262b2bef3b696c48864ad9[90] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 91, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[91] = I8d1e6fa299262b2bef3b696c48864ad9[91] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 92, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[92] = I8d1e6fa299262b2bef3b696c48864ad9[92] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 93, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[93] = I8d1e6fa299262b2bef3b696c48864ad9[93] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 94, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[94] = I8d1e6fa299262b2bef3b696c48864ad9[94] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 95, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[95] = I8d1e6fa299262b2bef3b696c48864ad9[95] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 96, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[96] = I8d1e6fa299262b2bef3b696c48864ad9[96] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 97, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[97] = I8d1e6fa299262b2bef3b696c48864ad9[97] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 98, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[98] = I8d1e6fa299262b2bef3b696c48864ad9[98] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 99, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[99] = I8d1e6fa299262b2bef3b696c48864ad9[99] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 100, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[100] = I8d1e6fa299262b2bef3b696c48864ad9[100] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 101, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[101] = I8d1e6fa299262b2bef3b696c48864ad9[101] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 102, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[102] = I8d1e6fa299262b2bef3b696c48864ad9[102] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 103, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[103] = I8d1e6fa299262b2bef3b696c48864ad9[103] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 104, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[104] = I8d1e6fa299262b2bef3b696c48864ad9[104] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 105, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[105] = I8d1e6fa299262b2bef3b696c48864ad9[105] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 106, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[106] = I8d1e6fa299262b2bef3b696c48864ad9[106] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 107, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[107] = I8d1e6fa299262b2bef3b696c48864ad9[107] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 108, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[108] = I8d1e6fa299262b2bef3b696c48864ad9[108] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 109, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[109] = I8d1e6fa299262b2bef3b696c48864ad9[109] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 110, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[110] = I8d1e6fa299262b2bef3b696c48864ad9[110] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 111, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[111] = I8d1e6fa299262b2bef3b696c48864ad9[111] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 112, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[112] = I8d1e6fa299262b2bef3b696c48864ad9[112] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 113, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[113] = I8d1e6fa299262b2bef3b696c48864ad9[113] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 114, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[114] = I8d1e6fa299262b2bef3b696c48864ad9[114] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 115, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[115] = I8d1e6fa299262b2bef3b696c48864ad9[115] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 116, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[116] = I8d1e6fa299262b2bef3b696c48864ad9[116] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 117, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[117] = I8d1e6fa299262b2bef3b696c48864ad9[117] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 118, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[118] = I8d1e6fa299262b2bef3b696c48864ad9[118] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 119, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[119] = I8d1e6fa299262b2bef3b696c48864ad9[119] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 120, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[120] = I8d1e6fa299262b2bef3b696c48864ad9[120] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 121, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[121] = I8d1e6fa299262b2bef3b696c48864ad9[121] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 122, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[122] = I8d1e6fa299262b2bef3b696c48864ad9[122] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 123, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[123] = I8d1e6fa299262b2bef3b696c48864ad9[123] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 124, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[124] = I8d1e6fa299262b2bef3b696c48864ad9[124] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 125, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[125] = I8d1e6fa299262b2bef3b696c48864ad9[125] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 126, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[126] = I8d1e6fa299262b2bef3b696c48864ad9[126] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 127, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[127] = I8d1e6fa299262b2bef3b696c48864ad9[127] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 128, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[128] = I8d1e6fa299262b2bef3b696c48864ad9[128] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 129, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[129] = I8d1e6fa299262b2bef3b696c48864ad9[129] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 130, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[130] = I8d1e6fa299262b2bef3b696c48864ad9[130] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 131, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[131] = I8d1e6fa299262b2bef3b696c48864ad9[131] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 132, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[132] = I8d1e6fa299262b2bef3b696c48864ad9[132] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 133, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[133] = I8d1e6fa299262b2bef3b696c48864ad9[133] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 134, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[134] = I8d1e6fa299262b2bef3b696c48864ad9[134] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 135, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[135] = I8d1e6fa299262b2bef3b696c48864ad9[135] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 136, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[136] = I8d1e6fa299262b2bef3b696c48864ad9[136] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 137, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[137] = I8d1e6fa299262b2bef3b696c48864ad9[137] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 138, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[138] = I8d1e6fa299262b2bef3b696c48864ad9[138] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 139, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[139] = I8d1e6fa299262b2bef3b696c48864ad9[139] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 140, 1,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[140] = I8d1e6fa299262b2bef3b696c48864ad9[140] ^ 1; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 141, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[141] = I8d1e6fa299262b2bef3b696c48864ad9[141] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 142, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[142] = I8d1e6fa299262b2bef3b696c48864ad9[142] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 143, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[143] = I8d1e6fa299262b2bef3b696c48864ad9[143] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 144, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[144] = I8d1e6fa299262b2bef3b696c48864ad9[144] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 145, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[145] = I8d1e6fa299262b2bef3b696c48864ad9[145] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 146, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[146] = I8d1e6fa299262b2bef3b696c48864ad9[146] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 147, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[147] = I8d1e6fa299262b2bef3b696c48864ad9[147] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 148, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[148] = I8d1e6fa299262b2bef3b696c48864ad9[148] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 149, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[149] = I8d1e6fa299262b2bef3b696c48864ad9[149] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 150, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[150] = I8d1e6fa299262b2bef3b696c48864ad9[150] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 151, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[151] = I8d1e6fa299262b2bef3b696c48864ad9[151] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 152, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[152] = I8d1e6fa299262b2bef3b696c48864ad9[152] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 153, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[153] = I8d1e6fa299262b2bef3b696c48864ad9[153] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 154, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[154] = I8d1e6fa299262b2bef3b696c48864ad9[154] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 155, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[155] = I8d1e6fa299262b2bef3b696c48864ad9[155] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 156, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[156] = I8d1e6fa299262b2bef3b696c48864ad9[156] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 157, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[157] = I8d1e6fa299262b2bef3b696c48864ad9[157] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 158, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[158] = I8d1e6fa299262b2bef3b696c48864ad9[158] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 159, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[159] = I8d1e6fa299262b2bef3b696c48864ad9[159] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 160, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[160] = I8d1e6fa299262b2bef3b696c48864ad9[160] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 161, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[161] = I8d1e6fa299262b2bef3b696c48864ad9[161] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 162, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[162] = I8d1e6fa299262b2bef3b696c48864ad9[162] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 163, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[163] = I8d1e6fa299262b2bef3b696c48864ad9[163] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 164, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[164] = I8d1e6fa299262b2bef3b696c48864ad9[164] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 165, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[165] = I8d1e6fa299262b2bef3b696c48864ad9[165] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 166, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[166] = I8d1e6fa299262b2bef3b696c48864ad9[166] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 167, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[167] = I8d1e6fa299262b2bef3b696c48864ad9[167] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 168, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[168] = I8d1e6fa299262b2bef3b696c48864ad9[168] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 169, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[169] = I8d1e6fa299262b2bef3b696c48864ad9[169] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 170, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[170] = I8d1e6fa299262b2bef3b696c48864ad9[170] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 171, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[171] = I8d1e6fa299262b2bef3b696c48864ad9[171] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 172, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[172] = I8d1e6fa299262b2bef3b696c48864ad9[172] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 173, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[173] = I8d1e6fa299262b2bef3b696c48864ad9[173] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 174, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[174] = I8d1e6fa299262b2bef3b696c48864ad9[174] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 175, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[175] = I8d1e6fa299262b2bef3b696c48864ad9[175] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 176, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[176] = I8d1e6fa299262b2bef3b696c48864ad9[176] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 177, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[177] = I8d1e6fa299262b2bef3b696c48864ad9[177] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 178, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[178] = I8d1e6fa299262b2bef3b696c48864ad9[178] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 179, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[179] = I8d1e6fa299262b2bef3b696c48864ad9[179] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 180, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[180] = I8d1e6fa299262b2bef3b696c48864ad9[180] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 181, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[181] = I8d1e6fa299262b2bef3b696c48864ad9[181] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 182, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[182] = I8d1e6fa299262b2bef3b696c48864ad9[182] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 183, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[183] = I8d1e6fa299262b2bef3b696c48864ad9[183] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 184, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[184] = I8d1e6fa299262b2bef3b696c48864ad9[184] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 185, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[185] = I8d1e6fa299262b2bef3b696c48864ad9[185] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 186, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[186] = I8d1e6fa299262b2bef3b696c48864ad9[186] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 187, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[187] = I8d1e6fa299262b2bef3b696c48864ad9[187] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 188, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[188] = I8d1e6fa299262b2bef3b696c48864ad9[188] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 189, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[189] = I8d1e6fa299262b2bef3b696c48864ad9[189] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 190, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[190] = I8d1e6fa299262b2bef3b696c48864ad9[190] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 191, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[191] = I8d1e6fa299262b2bef3b696c48864ad9[191] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 192, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[192] = I8d1e6fa299262b2bef3b696c48864ad9[192] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 193, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[193] = I8d1e6fa299262b2bef3b696c48864ad9[193] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 194, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[194] = I8d1e6fa299262b2bef3b696c48864ad9[194] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 195, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[195] = I8d1e6fa299262b2bef3b696c48864ad9[195] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 196, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[196] = I8d1e6fa299262b2bef3b696c48864ad9[196] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 197, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[197] = I8d1e6fa299262b2bef3b696c48864ad9[197] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 198, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[198] = I8d1e6fa299262b2bef3b696c48864ad9[198] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 199, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[199] = I8d1e6fa299262b2bef3b696c48864ad9[199] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 200, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[200] = I8d1e6fa299262b2bef3b696c48864ad9[200] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 201, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[201] = I8d1e6fa299262b2bef3b696c48864ad9[201] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 202, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[202] = I8d1e6fa299262b2bef3b696c48864ad9[202] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 203, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[203] = I8d1e6fa299262b2bef3b696c48864ad9[203] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 204, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[204] = I8d1e6fa299262b2bef3b696c48864ad9[204] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 205, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[205] = I8d1e6fa299262b2bef3b696c48864ad9[205] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 206, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[206] = I8d1e6fa299262b2bef3b696c48864ad9[206] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
       $display ("Icb5e100e5a9a3e7f6d1fd97512215282 bit [%0d]:%0d I83a7411fde733c403108d6608a156e2c:%0d", 207, 0,Ie18a4d4830028f90f158755e5e80fec5);
       I81dab9b4f78627240b44ac785b16acf9[207] = I8d1e6fa299262b2bef3b696c48864ad9[207] ^ 0; //Icb5e100e5a9a3e7f6d1fd97512215282 I350e6018b5636ab1e90720fed9694ccf
       Ie18a4d4830028f90f158755e5e80fec5++;
         tmp_bit[0] = 1;
         tmp_bit[1] = 1;
         tmp_bit[2] = 0;
         tmp_bit[3] = 1;
         tmp_bit[4] = 0;
         tmp_bit[5] = 0;
         tmp_bit[6] = 0;
         tmp_bit[7] = 0;
         tmp_bit[8] = 0;
         tmp_bit[9] = 1;
         tmp_bit[10] = 1;
         tmp_bit[11] = 1;
         tmp_bit[12] = 1;
         tmp_bit[13] = 1;
         tmp_bit[14] = 0;
         tmp_bit[15] = 1;
         tmp_bit[16] = 0;
         tmp_bit[17] = 0;
         tmp_bit[18] = 1;
         tmp_bit[19] = 0;
         tmp_bit[20] = 1;
         tmp_bit[21] = 1;
         tmp_bit[22] = 0;
         tmp_bit[23] = 0;
         tmp_bit[24] = 0;
         tmp_bit[25] = 1;
         tmp_bit[26] = 1;
         tmp_bit[27] = 0;
         tmp_bit[28] = 0;
         tmp_bit[29] = 1;
         tmp_bit[30] = 1;
         tmp_bit[31] = 1;
         tmp_bit[32] = 0;
         tmp_bit[33] = 0;
         tmp_bit[34] = 1;
         tmp_bit[35] = 0;
         tmp_bit[36] = 0;
         tmp_bit[37] = 0;
         tmp_bit[38] = 0;
         tmp_bit[39] = 0;
         tmp_bit[40] = 1;
         tmp_bit[41] = 0;
         tmp_bit[42] = 0;
         tmp_bit[43] = 1;
         tmp_bit[44] = 1;
         tmp_bit[45] = 1;
         tmp_bit[46] = 1;
         tmp_bit[47] = 0;
         tmp_bit[48] = 0;
         tmp_bit[49] = 1;
         tmp_bit[50] = 1;
         tmp_bit[51] = 0;
         tmp_bit[52] = 1;
         tmp_bit[53] = 1;
         tmp_bit[54] = 0;
         tmp_bit[55] = 1;
         tmp_bit[56] = 1;
         tmp_bit[57] = 0;
         tmp_bit[58] = 0;
         tmp_bit[59] = 1;
         tmp_bit[60] = 0;
         tmp_bit[61] = 0;
         tmp_bit[62] = 0;
         tmp_bit[63] = 1;
         tmp_bit[64] = 0;
         tmp_bit[65] = 1;
         tmp_bit[66] = 1;
         tmp_bit[67] = 1;
         tmp_bit[68] = 1;
         tmp_bit[69] = 1;
         tmp_bit[70] = 1;
         tmp_bit[71] = 1;
         tmp_bit[72] = 0;
         tmp_bit[73] = 0;
         tmp_bit[74] = 1;
         tmp_bit[75] = 0;
         tmp_bit[76] = 0;
         tmp_bit[77] = 0;
         tmp_bit[78] = 0;
         tmp_bit[79] = 0;
         tmp_bit[80] = 0;
         tmp_bit[81] = 1;
         tmp_bit[82] = 1;
         tmp_bit[83] = 0;
         tmp_bit[84] = 0;
         tmp_bit[85] = 0;
         tmp_bit[86] = 0;
         tmp_bit[87] = 0;
         tmp_bit[88] = 0;
         tmp_bit[89] = 1;
         tmp_bit[90] = 0;
         tmp_bit[91] = 1;
         tmp_bit[92] = 0;
         tmp_bit[93] = 0;
         tmp_bit[94] = 0;
         tmp_bit[95] = 0;
         tmp_bit[96] = 0;
         tmp_bit[97] = 0;
         tmp_bit[98] = 0;
         tmp_bit[99] = 0;
         tmp_bit[100] = 1;
         tmp_bit[101] = 1;
         tmp_bit[102] = 1;
         tmp_bit[103] = 1;
         tmp_bit[104] = 0;
         tmp_bit[105] = 1;
         tmp_bit[106] = 1;
         tmp_bit[107] = 1;
         tmp_bit[108] = 0;
         tmp_bit[109] = 0;
         tmp_bit[110] = 0;
         tmp_bit[111] = 1;
         tmp_bit[112] = 1;
         tmp_bit[113] = 0;
         tmp_bit[114] = 0;
         tmp_bit[115] = 1;
         tmp_bit[116] = 1;
         tmp_bit[117] = 1;
         tmp_bit[118] = 1;
         tmp_bit[119] = 0;
         tmp_bit[120] = 1;
         tmp_bit[121] = 0;
         tmp_bit[122] = 0;
         tmp_bit[123] = 1;
         tmp_bit[124] = 0;
         tmp_bit[125] = 0;
         tmp_bit[126] = 1;
         tmp_bit[127] = 1;
         tmp_bit[128] = 1;
         tmp_bit[129] = 0;
         tmp_bit[130] = 1;
         tmp_bit[131] = 0;
         tmp_bit[132] = 0;
         tmp_bit[133] = 0;
         tmp_bit[134] = 1;
         tmp_bit[135] = 1;
         tmp_bit[136] = 1;
         tmp_bit[137] = 0;
         tmp_bit[138] = 1;
         tmp_bit[139] = 1;
         tmp_bit[140] = 1;
         tmp_bit[141] = 0;
         tmp_bit[142] = 0;
         tmp_bit[143] = 1;
         tmp_bit[144] = 0;
         tmp_bit[145] = 1;
         tmp_bit[146] = 0;
         tmp_bit[147] = 1;
         tmp_bit[148] = 1;
         tmp_bit[149] = 1;
         tmp_bit[150] = 1;
         tmp_bit[151] = 0;
         tmp_bit[152] = 1;
         tmp_bit[153] = 0;
         tmp_bit[154] = 0;
         tmp_bit[155] = 0;
         tmp_bit[156] = 0;
         tmp_bit[157] = 1;
         tmp_bit[158] = 0;
         tmp_bit[159] = 1;
         tmp_bit[160] = 1;
         tmp_bit[161] = 0;
         tmp_bit[162] = 0;
         tmp_bit[163] = 1;
         tmp_bit[164] = 0;
         tmp_bit[165] = 0;
         tmp_bit[166] = 1;
         tmp_bit[167] = 1;
         tmp_bit[168] = 0;
         tmp_bit[169] = 0;
         tmp_bit[170] = 1;
         tmp_bit[171] = 0;
         tmp_bit[172] = 1;
         tmp_bit[173] = 1;
         tmp_bit[174] = 0;
         tmp_bit[175] = 0;
         tmp_bit[176] = 1;
         tmp_bit[177] = 0;
         tmp_bit[178] = 1;
         tmp_bit[179] = 1;
         tmp_bit[180] = 1;
         tmp_bit[181] = 0;
         tmp_bit[182] = 1;
         tmp_bit[183] = 1;
         tmp_bit[184] = 1;
         tmp_bit[185] = 1;
         tmp_bit[186] = 0;
         tmp_bit[187] = 1;
         tmp_bit[188] = 0;
         tmp_bit[189] = 0;
         tmp_bit[190] = 0;
         tmp_bit[191] = 0;
         tmp_bit[192] = 1;
         tmp_bit[193] = 0;
         tmp_bit[194] = 0;
         tmp_bit[195] = 0;
         tmp_bit[196] = 0;
         tmp_bit[197] = 0;
         tmp_bit[198] = 0;
         tmp_bit[199] = 0;
         tmp_bit[200] = 0;
         tmp_bit[201] = 0;
         tmp_bit[202] = 1;
         tmp_bit[203] = 0;
         tmp_bit[204] = 0;
         tmp_bit[205] = 0;
         tmp_bit[206] = 1;
         tmp_bit[207] = 0;
     repeat (1) @ (posedge clk);
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[0] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 0, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 0, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[1] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 1, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 1, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[2] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 2, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 2, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[3] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 3, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 3, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[4] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 4, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 4, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[5] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 5, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 5, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[6] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 6, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 6, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[7] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 7, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 7, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[8] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 8, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 8, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[9] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 9, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 9, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[10] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 10, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 10, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[11] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 11, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 11, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[12] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 12, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 12, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[13] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 13, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 13, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[14] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 14, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 14, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[15] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 15, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 15, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[16] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 16, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 16, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[17] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 17, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 17, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[18] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 18, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 18, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[19] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 19, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 19, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[20] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 20, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 20, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[21] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 21, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 21, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[22] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 22, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 22, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[23] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 23, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 23, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[24] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 24, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 24, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[25] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 25, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 25, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[26] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 26, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 26, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[27] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 27, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 27, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[28] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 28, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 28, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[29] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 29, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 29, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[30] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 30, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 30, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[31] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 31, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 31, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[32] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 32, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 32, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[33] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 33, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 33, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[34] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 34, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 34, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[35] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 35, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 35, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[36] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 36, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 36, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[37] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 37, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 37, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[38] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 38, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 38, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[39] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 39, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 39, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[40] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 40, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 40, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[41] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 41, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 41, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[42] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 42, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 42, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[43] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 43, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 43, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[44] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 44, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 44, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[45] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 45, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 45, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[46] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 46, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 46, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[47] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 47, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 47, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[48] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 48, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 48, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[49] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 49, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 49, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[50] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 50, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 50, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[51] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 51, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 51, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[52] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 52, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 52, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[53] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 53, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 53, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[54] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 54, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 54, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[55] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 55, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 55, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[56] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 56, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 56, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[57] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 57, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 57, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[58] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 58, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 58, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[59] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 59, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 59, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[60] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 60, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 60, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[61] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 61, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 61, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[62] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 62, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 62, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[63] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 63, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 63, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[64] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 64, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 64, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[65] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 65, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 65, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[66] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 66, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 66, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[67] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 67, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 67, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[68] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 68, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 68, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[69] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 69, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 69, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[70] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 70, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 70, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[71] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 71, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 71, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[72] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 72, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 72, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[73] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 73, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 73, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[74] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 74, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 74, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[75] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 75, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 75, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[76] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 76, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 76, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[77] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 77, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 77, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[78] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 78, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 78, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[79] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 79, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 79, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[80] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 80, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 80, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[81] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 81, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 81, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[82] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 82, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 82, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[83] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 83, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 83, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[84] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 84, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 84, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[85] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 85, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 85, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[86] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 86, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 86, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[87] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 87, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 87, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[88] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 88, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 88, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[89] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 89, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 89, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[90] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 90, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 90, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[91] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 91, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 91, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[92] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 92, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 92, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[93] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 93, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 93, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[94] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 94, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 94, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[95] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 95, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 95, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[96] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 96, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 96, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[97] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 97, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 97, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[98] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 98, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 98, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[99] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 99, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 99, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[100] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 100, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 100, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[101] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 101, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 101, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[102] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 102, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 102, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[103] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 103, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 103, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[104] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 104, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 104, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[105] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 105, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 105, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[106] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 106, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 106, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[107] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 107, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 107, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[108] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 108, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 108, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[109] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 109, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 109, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[110] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 110, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 110, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[111] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 111, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 111, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[112] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 112, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 112, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[113] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 113, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 113, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[114] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 114, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 114, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[115] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 115, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 115, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[116] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 116, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 116, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[117] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 117, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 117, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[118] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 118, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 118, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[119] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 119, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 119, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[120] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 120, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 120, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[121] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 121, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 121, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[122] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 122, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 122, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[123] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 123, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 123, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[124] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 124, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 124, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[125] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 125, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 125, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[126] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 126, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 126, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[127] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 127, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 127, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[128] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 128, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 128, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[129] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 129, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 129, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[130] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 130, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 130, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[131] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 131, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 131, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[132] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 132, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 132, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[133] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 133, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 133, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[134] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 134, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 134, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[135] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 135, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 135, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[136] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 136, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 136, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[137] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 137, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 137, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[138] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 138, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 138, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[139] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 139, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 139, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[140] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 140, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 140, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[141] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 141, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 141, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[142] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 142, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 142, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[143] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 143, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 143, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[144] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 144, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 144, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[145] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 145, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 145, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[146] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 146, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 146, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[147] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 147, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 147, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[148] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 148, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 148, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[149] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 149, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 149, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[150] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 150, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 150, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[151] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 151, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 151, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[152] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 152, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 152, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[153] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 153, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 153, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[154] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 154, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 154, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[155] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 155, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 155, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[156] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 156, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 156, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[157] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 157, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 157, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[158] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 158, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 158, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[159] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 159, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 159, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[160] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 160, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 160, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[161] ;
         if ( 1 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 161, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",1, 161, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[162] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 162, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 162, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[163] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 163, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 163, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[164] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 164, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 164, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[165] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 165, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 165, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[166] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 166, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 166, I798dd71209184f626a7f6bed517aa125 );
         end
         I798dd71209184f626a7f6bed517aa125 = ~  syndrome[167] ;
         if ( 0 == I798dd71209184f626a7f6bed517aa125 ) begin
              $display ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 167, I798dd71209184f626a7f6bed517aa125 );
         end else begin
              $error   ("syndrome Iebc6097498b06421e2759a773c992ed3:%0d syndrome[%0d]:%0d",0, 167, I798dd71209184f626a7f6bed517aa125 );
         end
     repeat (1) @ (posedge clk);
     $finish;

     for (int I865c0c0b4ab0e063e5caa3387c1a8741=0;I865c0c0b4ab0e063e5caa3387c1a8741<NN;I865c0c0b4ab0e063e5caa3387c1a8741++) begin
            if (I81dab9b4f78627240b44ac785b16acf9[I865c0c0b4ab0e063e5caa3387c1a8741]) begin
                 I61e23fc401e882840b471b3b125a68a9  [I865c0c0b4ab0e063e5caa3387c1a8741] <= 2'b11;  // Icfd8f331d281b0da79e7c6ed6988243c 1: -1 === 2'b11
                                    // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 1 If44b5337a5f63ffc29f578e9a8c52b9b -1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b11
            end else begin
                 I61e23fc401e882840b471b3b125a68a9  [I865c0c0b4ab0e063e5caa3387c1a8741] <= 2'b01;  // Icfd8f331d281b0da79e7c6ed6988243c 0: 1  === 2'b01
                                    // I2063c1608d6e0baf80249c42e2be5804 I8bf8854bebe108183caeb845c7676ae4 0 If44b5337a5f63ffc29f578e9a8c52b9b 1 I13b5bfe96f3e2fe411c9f66f4a582adf Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 2'b01
            end
     end
     for (int I865c0c0b4ab0e063e5caa3387c1a8741=0;I865c0c0b4ab0e063e5caa3387c1a8741<MM;I865c0c0b4ab0e063e5caa3387c1a8741++) begin
         exp_syn [I865c0c0b4ab0e063e5caa3387c1a8741] <= 1'b1;
     end

  end




  repeat (4) @ (posedge clk);
  Iea2b2676c28c0db26d39331a336c6b92                          <= 1'b1;
  repeat (1) @ (posedge clk);
  Iea2b2676c28c0db26d39331a336c6b92                          <= 1'b0;
  repeat (20) @(posedge clk);
  $display("I4f62dc0a0e700849a9987d10e9dc369b:Ib3508db383796b91f1628675de826704 I4f33252742282f871b0617168156fd55 I90272dda245ae1fb3cf197e91a8689dc :%0d %t", Ifb48ed869c44bdc930da7ccc778d5014, $time);
  repeat (20) @(posedge clk);
  $finish();
end


assign percent_probability_int = 32'd 206;

initial
begin
`ifdef IVERILOG
          $dumpfile("sntc_ldpc_syndrome_tb.I935c34f94bcb203a6a5a2255c3cebffa");
          $dumpvars(0, sntc_ldpc_syndrome_tb);
`endif
  repeat (600) @(posedge clk);
end

initial
begin
  forever begin
      if (I7de33615d7fbc1cb7bc608d12f1993d2[1]) begin
         $display("Iba06facad762a0a1ec4f0d5bf31b6b3d end If910ff3a8628ebda9c67ed678703fd7d");
         if (I7de33615d7fbc1cb7bc608d12f1993d2[0]) begin
            $display("I269f3d1562cbd15624e7d2c4b10122e3: I74cac558072300385f7ab4dff7465e3c If00bbb7747929fafa9d1afd071dba78e");
         end else begin
            $error("Ib9e14d9b2886bcff408b85aefa780419: I74cac558072300385f7ab4dff7465e3c not If00bbb7747929fafa9d1afd071dba78e");
         end
         $finish();
      end
      repeat (1) @(posedge clk);
  end
end

`endif




`ifdef ENCRYPT
`endif

endmodule

//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.100000 I7290d6b1f1458098d2f225877e609ba6:2.197225 percent_probability_int:'d141

 //Ic07b0b4d7660314f711a68fc47c4ab38 I48d8d6f5a3efbf52837d6b788a22859a valid Ic13367945d5d4c91047b3b50234aa7ab Ic47d187067c6cf953245f128b5fde62a
//y_int:
 //44010bdd34c9a17a9dc5c9798ef00a0604fe89b67904e634be0b
//Iebc6097498b06421e2759a773c992ed3:
 //0200400200100008100880c0000680200320002200
//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.038462 I7290d6b1f1458098d2f225877e609ba6:3.218876 percent_probability_int:'d206
