 reg  ['h3ff:0] [$clog2('h7000+1)-1:0] Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441 ;
