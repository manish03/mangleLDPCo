 parameter flogtanh_WDTH =  20 ;
 reg  [flogtanh_WDTH -1 :0] flogtanh_sel ;
 reg  [$clog2('h7000+1)-1:0] I0ef7780b478bfb05e8c9bf2fcea00183 ;
