//`include "GF2_LDPC_fgallag_0x00012_assign_inc.sv"
//always_comb begin
              I6be0bfc1327465230710d1b067b706d4['h00000] = 
          (!fgallag_sel['h00012]) ? 
                       I34f69b29975fc71eeee92e6ac4210723['h00000] : //%
                       I34f69b29975fc71eeee92e6ac4210723['h00001] ;
//end
