              I5615abbd072d30da52163f16f1980957 = 
          (!flogtanh_sel[4]) ? 
                       I869ad51812ced1ce31815a7ccaf5578d: 
                       I6442979212fb9e03df3685a28065f02e;
              Ie7e694e2f86689b06efbd2eb66c5ffd8 = 
          (!flogtanh_sel[4]) ? 
                       I5e2d92b7f01402ec98771a9026c756e5: 
                       I3050b73b4bf3bb60e38178a3a372231f;
              Id0287bb263a65d5eea34cbd5be2cfe3d = 
          (!flogtanh_sel[4]) ? 
                       I32f1d36a7d8d44da0bc6d3ad8d2a1153: 
                       I7637d7cc7dc2189e17cce002a981082a;
              Ic223bac65f3241d30afc2e21178eebfc = 
          (!flogtanh_sel[4]) ? 
                       I0cb1cf10cb15dd8c1066f460f67538c2: 
                       Ifbe06c2706fb89aaa251789703159e25;
              I22794d7d1503d8cf477ad8b189d53ace = 
          (!flogtanh_sel[4]) ? 
                       I8fe4558357f35c3e71ab801b22392c83: 
                       Ic6a2f31a403a6389f0d7df052a5cfdec;
              I8ccd9901d0629218945ab24f6eea34a3 = 
          (!flogtanh_sel[4]) ? 
                       I96b2c098a97cd3303228da6f6484e240: 
                       I9d07ffc430043e95f348f4d05d3f6dbb;
              Ifdeb82639682ca4a87f76e40a181bf79 = 
          (!flogtanh_sel[4]) ? 
                       I4cd469fecb0f25820f04091a44c50b61: 
                       Ib7fe035c4d2cc2f25edc04489db7a532;
              Ib1879574e569ce9d6787132cc87e8de4 = 
          (!flogtanh_sel[4]) ? 
                       I923a9ae3ead074bc3abd711b3378060d: 
                       I53c4fe7b76ec5282e86c2fb100bb6b18;
              Ifbb918c9c8ed9c0de0d1fd1e02eccd4d = 
          (!flogtanh_sel[4]) ? 
                       Ib1f88a9e7696e0798fbeedbbd1aaaf92: 
                       Iabe16f9be9c25cd6e4c2b63984a7e09b;
               Ib230198837d881f6349f181cf4b3c4c8 =  I606e85239115132c5e6281b7ed7ec81a ;
               I1a07a0d5e3768a4ecf4c56f6698fef63 =  I5f13934441008d491b64e006c2704a7f ;
              I55ff759485b4e816fac06d20ac5b2790 = 
          (!flogtanh_sel[4]) ? 
                       I33399cd8c4a4774d52f0ff4940f8321e: 
                       I2abe8717ff4ddfa416d7b2cb47edf15d;
