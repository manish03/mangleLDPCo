 reg  ['h1fff:0] [$clog2('h7000+1)-1:0] Ic18a6d922901eba6fa14d7b0fce00db5418ec3266b6efe12d09f4bf837920f3f ;
