//`include "GF2_LDPC_flogtanh_0x00006_assign_inc.sv"
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00000] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00000] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00001] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00001] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00002] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00003] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00002] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00004] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00005] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00003] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00006] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00007] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00004] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00008] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00009] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00005] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00006] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00007] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00008] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00010] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00011] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00009] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00012] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00013] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000a] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00014] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00015] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000b] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00016] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00017] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000c] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00018] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00019] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000d] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0000f] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00010] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00020] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00021] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00011] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00022] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00023] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00012] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00024] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00025] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00013] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00026] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00027] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00014] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00028] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00029] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00015] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00016] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00017] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00018] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00030] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00031] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00019] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00032] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00033] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001a] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00034] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00035] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001b] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00036] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00037] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001c] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00038] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00039] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001d] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0001f] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00020] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00040] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00041] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00021] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00042] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00043] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00022] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00044] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00045] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00023] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00046] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00047] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00024] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00048] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00049] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00025] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00026] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00027] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00028] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00050] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00051] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00029] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00052] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00053] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002a] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00054] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00055] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002b] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00056] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00057] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002c] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00058] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00059] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002d] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0002f] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00030] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00060] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00061] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00031] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00062] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00063] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00032] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00064] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00065] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00033] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00066] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00067] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00034] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00068] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00069] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00035] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00036] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00037] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00038] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00070] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00071] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00039] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00072] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00073] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003a] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00074] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00075] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003b] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00076] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00077] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003c] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00078] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00079] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003d] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0003f] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00040] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00080] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00081] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00041] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00082] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00083] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00042] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00084] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00085] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00043] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00086] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00087] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00044] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00088] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00089] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00045] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00046] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00047] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00048] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00090] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00091] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00049] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00092] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00093] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004a] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00094] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00095] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004b] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00096] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00097] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004c] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00098] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00099] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004d] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009a] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009b] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009c] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009d] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0004f] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009e] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009f] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00050] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a0] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a1] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00051] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a2] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a3] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00052] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a4] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a5] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00053] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a6] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a7] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00054] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a8] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a9] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00055] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000aa] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ab] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00056] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ac] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ad] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00057] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ae] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000af] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00058] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b0] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b1] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00059] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b2] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b3] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005a] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b4] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b5] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005b] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b6] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b7] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005c] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b8] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b9] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ba] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bc] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bd] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0005f] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000be] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bf] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00060] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c0] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00061] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c2] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c3] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00062] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c4] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c5] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00063] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c6] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00064] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c8] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c9] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00065] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00066] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000cc] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00067] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ce] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000cf] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00068] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d0] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00069] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d2] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d3] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d8] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006d] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000da] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000db] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0006f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00070] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e0] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00071] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e2] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e3] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00072] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00073] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00074] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00075] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ea] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00076] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ec] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ed] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00077] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00078] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00079] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fa] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007e] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fc] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fd] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0007f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00080] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00100] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00081] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00102] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00082] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00104] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00083] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00106] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00084] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00108] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00085] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00086] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00087] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00088] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00110] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00089] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00112] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00114] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00116] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00118] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0008f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011e] ;
//end
//always_comb begin
              I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00090] = 
          (!flogtanh_sel['h00006]) ? 
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00120] : //%
                       I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00121] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00091] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00122] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00092] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00124] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00093] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00126] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00094] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00128] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00095] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00096] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00097] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00098] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00130] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00099] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00132] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00134] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00136] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00138] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0009f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00140] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00142] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00144] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00146] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00148] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00150] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00152] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00154] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00156] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00158] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00160] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00162] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00164] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00166] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00168] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00170] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00172] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00174] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00176] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00178] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00180] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00182] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00184] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00186] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00188] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00190] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00192] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00194] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00196] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00198] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h000ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00100] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00200] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00101] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00202] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00102] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00204] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00103] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00206] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00104] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00208] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00105] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00106] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00107] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00108] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00210] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00109] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00212] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00214] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00216] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00218] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0010f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00110] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00220] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00111] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00222] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00112] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00224] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00113] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00226] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00114] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00228] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00115] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00116] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00117] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00118] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00230] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00119] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00232] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00234] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00236] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00238] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0011f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00120] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00240] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00121] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00242] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00122] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00244] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00123] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00246] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00124] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00248] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00125] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00126] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00127] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00128] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00250] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00129] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00252] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00254] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00256] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00258] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0012f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00130] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00260] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00131] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00262] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00132] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00264] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00133] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00266] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00134] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00268] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00135] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00136] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00137] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00138] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00270] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00139] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00272] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00274] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00276] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00278] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0013f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00140] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00280] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00141] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00282] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00142] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00284] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00143] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00286] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00144] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00288] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00145] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00146] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00147] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00148] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00290] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00149] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00292] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00294] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00296] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00298] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0014f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00150] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00151] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00152] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00153] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00154] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00155] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00156] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00157] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00158] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00159] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0015f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00160] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00161] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00162] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00163] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00164] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00165] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00166] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00167] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00168] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00169] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0016f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00170] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00171] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00172] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00173] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00174] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00175] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00176] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00177] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00178] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00179] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0017f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00180] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00300] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00181] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00302] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00182] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00304] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00183] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00306] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00184] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00308] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00185] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00186] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00187] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00188] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00310] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00189] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00312] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00314] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00316] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00318] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0018f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00190] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00320] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00191] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00322] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00192] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00324] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00193] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00326] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00194] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00328] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00195] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00196] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00197] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00198] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00330] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00199] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00332] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00334] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00336] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00338] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0019f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00340] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00342] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00344] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00346] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00348] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00350] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00352] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00354] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00356] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00358] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00360] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00362] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00364] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00366] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00368] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00370] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00372] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00374] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00376] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00378] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00380] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00382] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00384] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00386] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00388] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00390] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00392] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00394] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00396] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00398] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h001ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00200] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00400] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00201] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00402] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00202] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00404] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00203] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00406] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00204] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00408] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00205] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00206] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00207] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00208] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00410] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00209] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00412] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00414] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00416] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00418] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0020f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00210] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00420] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00211] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00422] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00212] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00424] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00213] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00426] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00214] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00428] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00215] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00216] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00217] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00218] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00430] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00219] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00432] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00434] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00436] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00438] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0021f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00220] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00440] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00221] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00442] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00222] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00444] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00223] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00446] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00224] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00448] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00225] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00226] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00227] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00228] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00450] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00229] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00452] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00454] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00456] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00458] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0022f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00230] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00460] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00231] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00462] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00232] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00464] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00233] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00466] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00234] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00468] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00235] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00236] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00237] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00238] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00470] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00239] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00472] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00474] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00476] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00478] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0023f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00240] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00480] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00241] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00482] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00242] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00484] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00243] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00486] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00244] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00488] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00245] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00246] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00247] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00248] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00490] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00249] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00492] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00494] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00496] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00498] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0024f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00250] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00251] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00252] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00253] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00254] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00255] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00256] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00257] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00258] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00259] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0025f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00260] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00261] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00262] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00263] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00264] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00265] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00266] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00267] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00268] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00269] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0026f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00270] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00271] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00272] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00273] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00274] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00275] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00276] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00277] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00278] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00279] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0027f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00280] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00500] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00281] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00502] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00282] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00504] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00283] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00506] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00284] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00508] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00285] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00286] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00287] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00288] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00510] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00289] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00512] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00514] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00516] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00518] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0028f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00290] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00520] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00291] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00522] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00292] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00524] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00293] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00526] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00294] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00528] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00295] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00296] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00297] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00298] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00530] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00299] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00532] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00534] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00536] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00538] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0029f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00540] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00542] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00544] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00546] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00548] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00550] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00552] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00554] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00556] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00558] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00560] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00562] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00564] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00566] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00568] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00570] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00572] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00574] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00576] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00578] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00580] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00582] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00584] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00586] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00588] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00590] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00592] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00594] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00596] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00598] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h002ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00300] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00600] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00301] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00602] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00302] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00604] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00303] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00606] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00304] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00608] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00305] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00306] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00307] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00308] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00610] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00309] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00612] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00614] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00616] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00618] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0030f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00310] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00620] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00311] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00622] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00312] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00624] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00313] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00626] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00314] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00628] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00315] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00316] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00317] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00318] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00630] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00319] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00632] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00634] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00636] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00638] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0031f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00320] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00640] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00321] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00642] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00322] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00644] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00323] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00646] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00324] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00648] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00325] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00326] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00327] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00328] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00650] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00329] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00652] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00654] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00656] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00658] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0032f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00330] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00660] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00331] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00662] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00332] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00664] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00333] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00666] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00334] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00668] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00335] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00336] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00337] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00338] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00670] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00339] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00672] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00674] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00676] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00678] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0033f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00340] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00680] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00341] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00682] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00342] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00684] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00343] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00686] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00344] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00688] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00345] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00346] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00347] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00348] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00690] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00349] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00692] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00694] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00696] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00698] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0034f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00350] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00351] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00352] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00353] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00354] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00355] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00356] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00357] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00358] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00359] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0035f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00360] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00361] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00362] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00363] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00364] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00365] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00366] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00367] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00368] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00369] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0036f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00370] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00371] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00372] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00373] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00374] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00375] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00376] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00377] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00378] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00379] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0037f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00380] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00700] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00381] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00702] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00382] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00704] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00383] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00706] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00384] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00708] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00385] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00386] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00387] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00388] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00710] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00389] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00712] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00714] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00716] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00718] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0038f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00390] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00720] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00391] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00722] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00392] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00724] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00393] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00726] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00394] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00728] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00395] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00396] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00397] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00398] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00730] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00399] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00732] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00734] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00736] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00738] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0039f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00740] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00742] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00744] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00746] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00748] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00750] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00752] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00754] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00756] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00758] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00760] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00762] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00764] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00766] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00768] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00770] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00772] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00774] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00776] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00778] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00780] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00782] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00784] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00786] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00788] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00790] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00792] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00794] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00796] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00798] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h003ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00400] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00800] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00401] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00802] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00402] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00804] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00403] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00806] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00404] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00808] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00405] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00406] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00407] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00408] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00810] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00409] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00812] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00814] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00816] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00818] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0040f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00410] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00820] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00411] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00822] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00412] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00824] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00413] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00826] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00414] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00828] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00415] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00416] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00417] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00418] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00830] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00419] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00832] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00834] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00836] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00838] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0041f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00420] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00840] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00421] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00842] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00422] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00844] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00423] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00846] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00424] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00848] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00425] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00426] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00427] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00428] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00850] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00429] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00852] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00854] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00856] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00858] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0042f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00430] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00860] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00431] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00862] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00432] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00864] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00433] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00866] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00434] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00868] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00435] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00436] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00437] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00438] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00870] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00439] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00872] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00874] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00876] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00878] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0043f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00440] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00880] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00441] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00882] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00442] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00884] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00443] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00886] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00444] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00888] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00445] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00446] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00447] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00448] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00890] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00449] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00892] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00894] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00896] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00898] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0044f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00450] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00451] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00452] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00453] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00454] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00455] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00456] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00457] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00458] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00459] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0045f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00460] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00461] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00462] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00463] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00464] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00465] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00466] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00467] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00468] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00469] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0046f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00470] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00471] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00472] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00473] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00474] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00475] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00476] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00477] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00478] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00479] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0047f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00480] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00900] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00481] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00902] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00482] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00904] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00483] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00906] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00484] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00908] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00485] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00486] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00487] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00488] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00910] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00489] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00912] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00914] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00916] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00918] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0048f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00490] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00920] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00491] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00922] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00492] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00924] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00493] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00926] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00494] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00928] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00495] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00496] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00497] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00498] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00930] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00499] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00932] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00934] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00936] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00938] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0049f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00940] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00942] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00944] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00946] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00948] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00950] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00952] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00954] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00956] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00958] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00960] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00962] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00964] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00966] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00968] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00970] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00972] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00974] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00976] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00978] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00980] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00982] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00984] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00986] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00988] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00990] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00992] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00994] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00996] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00998] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h004ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00500] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00501] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00502] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00503] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00504] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00505] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00506] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00507] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00508] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00509] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0050f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00510] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00511] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00512] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00513] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00514] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00515] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00516] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00517] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00518] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00519] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0051f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00520] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00521] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00522] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00523] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00524] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00525] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00526] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00527] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00528] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00529] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0052f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00530] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00531] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00532] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00533] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00534] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00535] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00536] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00537] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00538] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00539] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0053f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00540] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00541] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00542] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00543] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00544] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00545] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00546] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00547] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00548] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00549] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0054f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00550] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00551] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00552] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00553] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00554] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00555] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aaa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00556] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00557] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00558] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00559] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0055f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00560] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00561] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00562] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00563] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00564] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00565] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00566] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00acc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00567] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ace] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00568] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00569] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ada] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00adc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0056f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ade] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00570] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00571] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00572] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00573] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00574] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00575] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00576] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00577] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00578] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00579] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0057f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00580] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00581] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00582] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00583] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00584] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00585] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00586] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00587] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00588] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00589] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0058f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00590] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00591] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00592] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00593] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00594] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00595] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00596] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00597] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00598] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00599] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0059f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00baa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bcc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bdc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h005ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00600] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00601] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00602] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00603] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00604] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00605] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00606] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00607] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00608] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00609] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0060f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00610] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00611] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00612] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00613] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00614] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00615] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00616] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00617] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00618] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00619] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0061f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00620] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00621] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00622] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00623] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00624] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00625] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00626] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00627] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00628] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00629] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0062f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00630] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00631] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00632] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00633] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00634] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00635] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00636] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00637] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00638] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00639] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0063f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00640] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00641] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00642] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00643] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00644] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00645] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00646] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00647] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00648] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00649] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0064f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00650] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00651] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00652] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00653] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00654] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00655] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00caa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00656] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00657] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00658] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00659] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0065f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00660] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00661] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00662] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00663] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00664] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00665] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00666] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ccc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00667] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00668] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00669] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cdc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0066f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00670] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00671] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00672] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00673] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00674] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00675] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00676] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00677] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00678] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00679] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0067f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00680] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00681] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00682] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00683] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00684] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00685] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00686] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00687] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00688] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00689] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0068f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00690] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00691] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00692] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00693] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00694] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00695] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00696] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00697] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00698] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00699] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0069f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00daa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dcc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ddc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h006ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00700] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00701] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00702] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00703] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00704] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00705] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00706] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00707] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00708] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00709] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0070f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00710] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00711] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00712] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00713] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00714] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00715] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00716] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00717] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00718] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00719] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0071f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00720] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00721] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00722] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00723] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00724] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00725] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00726] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00727] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00728] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00729] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0072f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00730] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00731] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00732] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00733] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00734] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00735] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00736] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00737] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00738] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00739] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0073f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00740] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00741] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00742] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00743] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00744] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00745] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00746] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00747] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00748] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00749] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0074f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00750] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00751] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00752] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00753] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00754] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00755] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eaa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00756] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00757] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00758] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00759] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0075f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00760] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00761] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00762] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00763] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00764] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00765] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00766] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ecc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00767] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ece] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00768] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00769] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00edc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0076f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ede] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00770] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00771] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00772] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00773] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00774] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00775] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00776] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00777] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00778] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00779] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0077f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00780] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00781] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00782] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00783] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00784] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00785] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00786] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00787] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00788] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00789] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0078f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00790] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00791] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00792] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00793] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00794] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00795] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00796] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00797] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00798] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00799] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0079f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00faa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fcc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fdc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h007ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00800] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01000] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00801] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01002] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00802] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01004] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00803] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01006] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00804] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01008] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00805] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00806] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00807] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00808] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01010] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00809] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01012] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01014] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01016] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01018] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0080f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00810] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01020] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00811] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01022] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00812] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01024] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00813] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01026] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00814] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01028] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00815] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00816] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00817] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00818] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01030] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00819] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01032] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01034] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01036] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01038] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0081f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00820] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01040] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00821] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01042] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00822] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01044] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00823] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01046] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00824] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01048] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00825] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00826] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00827] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00828] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01050] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00829] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01052] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01054] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01056] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01058] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0082f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00830] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01060] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00831] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01062] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00832] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01064] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00833] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01066] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00834] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01068] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00835] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00836] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00837] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00838] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01070] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00839] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01072] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01074] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01076] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01078] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0083f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00840] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01080] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00841] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01082] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00842] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01084] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00843] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01086] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00844] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01088] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00845] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00846] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00847] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00848] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01090] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00849] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01092] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01094] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01096] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01098] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0084f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00850] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00851] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00852] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00853] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00854] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00855] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00856] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00857] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00858] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00859] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0085f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00860] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00861] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00862] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00863] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00864] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00865] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00866] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00867] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00868] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00869] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0086f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00870] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00871] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00872] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00873] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00874] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00875] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00876] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00877] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00878] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00879] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0087f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00880] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01100] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00881] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01102] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00882] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01104] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00883] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01106] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00884] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01108] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00885] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00886] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00887] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00888] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01110] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00889] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01112] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01114] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01116] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01118] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0088f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00890] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01120] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00891] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01122] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00892] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01124] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00893] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01126] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00894] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01128] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00895] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00896] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00897] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00898] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01130] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00899] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01132] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01134] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01136] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01138] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0089f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01140] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01142] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01144] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01146] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01148] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01150] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01152] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01154] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01156] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01158] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01160] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01162] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01164] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01166] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01168] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01170] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01172] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01174] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01176] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01178] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01180] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01182] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01184] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01186] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01188] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01190] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01192] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01194] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01196] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01198] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h008ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00900] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01200] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00901] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01202] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00902] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01204] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00903] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01206] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00904] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01208] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00905] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00906] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00907] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00908] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01210] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00909] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01212] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01214] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01216] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01218] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0090f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00910] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01220] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00911] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01222] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00912] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01224] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00913] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01226] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00914] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01228] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00915] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00916] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00917] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00918] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01230] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00919] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01232] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01234] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01236] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01238] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0091f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00920] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01240] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00921] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01242] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00922] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01244] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00923] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01246] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00924] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01248] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00925] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00926] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00927] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00928] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01250] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00929] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01252] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01254] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01256] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01258] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0092f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00930] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01260] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00931] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01262] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00932] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01264] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00933] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01266] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00934] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01268] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00935] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00936] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00937] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00938] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01270] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00939] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01272] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01274] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01276] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01278] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0093f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00940] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01280] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00941] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01282] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00942] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01284] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00943] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01286] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00944] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01288] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00945] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00946] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00947] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00948] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01290] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00949] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01292] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01294] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01296] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01298] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0094f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00950] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00951] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00952] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00953] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00954] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00955] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00956] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00957] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00958] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00959] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0095f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00960] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00961] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00962] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00963] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00964] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00965] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00966] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00967] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00968] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00969] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0096f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00970] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00971] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00972] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00973] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00974] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00975] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00976] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00977] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00978] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00979] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0097f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00980] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01300] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00981] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01302] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00982] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01304] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00983] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01306] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00984] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01308] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00985] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00986] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00987] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00988] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01310] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00989] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01312] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01314] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01316] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01318] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0098f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00990] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01320] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00991] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01322] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00992] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01324] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00993] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01326] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00994] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01328] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00995] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00996] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00997] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00998] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01330] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00999] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01332] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01334] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01336] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01338] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h0099f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01340] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01342] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01344] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01346] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01348] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01350] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009a9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01352] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009aa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01354] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01356] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01358] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009af] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01360] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01362] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01364] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01366] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01368] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01370] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009b9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01372] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01374] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009bb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01376] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009bc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01378] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009bd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009be] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009bf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01380] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01382] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01384] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01386] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01388] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01390] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009c9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01392] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01394] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009cb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01396] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009cc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01398] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009cd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009cf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009d9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009da] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009db] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009dc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009dd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009de] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009df] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009e9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009eb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009f9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009fe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h009ff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a00] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01400] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a01] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01402] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a02] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01404] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a03] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01406] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a04] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01408] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a05] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a06] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a07] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a08] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01410] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a09] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01412] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01414] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01416] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01418] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a0f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a10] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01420] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a11] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01422] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a12] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01424] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a13] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01426] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a14] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01428] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a15] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a16] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a17] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a18] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01430] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a19] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01432] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01434] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01436] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01438] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a1f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a20] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01440] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a21] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01442] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a22] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01444] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a23] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01446] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a24] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01448] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a25] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a26] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a27] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a28] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01450] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a29] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01452] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01454] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01456] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01458] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a2f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a30] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01460] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a31] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01462] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a32] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01464] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a33] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01466] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a34] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01468] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a35] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a36] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a37] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a38] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01470] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a39] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01472] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01474] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01476] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01478] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a3f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a40] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01480] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a41] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01482] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a42] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01484] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a43] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01486] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a44] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01488] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a45] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a46] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a47] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a48] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01490] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a49] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01492] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01494] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01496] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01498] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a4f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a50] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a51] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a52] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a53] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a54] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a55] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a56] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a57] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a58] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a59] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a5f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a60] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a61] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a62] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a63] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a64] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a65] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a66] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a67] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a68] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a69] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a6f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a70] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a71] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a72] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a73] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a74] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a75] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a76] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a77] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a78] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a79] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a7f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a80] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01500] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a81] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01502] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a82] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01504] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a83] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01506] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a84] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01508] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a85] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a86] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a87] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a88] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01510] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a89] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01512] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01514] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01516] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01518] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a8f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a90] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01520] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a91] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01522] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a92] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01524] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a93] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01526] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a94] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01528] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a95] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a96] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a97] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a98] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01530] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a99] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01532] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01534] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01536] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01538] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00a9f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01540] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01542] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01544] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01546] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01548] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01550] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aa9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01552] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aaa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01554] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01556] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01558] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aaf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01560] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01562] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01564] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01566] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01568] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01570] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ab9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01572] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01574] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01576] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01578] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00abf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01580] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01582] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01584] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01586] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01588] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01590] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ac9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01592] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01594] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00acb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01596] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00acc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01598] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00acd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ace] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00acf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ad9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ada] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00adb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00adc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00add] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ade] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00adf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ae9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aeb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00af9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00afe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00aff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b00] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01600] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b01] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01602] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b02] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01604] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b03] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01606] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b04] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01608] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b05] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b06] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b07] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b08] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01610] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b09] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01612] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01614] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01616] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01618] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b0f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b10] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01620] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b11] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01622] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b12] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01624] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b13] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01626] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b14] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01628] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b15] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b16] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b17] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b18] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01630] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b19] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01632] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01634] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01636] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01638] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b1f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b20] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01640] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b21] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01642] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b22] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01644] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b23] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01646] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b24] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01648] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b25] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b26] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b27] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b28] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01650] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b29] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01652] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01654] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01656] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01658] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b2f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b30] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01660] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b31] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01662] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b32] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01664] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b33] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01666] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b34] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01668] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b35] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b36] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b37] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b38] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01670] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b39] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01672] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01674] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01676] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01678] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b3f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b40] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01680] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b41] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01682] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b42] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01684] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b43] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01686] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b44] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01688] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b45] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b46] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b47] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b48] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01690] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b49] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01692] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01694] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01696] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01698] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b4f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b50] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b51] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b52] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b53] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b54] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b55] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b56] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b57] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b58] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b59] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b5f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b60] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b61] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b62] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b63] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b64] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b65] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b66] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b67] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b68] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b69] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b6f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b70] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b71] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b72] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b73] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b74] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b75] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b76] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b77] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b78] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b79] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b7f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b80] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01700] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b81] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01702] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b82] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01704] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b83] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01706] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b84] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01708] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b85] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b86] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b87] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b88] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01710] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b89] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01712] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01714] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01716] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01718] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b8f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b90] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01720] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b91] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01722] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b92] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01724] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b93] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01726] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b94] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01728] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b95] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b96] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b97] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b98] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01730] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b99] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01732] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01734] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01736] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01738] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00b9f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01740] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01742] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01744] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01746] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01748] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01750] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ba9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01752] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00baa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01754] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01756] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01758] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00baf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01760] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01762] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01764] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01766] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01768] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01770] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bb9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01772] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01774] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01776] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01778] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bbf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01780] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01782] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01784] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01786] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01788] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01790] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bc9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01792] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01794] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bcb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01796] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bcc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01798] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bcd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bcf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bd9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bda] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bdb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bdc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bdd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bde] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bdf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00be9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00beb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bf9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bfe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00bff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c00] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01800] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c01] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01802] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c02] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01804] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c03] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01806] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c04] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01808] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c05] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c06] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c07] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c08] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01810] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c09] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01812] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01814] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01816] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01818] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c0f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c10] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01820] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c11] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01822] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c12] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01824] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c13] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01826] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c14] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01828] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c15] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c16] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c17] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c18] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01830] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c19] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01832] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01834] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01836] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01838] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c1f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c20] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01840] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c21] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01842] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c22] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01844] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c23] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01846] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c24] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01848] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c25] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c26] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c27] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c28] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01850] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c29] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01852] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01854] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01856] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01858] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c2f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c30] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01860] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c31] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01862] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c32] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01864] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c33] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01866] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c34] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01868] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c35] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c36] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c37] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c38] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01870] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c39] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01872] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01874] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01876] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01878] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c3f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c40] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01880] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c41] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01882] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c42] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01884] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c43] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01886] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c44] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01888] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c45] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c46] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c47] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c48] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01890] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c49] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01892] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01894] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01896] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01898] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c4f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c50] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c51] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c52] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c53] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c54] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c55] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c56] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c57] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c58] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c59] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c5f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c60] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c61] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c62] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c63] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c64] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c65] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c66] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c67] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c68] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c69] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c6f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c70] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c71] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c72] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c73] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c74] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c75] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c76] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c77] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c78] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c79] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c7f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c80] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01900] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c81] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01902] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c82] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01904] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c83] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01906] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c84] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01908] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c85] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c86] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c87] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c88] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01910] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c89] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01912] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01914] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01916] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01918] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c8f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c90] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01920] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c91] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01922] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c92] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01924] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c93] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01926] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c94] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01928] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c95] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c96] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c97] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c98] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01930] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c99] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01932] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01934] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01936] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01938] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00c9f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01940] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01942] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01944] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01946] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01948] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01950] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ca9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01952] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00caa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01954] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01956] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01958] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00caf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01960] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01962] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01964] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01966] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01968] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01970] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cb9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01972] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01974] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01976] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01978] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cbf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01980] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01982] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01984] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01986] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01988] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01990] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cc9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01992] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01994] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ccb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01996] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ccc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01998] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ccd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ccf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019aa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cd9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cda] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cdb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cdc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cdd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cde] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019bc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cdf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019be] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019cc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ce9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ceb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ced] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019da] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019dc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019de] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cf9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cfe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00cff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d00] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d01] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d02] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d03] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d04] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d05] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d06] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d07] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d08] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d09] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d0f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d10] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d11] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d12] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d13] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d14] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d15] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d16] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d17] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d18] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d19] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d1f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d20] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d21] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d22] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d23] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d24] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d25] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d26] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d27] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d28] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d29] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d2f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d30] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d31] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d32] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d33] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d34] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d35] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d36] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d37] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d38] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d39] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d3f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d40] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d41] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d42] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d43] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d44] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d45] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d46] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d47] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d48] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d49] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d4f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d50] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d51] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d52] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d53] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d54] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d55] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aaa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d56] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d57] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d58] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d59] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d5f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d60] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d61] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d62] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d63] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d64] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d65] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d66] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01acc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d67] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ace] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d68] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d69] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ada] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01adc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d6f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ade] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d70] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d71] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d72] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d73] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d74] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d75] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d76] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d77] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d78] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d79] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d7f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d80] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d81] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d82] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d83] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d84] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d85] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d86] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d87] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d88] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d89] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d8f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d90] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d91] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d92] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d93] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d94] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d95] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d96] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d97] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d98] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d99] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00d9f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00da9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00daa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00daf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00db9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dbf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dc9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dcb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dcc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dcd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dcf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01baa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dd9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dda] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ddb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ddc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ddd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dde] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ddf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bcc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00de9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00deb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ded] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bdc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00def] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00df9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dfe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00dff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e00] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e01] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e02] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e03] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e04] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e05] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e06] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e07] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e08] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e09] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e0f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e10] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e11] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e12] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e13] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e14] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e15] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e16] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e17] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e18] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e19] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e1f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e20] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e21] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e22] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e23] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e24] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e25] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e26] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e27] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e28] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e29] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e2f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e30] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e31] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e32] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e33] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e34] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e35] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e36] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e37] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e38] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e39] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e3f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e40] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e41] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e42] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e43] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e44] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e45] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e46] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e47] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e48] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e49] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e4f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e50] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e51] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e52] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e53] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e54] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e55] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01caa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e56] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e57] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e58] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e59] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e5f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e60] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e61] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e62] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e63] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e64] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e65] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e66] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ccc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e67] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e68] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e69] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cdc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e6f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e70] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e71] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e72] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e73] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e74] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e75] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e76] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e77] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e78] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e79] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e7f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e80] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e81] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e82] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e83] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e84] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e85] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e86] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e87] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e88] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e89] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e8f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e90] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e91] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e92] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e93] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e94] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e95] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e96] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e97] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e98] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e99] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00e9f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ea9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eaa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ead] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eaf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eb9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ebf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ec9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ecb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ecc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ecd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ece] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ecf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01daa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ed9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eda] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00edb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00edc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00edd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ede] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00edf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dcc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ee9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eeb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ddc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ef9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00efe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00eff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f00] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f01] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f02] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f03] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f04] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f05] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f06] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f07] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f08] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f09] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f0f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f10] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f11] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f12] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f13] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f14] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f15] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f16] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f17] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f18] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f19] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f1f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f20] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f21] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f22] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f23] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f24] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f25] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f26] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f27] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f28] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f29] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f2f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f30] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f31] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f32] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f33] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f34] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f35] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f36] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f37] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f38] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f39] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f3f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f40] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f41] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f42] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f43] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f44] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f45] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f46] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f47] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f48] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f49] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f4f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f50] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f51] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f52] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f53] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f54] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f55] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eaa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f56] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f57] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f58] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f59] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f5f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f60] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f61] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f62] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f63] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f64] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f65] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f66] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ecc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f67] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ece] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f68] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f69] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01edc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f6f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ede] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f70] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f71] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f72] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f73] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f74] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f75] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f76] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f77] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f78] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f79] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f7f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f80] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f00] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f81] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f02] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f82] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f04] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f83] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f06] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f84] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f08] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f85] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f86] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f87] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f88] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f10] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f89] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f12] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f14] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f16] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f18] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f8f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f90] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f20] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f91] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f22] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f92] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f24] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f93] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f26] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f94] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f28] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f95] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f96] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f97] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f98] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f30] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f99] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f32] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9a] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f34] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9b] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f36] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9c] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f38] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9d] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9e] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00f9f] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f40] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f42] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f44] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f46] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f48] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f50] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fa9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f52] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00faa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f54] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fab] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f56] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fac] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f58] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fad] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fae] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00faf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f60] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f62] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f64] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f66] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f68] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f70] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fb9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f72] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fba] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f74] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f76] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f78] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fbf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f80] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f82] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f84] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f86] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f88] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f90] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fc9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f92] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fca] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f94] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fcb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f96] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fcc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f98] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fcd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9a] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fce] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9c] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fcf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9e] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01faa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fac] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fae] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fd9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fda] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fdb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fdc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fdd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fba] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fde] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fdf] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbe] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fca] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fcc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fce] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fe9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fea] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00feb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fec] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fed] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fda] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fee] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fdc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fef] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fde] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff0] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff1] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff2] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff3] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff4] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff5] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fea] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff6] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fec] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff7] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fee] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff8] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff0] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ff9] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff2] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffa] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff4] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffb] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff6] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffc] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff8] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffd] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffa] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00ffe] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffc] ;
//end
//always_comb begin // 
               I067cf36cf447510cb166aa42d93fc80279a816ddb8415245a2824f43cc242a5e['h00fff] =  I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffe] ;
//end
