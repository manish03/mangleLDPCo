//`include "GF2_LDPC_fgallag_0x00008_assign_inc.sv"
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00000] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00000] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00001] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00001] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00002] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00003] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00002] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00004] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00005] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00003] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00006] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00007] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00004] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00008] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00009] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00005] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000a] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000b] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00006] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000c] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000d] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00007] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000e] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000f] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00008] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00010] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00011] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00009] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00012] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00013] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000a] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00014] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00015] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000b] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00016] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00017] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000c] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00018] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00019] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000d] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001a] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001b] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000e] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001c] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001d] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0000f] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001e] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001f] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00010] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00020] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00021] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00011] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00022] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00023] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00012] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00024] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00025] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00013] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00026] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00027] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00014] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00028] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00029] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00015] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002a] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002b] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00016] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002c] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002d] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00017] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002e] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002f] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00018] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00030] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00031] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00019] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00032] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00033] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001a] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00034] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00035] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001b] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00036] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00037] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001c] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00038] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00039] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001d] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003a] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003b] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003c] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0001f] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003e] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003f] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00020] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00040] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00021] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00042] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00022] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00044] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00023] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00046] ;
//end
//always_comb begin
              I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00024] = 
          (!fgallag_sel['h00008]) ? 
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00048] : //%
                       I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00049] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00025] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00026] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00027] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00028] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00050] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00029] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00052] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00054] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00056] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00058] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0002f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00030] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00060] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00031] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00062] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00032] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00064] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00033] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00066] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00034] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00068] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00035] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00036] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00037] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00038] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00070] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00039] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00072] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00074] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00076] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00078] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0003f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00040] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00080] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00041] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00082] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00042] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00084] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00043] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00086] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00044] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00088] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00045] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00046] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00047] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00048] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00090] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00049] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00092] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00094] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00096] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00098] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0004f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00050] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00051] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00052] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00053] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00054] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00055] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00056] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00057] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00058] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00059] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0005f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00060] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00061] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00062] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00063] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00064] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00065] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00066] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00067] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00068] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00069] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0006f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00070] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00071] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00072] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00073] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00074] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00075] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00076] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00077] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00078] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00079] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0007f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00080] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00100] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00081] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00102] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00082] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00104] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00083] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00106] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00084] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00108] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00085] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00086] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00087] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00088] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00110] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00089] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00112] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00114] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00116] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00118] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0008f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00090] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00120] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00091] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00122] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00092] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00124] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00093] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00126] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00094] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00128] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00095] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00096] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00097] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00098] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00130] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00099] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00132] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00134] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00136] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00138] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0009f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00140] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00142] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00144] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00146] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00148] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00150] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000a9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00152] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000aa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00154] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ab] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00156] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ac] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00158] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ad] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ae] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000af] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00160] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00162] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00164] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00166] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00168] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00170] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000b9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00172] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ba] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00174] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000bb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00176] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000bc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00178] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000bd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000be] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000bf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00180] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00182] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00184] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00186] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00188] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00190] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000c9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00192] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ca] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00194] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000cb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00196] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000cc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00198] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000cd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ce] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000cf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000d9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000da] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000db] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000dc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000dd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000de] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000df] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000e9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ea] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000eb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ec] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ed] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ee] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ef] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000f9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000fe] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h000ff] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00100] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00200] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00101] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00202] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00102] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00204] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00103] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00206] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00104] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00208] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00105] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00106] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00107] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00108] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00210] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00109] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00212] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00214] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00216] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00218] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0010f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00110] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00220] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00111] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00222] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00112] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00224] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00113] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00226] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00114] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00228] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00115] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00116] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00117] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00118] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00230] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00119] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00232] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00234] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00236] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00238] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0011f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00120] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00240] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00121] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00242] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00122] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00244] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00123] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00246] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00124] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00248] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00125] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00126] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00127] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00128] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00250] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00129] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00252] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00254] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00256] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00258] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0012f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00130] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00260] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00131] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00262] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00132] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00264] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00133] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00266] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00134] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00268] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00135] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00136] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00137] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00138] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00270] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00139] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00272] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00274] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00276] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00278] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0013f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00140] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00280] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00141] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00282] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00142] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00284] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00143] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00286] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00144] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00288] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00145] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00146] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00147] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00148] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00290] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00149] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00292] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00294] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00296] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00298] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0014f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00150] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00151] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00152] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00153] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00154] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00155] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00156] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00157] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00158] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00159] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0015f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00160] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00161] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00162] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00163] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00164] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00165] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00166] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00167] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00168] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00169] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0016f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00170] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00171] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00172] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00173] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00174] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00175] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00176] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00177] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00178] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00179] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0017f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00180] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00300] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00181] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00302] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00182] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00304] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00183] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00306] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00184] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00308] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00185] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00186] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00187] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00188] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00310] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00189] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00312] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00314] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00316] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00318] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0018f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00190] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00320] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00191] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00322] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00192] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00324] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00193] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00326] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00194] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00328] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00195] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00196] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00197] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00198] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00330] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00199] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00332] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00334] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00336] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00338] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0019f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00340] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00342] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00344] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00346] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00348] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00350] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001a9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00352] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001aa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00354] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ab] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00356] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ac] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00358] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ad] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ae] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001af] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00360] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00362] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00364] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00366] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00368] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00370] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001b9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00372] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ba] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00374] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001bb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00376] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001bc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00378] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001bd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001be] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001bf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00380] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00382] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00384] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00386] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00388] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00390] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001c9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00392] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ca] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00394] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001cb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00396] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001cc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00398] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001cd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ce] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001cf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001d9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001da] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001db] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001dc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001dd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001de] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001df] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001e9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ea] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001eb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ec] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ed] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ee] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ef] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001f9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001fe] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h001ff] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00200] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00400] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00201] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00402] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00202] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00404] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00203] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00406] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00204] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00408] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00205] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00206] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00207] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00208] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00410] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00209] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00412] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00414] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00416] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00418] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0020f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00210] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00420] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00211] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00422] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00212] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00424] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00213] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00426] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00214] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00428] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00215] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00216] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00217] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00218] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00430] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00219] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00432] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00434] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00436] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00438] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0021f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00220] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00440] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00221] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00442] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00222] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00444] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00223] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00446] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00224] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00448] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00225] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00226] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00227] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00228] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00450] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00229] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00452] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00454] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00456] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00458] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0022f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00230] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00460] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00231] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00462] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00232] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00464] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00233] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00466] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00234] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00468] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00235] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00236] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00237] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00238] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00470] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00239] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00472] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00474] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00476] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00478] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0023f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00240] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00480] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00241] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00482] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00242] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00484] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00243] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00486] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00244] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00488] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00245] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00246] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00247] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00248] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00490] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00249] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00492] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00494] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00496] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00498] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0024f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00250] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00251] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00252] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00253] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00254] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00255] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00256] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00257] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00258] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00259] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0025f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00260] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00261] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00262] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00263] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00264] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00265] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00266] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00267] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00268] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00269] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0026f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00270] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00271] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00272] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00273] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00274] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00275] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00276] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00277] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00278] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00279] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0027f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00280] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00500] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00281] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00502] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00282] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00504] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00283] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00506] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00284] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00508] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00285] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00286] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00287] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00288] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00510] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00289] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00512] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00514] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00516] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00518] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0028f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00290] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00520] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00291] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00522] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00292] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00524] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00293] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00526] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00294] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00528] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00295] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00296] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00297] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00298] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00530] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00299] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00532] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00534] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00536] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00538] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0029f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00540] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00542] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00544] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00546] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00548] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00550] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002a9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00552] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002aa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00554] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ab] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00556] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ac] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00558] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ad] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ae] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002af] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00560] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00562] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00564] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00566] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00568] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00570] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002b9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00572] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ba] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00574] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002bb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00576] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002bc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00578] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002bd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002be] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002bf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00580] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00582] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00584] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00586] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00588] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00590] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002c9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00592] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ca] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00594] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002cb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00596] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002cc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00598] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002cd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ce] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002cf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002d9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002da] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002db] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002dc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002dd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002de] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002df] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002e9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ea] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002eb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ec] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ed] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ee] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ef] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002f9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002fe] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h002ff] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00300] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00600] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00301] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00602] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00302] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00604] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00303] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00606] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00304] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00608] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00305] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00306] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00307] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00308] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00610] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00309] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00612] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00614] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00616] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00618] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0030f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00310] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00620] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00311] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00622] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00312] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00624] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00313] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00626] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00314] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00628] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00315] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00316] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00317] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00318] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00630] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00319] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00632] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00634] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00636] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00638] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0031f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00320] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00640] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00321] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00642] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00322] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00644] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00323] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00646] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00324] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00648] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00325] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00326] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00327] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00328] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00650] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00329] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00652] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00654] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00656] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00658] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0032f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00330] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00660] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00331] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00662] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00332] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00664] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00333] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00666] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00334] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00668] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00335] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00336] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00337] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00338] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00670] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00339] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00672] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00674] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00676] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00678] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0033f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00340] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00680] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00341] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00682] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00342] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00684] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00343] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00686] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00344] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00688] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00345] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00346] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00347] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00348] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00690] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00349] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00692] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00694] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00696] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00698] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0034f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00350] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00351] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00352] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00353] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00354] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00355] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00356] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00357] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00358] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00359] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0035f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00360] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00361] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00362] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00363] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00364] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00365] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00366] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00367] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00368] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00369] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0036f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00370] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00371] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00372] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00373] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00374] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00375] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00376] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00377] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00378] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00379] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0037f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fe] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00380] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00700] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00381] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00702] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00382] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00704] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00383] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00706] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00384] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00708] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00385] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00386] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00387] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00388] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00710] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00389] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00712] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00714] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00716] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00718] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0038f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00390] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00720] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00391] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00722] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00392] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00724] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00393] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00726] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00394] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00728] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00395] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00396] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00397] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00398] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00730] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h00399] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00732] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039a] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00734] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039b] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00736] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039c] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00738] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039d] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039e] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h0039f] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00740] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00742] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00744] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00746] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00748] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00750] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003a9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00752] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003aa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00754] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ab] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00756] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ac] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00758] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ad] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ae] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003af] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00760] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00762] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00764] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00766] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00768] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00770] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003b9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00772] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ba] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00774] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003bb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00776] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003bc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00778] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003bd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003be] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003bf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00780] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00782] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00784] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00786] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00788] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00790] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003c9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00792] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ca] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00794] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003cb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00796] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003cc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00798] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003cd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079a] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ce] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079c] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003cf] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079e] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007aa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ac] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ae] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003d9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003da] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003db] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003dc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003dd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ba] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003de] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007bc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003df] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007be] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ca] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007cc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ce] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003e9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ea] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003eb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ec] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ed] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007da] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ee] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007dc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ef] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007de] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f0] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f1] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f2] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f3] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f4] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f5] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ea] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f6] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ec] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f7] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ee] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f8] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f0] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003f9] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f2] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fa] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f4] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fb] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f6] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fc] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f8] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fd] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fa] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003fe] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fc] ;
//end
//always_comb begin // 
               I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322['h003ff] =  I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fe] ;
//end
