 reg  ['h1f:0] [$clog2('h7000+1)-1:0] I1f3af771a6bf6da6d9e448fb87a2d186 ;
