 reg  ['h1:0] [$clog2('h7000+1)-1:0] Ic7e91188980d728ad34dbe693d9a6e04 ;
