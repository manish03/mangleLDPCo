//`include "GF2_LDPC_flogtanh_0x00007_assign_inc.sv"
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00000] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00000] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00001] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00001] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00002] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00003] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00002] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00004] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00005] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00003] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00006] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00007] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00004] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00008] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00009] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00005] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000a] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000b] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00006] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000d] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00007] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000f] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00008] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00010] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00011] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00009] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00012] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00013] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0000a] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00014] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00015] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0000b] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00016] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00017] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0000c] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00018] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00019] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0000d] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001a] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001b] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0000e] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001d] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0000f] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001f] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00010] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00020] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00021] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00011] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00022] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00023] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00012] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00024] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00025] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00013] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00026] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00027] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00014] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00028] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00029] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00015] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002a] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002b] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00016] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002d] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00017] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002f] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00018] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00030] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00031] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00019] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00032] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00033] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0001a] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00034] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00035] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0001b] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00036] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00037] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0001c] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00038] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00039] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0001d] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003a] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003b] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0001e] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003d] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0001f] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003f] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00020] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00040] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00041] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00021] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00042] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00043] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00022] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00044] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00045] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00023] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00046] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00047] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00024] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00048] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00049] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00025] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004a] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004b] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00026] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004d] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00027] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004f] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00028] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00050] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00051] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00029] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00052] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00053] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0002a] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00054] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00055] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0002b] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00056] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00057] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0002c] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00058] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00059] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0002d] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005a] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005b] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0002e] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005d] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0002f] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005f] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00030] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00060] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00061] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00031] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00062] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00063] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00032] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00064] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00065] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00033] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00066] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00067] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00034] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00068] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00069] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00035] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006a] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00036] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006c] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006d] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00037] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006e] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00038] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00070] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00071] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00039] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00072] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0003a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00074] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0003b] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00076] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00077] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0003c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00078] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0003d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0003e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007c] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h0003f] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007e] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007f] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00040] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00080] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00041] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00082] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00042] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00084] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00043] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00086] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00044] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00088] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00045] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00046] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00047] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008e] ;
//end
//always_comb begin
              I38e438ab568822a1c40149a2acc5d876['h00048] = 
          (!flogtanh_sel['h00007]) ? 
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00090] : //%
                       I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00091] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00049] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00092] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0004a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00094] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0004b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00096] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0004c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00098] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0004d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0004e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0004f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00050] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00051] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00052] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00053] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00054] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00055] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00056] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00057] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00058] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00059] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0005a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0005b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0005c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0005d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0005e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0005f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00060] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00061] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00062] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00063] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00064] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00065] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00066] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00067] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00068] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00069] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0006a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0006b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0006c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0006d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0006e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0006f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00070] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00071] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00072] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00073] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00074] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00075] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00076] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00077] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00078] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00079] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0007a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0007b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0007c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0007d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0007e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0007f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00080] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00100] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00081] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00102] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00082] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00104] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00083] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00106] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00084] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00108] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00085] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00086] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00087] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00088] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00110] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00089] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00112] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0008a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00114] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0008b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00116] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0008c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00118] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0008d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0008e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0008f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00090] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00120] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00091] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00122] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00092] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00124] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00093] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00126] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00094] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00128] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00095] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00096] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00097] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00098] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00130] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00099] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00132] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0009a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00134] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0009b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00136] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0009c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00138] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0009d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0009e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0009f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00140] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00142] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00144] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00146] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00148] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00150] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00152] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00154] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00156] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00158] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00160] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00162] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00164] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00166] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00168] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00170] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00172] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00174] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00176] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00178] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00180] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00182] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00184] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00186] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00188] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00190] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00192] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00194] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00196] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00198] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h000ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00100] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00200] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00101] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00202] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00102] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00204] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00103] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00206] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00104] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00208] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00105] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00106] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00107] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00108] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00210] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00109] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00212] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0010a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00214] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0010b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00216] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0010c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00218] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0010d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0010e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0010f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00110] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00220] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00111] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00222] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00112] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00224] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00113] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00226] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00114] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00228] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00115] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00116] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00117] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00118] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00230] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00119] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00232] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0011a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00234] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0011b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00236] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0011c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00238] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0011d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0011e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0011f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00120] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00240] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00121] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00242] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00122] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00244] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00123] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00246] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00124] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00248] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00125] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00126] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00127] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00128] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00250] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00129] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00252] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0012a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00254] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0012b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00256] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0012c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00258] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0012d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0012e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0012f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00130] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00260] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00131] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00262] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00132] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00264] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00133] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00266] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00134] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00268] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00135] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00136] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00137] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00138] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00270] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00139] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00272] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0013a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00274] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0013b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00276] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0013c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00278] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0013d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0013e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0013f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00140] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00280] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00141] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00282] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00142] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00284] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00143] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00286] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00144] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00288] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00145] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00146] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00147] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00148] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00290] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00149] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00292] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0014a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00294] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0014b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00296] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0014c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00298] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0014d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0014e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0014f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00150] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00151] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00152] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00153] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00154] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00155] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00156] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00157] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00158] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00159] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0015a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0015b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0015c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0015d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0015e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0015f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00160] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00161] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00162] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00163] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00164] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00165] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00166] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00167] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00168] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00169] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0016a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0016b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0016c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0016d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0016e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0016f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00170] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00171] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00172] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00173] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00174] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00175] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00176] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00177] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00178] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00179] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0017a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0017b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0017c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0017d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0017e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0017f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00180] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00300] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00181] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00302] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00182] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00304] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00183] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00306] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00184] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00308] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00185] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00186] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00187] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00188] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00310] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00189] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00312] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0018a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00314] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0018b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00316] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0018c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00318] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0018d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0018e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0018f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00190] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00320] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00191] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00322] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00192] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00324] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00193] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00326] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00194] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00328] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00195] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00196] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00197] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00198] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00330] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00199] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00332] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0019a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00334] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0019b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00336] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0019c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00338] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0019d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0019e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0019f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00340] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00342] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00344] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00346] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00348] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00350] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00352] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00354] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00356] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00358] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00360] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00362] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00364] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00366] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00368] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00370] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00372] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00374] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00376] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00378] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00380] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00382] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00384] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00386] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00388] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00390] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00392] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00394] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00396] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00398] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h001ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00200] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00400] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00201] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00402] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00202] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00404] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00203] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00406] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00204] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00408] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00205] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00206] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00207] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00208] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00410] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00209] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00412] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0020a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00414] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0020b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00416] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0020c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00418] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0020d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0020e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0020f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00210] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00420] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00211] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00422] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00212] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00424] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00213] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00426] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00214] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00428] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00215] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00216] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00217] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00218] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00430] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00219] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00432] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0021a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00434] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0021b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00436] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0021c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00438] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0021d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0021e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0021f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00220] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00440] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00221] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00442] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00222] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00444] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00223] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00446] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00224] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00448] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00225] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00226] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00227] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00228] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00450] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00229] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00452] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0022a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00454] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0022b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00456] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0022c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00458] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0022d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0022e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0022f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00230] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00460] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00231] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00462] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00232] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00464] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00233] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00466] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00234] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00468] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00235] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00236] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00237] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00238] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00470] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00239] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00472] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0023a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00474] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0023b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00476] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0023c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00478] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0023d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0023e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0023f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00240] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00480] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00241] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00482] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00242] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00484] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00243] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00486] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00244] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00488] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00245] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00246] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00247] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00248] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00490] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00249] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00492] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0024a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00494] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0024b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00496] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0024c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00498] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0024d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0024e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0024f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00250] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00251] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00252] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00253] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00254] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00255] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00256] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00257] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00258] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00259] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0025a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0025b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0025c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0025d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0025e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0025f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00260] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00261] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00262] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00263] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00264] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00265] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00266] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00267] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00268] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00269] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0026a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0026b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0026c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0026d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0026e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0026f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00270] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00271] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00272] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00273] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00274] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00275] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00276] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00277] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00278] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00279] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0027a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0027b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0027c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0027d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0027e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0027f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00280] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00500] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00281] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00502] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00282] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00504] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00283] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00506] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00284] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00508] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00285] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00286] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00287] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00288] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00510] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00289] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00512] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0028a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00514] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0028b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00516] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0028c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00518] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0028d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0028e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0028f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00290] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00520] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00291] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00522] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00292] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00524] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00293] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00526] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00294] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00528] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00295] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00296] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00297] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00298] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00530] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00299] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00532] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0029a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00534] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0029b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00536] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0029c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00538] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0029d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0029e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0029f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00540] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00542] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00544] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00546] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00548] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00550] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00552] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00554] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00556] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00558] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00560] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00562] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00564] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00566] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00568] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00570] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00572] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00574] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00576] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00578] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00580] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00582] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00584] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00586] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00588] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00590] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00592] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00594] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00596] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00598] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h002ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00300] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00600] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00301] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00602] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00302] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00604] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00303] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00606] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00304] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00608] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00305] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00306] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00307] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00308] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00610] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00309] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00612] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0030a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00614] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0030b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00616] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0030c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00618] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0030d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0030e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0030f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00310] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00620] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00311] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00622] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00312] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00624] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00313] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00626] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00314] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00628] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00315] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00316] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00317] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00318] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00630] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00319] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00632] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0031a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00634] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0031b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00636] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0031c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00638] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0031d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0031e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0031f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00320] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00640] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00321] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00642] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00322] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00644] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00323] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00646] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00324] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00648] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00325] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00326] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00327] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00328] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00650] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00329] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00652] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0032a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00654] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0032b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00656] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0032c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00658] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0032d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0032e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0032f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00330] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00660] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00331] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00662] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00332] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00664] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00333] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00666] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00334] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00668] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00335] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00336] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00337] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00338] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00670] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00339] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00672] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0033a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00674] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0033b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00676] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0033c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00678] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0033d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0033e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0033f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00340] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00680] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00341] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00682] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00342] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00684] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00343] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00686] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00344] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00688] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00345] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00346] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00347] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00348] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00690] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00349] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00692] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0034a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00694] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0034b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00696] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0034c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00698] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0034d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0034e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0034f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00350] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00351] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00352] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00353] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00354] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00355] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00356] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00357] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00358] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00359] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0035a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0035b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0035c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0035d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0035e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0035f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00360] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00361] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00362] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00363] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00364] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00365] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00366] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00367] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00368] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00369] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0036a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0036b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0036c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0036d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0036e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0036f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00370] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00371] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00372] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00373] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00374] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00375] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00376] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00377] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00378] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00379] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0037a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0037b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0037c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0037d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0037e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0037f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00380] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00700] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00381] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00702] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00382] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00704] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00383] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00706] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00384] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00708] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00385] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00386] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00387] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00388] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00710] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00389] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00712] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0038a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00714] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0038b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00716] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0038c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00718] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0038d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0038e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0038f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00390] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00720] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00391] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00722] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00392] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00724] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00393] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00726] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00394] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00728] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00395] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00396] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00397] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00398] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00730] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00399] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00732] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0039a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00734] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0039b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00736] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0039c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00738] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0039d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0039e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0039f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00740] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00742] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00744] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00746] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00748] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00750] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00752] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00754] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00756] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00758] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00760] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00762] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00764] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00766] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00768] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00770] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00772] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00774] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00776] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00778] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00780] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00782] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00784] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00786] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00788] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00790] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00792] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00794] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00796] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00798] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h003ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00400] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00800] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00401] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00802] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00402] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00804] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00403] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00806] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00404] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00808] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00405] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00406] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00407] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00408] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00810] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00409] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00812] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0040a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00814] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0040b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00816] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0040c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00818] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0040d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0040e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0040f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00410] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00820] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00411] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00822] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00412] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00824] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00413] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00826] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00414] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00828] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00415] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00416] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00417] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00418] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00830] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00419] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00832] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0041a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00834] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0041b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00836] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0041c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00838] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0041d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0041e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0041f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00420] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00840] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00421] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00842] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00422] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00844] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00423] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00846] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00424] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00848] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00425] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00426] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00427] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00428] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00850] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00429] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00852] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0042a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00854] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0042b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00856] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0042c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00858] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0042d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0042e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0042f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00430] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00860] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00431] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00862] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00432] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00864] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00433] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00866] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00434] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00868] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00435] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00436] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00437] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00438] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00870] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00439] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00872] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0043a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00874] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0043b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00876] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0043c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00878] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0043d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0043e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0043f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00440] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00880] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00441] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00882] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00442] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00884] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00443] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00886] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00444] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00888] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00445] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00446] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00447] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00448] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00890] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00449] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00892] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0044a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00894] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0044b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00896] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0044c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00898] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0044d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0044e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0044f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00450] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00451] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00452] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00453] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00454] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00455] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00456] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00457] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00458] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00459] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0045a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0045b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0045c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0045d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0045e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0045f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00460] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00461] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00462] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00463] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00464] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00465] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00466] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00467] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00468] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00469] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0046a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0046b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0046c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0046d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0046e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0046f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00470] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00471] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00472] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00473] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00474] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00475] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00476] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00477] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00478] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00479] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0047a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0047b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0047c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0047d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0047e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0047f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00480] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00900] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00481] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00902] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00482] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00904] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00483] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00906] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00484] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00908] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00485] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00486] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00487] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00488] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00910] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00489] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00912] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0048a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00914] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0048b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00916] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0048c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00918] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0048d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0048e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0048f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00490] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00920] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00491] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00922] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00492] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00924] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00493] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00926] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00494] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00928] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00495] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00496] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00497] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00498] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00930] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00499] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00932] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0049a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00934] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0049b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00936] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0049c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00938] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0049d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0049e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0049f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00940] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00942] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00944] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00946] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00948] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00950] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00952] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00954] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00956] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00958] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00960] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00962] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00964] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00966] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00968] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00970] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00972] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00974] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00976] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00978] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00980] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00982] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00984] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00986] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00988] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00990] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00992] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00994] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00996] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00998] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009aa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009bc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009be] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009cc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009da] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009dc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009de] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h004ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00500] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a00] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00501] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a02] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00502] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a04] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00503] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a06] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00504] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a08] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00505] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00506] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00507] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00508] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a10] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00509] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a12] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0050a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a14] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0050b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a16] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0050c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a18] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0050d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0050e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0050f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00510] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a20] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00511] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a22] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00512] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a24] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00513] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a26] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00514] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a28] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00515] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00516] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00517] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00518] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a30] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00519] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a32] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0051a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a34] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0051b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a36] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0051c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a38] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0051d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0051e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0051f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00520] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a40] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00521] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a42] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00522] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a44] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00523] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a46] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00524] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a48] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00525] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00526] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00527] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00528] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a50] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00529] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a52] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0052a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a54] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0052b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a56] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0052c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a58] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0052d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0052e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0052f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00530] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a60] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00531] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a62] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00532] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a64] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00533] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a66] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00534] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a68] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00535] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00536] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00537] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00538] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a70] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00539] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a72] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0053a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a74] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0053b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a76] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0053c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a78] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0053d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0053e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0053f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00540] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a80] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00541] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a82] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00542] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a84] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00543] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a86] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00544] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a88] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00545] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00546] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00547] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00548] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a90] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00549] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a92] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0054a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a94] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0054b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a96] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0054c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a98] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0054d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0054e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0054f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00550] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00551] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00552] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00553] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00554] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00555] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aaa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00556] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00557] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00558] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00559] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0055a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0055b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0055c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0055d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0055e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0055f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00560] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00561] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00562] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00563] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00564] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00565] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00566] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00acc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00567] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ace] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00568] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00569] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0056a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0056b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0056c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0056d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ada] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0056e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00adc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0056f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ade] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00570] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00571] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00572] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00573] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00574] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00575] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00576] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00577] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00578] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00579] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0057a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0057b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0057c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0057d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0057e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0057f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00580] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b00] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00581] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b02] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00582] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b04] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00583] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b06] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00584] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b08] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00585] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00586] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00587] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00588] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b10] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00589] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b12] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0058a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b14] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0058b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b16] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0058c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b18] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0058d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0058e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0058f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00590] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b20] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00591] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b22] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00592] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b24] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00593] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b26] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00594] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b28] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00595] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00596] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00597] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00598] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b30] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00599] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b32] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0059a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b34] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0059b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b36] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0059c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b38] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0059d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0059e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0059f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b40] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b42] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b44] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b46] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b48] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b50] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b52] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b54] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b56] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b58] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b60] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b62] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b64] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b66] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b68] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b70] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b72] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b74] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b76] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b78] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b80] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b82] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b84] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b86] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b88] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b90] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b92] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b94] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b96] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b98] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00baa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bcc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bda] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bdc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bde] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h005ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00600] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c00] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00601] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c02] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00602] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c04] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00603] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c06] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00604] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c08] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00605] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00606] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00607] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00608] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c10] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00609] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c12] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0060a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c14] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0060b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c16] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0060c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c18] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0060d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0060e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0060f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00610] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c20] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00611] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c22] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00612] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c24] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00613] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c26] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00614] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c28] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00615] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00616] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00617] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00618] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c30] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00619] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c32] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0061a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c34] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0061b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c36] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0061c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c38] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0061d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0061e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0061f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00620] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c40] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00621] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c42] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00622] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c44] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00623] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c46] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00624] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c48] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00625] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00626] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00627] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00628] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c50] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00629] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c52] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0062a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c54] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0062b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c56] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0062c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c58] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0062d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0062e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0062f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00630] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c60] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00631] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c62] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00632] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c64] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00633] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c66] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00634] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c68] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00635] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00636] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00637] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00638] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c70] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00639] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c72] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0063a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c74] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0063b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c76] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0063c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c78] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0063d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0063e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0063f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00640] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c80] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00641] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c82] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00642] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c84] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00643] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c86] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00644] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c88] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00645] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00646] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00647] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00648] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c90] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00649] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c92] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0064a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c94] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0064b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c96] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0064c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c98] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0064d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0064e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0064f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00650] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00651] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00652] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00653] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00654] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00655] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00caa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00656] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00657] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00658] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00659] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0065a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0065b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0065c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0065d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0065e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0065f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00660] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00661] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00662] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00663] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00664] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00665] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00666] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ccc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00667] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00668] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00669] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0066a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0066b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0066c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0066d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cda] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0066e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cdc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0066f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cde] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00670] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00671] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00672] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00673] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00674] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00675] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00676] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00677] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00678] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00679] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0067a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0067b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0067c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0067d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0067e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0067f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00680] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d00] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00681] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d02] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00682] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d04] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00683] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d06] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00684] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d08] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00685] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00686] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00687] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00688] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d10] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00689] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d12] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0068a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d14] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0068b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d16] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0068c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d18] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0068d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0068e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0068f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00690] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d20] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00691] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d22] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00692] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d24] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00693] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d26] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00694] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d28] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00695] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00696] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00697] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00698] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d30] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00699] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d32] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0069a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d34] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0069b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d36] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0069c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d38] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0069d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0069e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0069f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d40] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d42] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d44] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d46] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d48] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d50] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d52] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d54] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d56] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d58] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d60] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d62] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d64] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d66] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d68] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d70] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d72] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d74] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d76] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d78] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d80] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d82] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d84] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d86] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d88] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d90] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d92] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d94] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d96] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d98] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00daa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dcc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dda] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ddc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dde] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h006ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00700] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e00] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00701] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e02] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00702] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e04] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00703] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e06] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00704] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e08] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00705] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00706] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00707] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00708] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e10] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00709] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e12] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0070a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e14] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0070b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e16] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0070c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e18] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0070d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0070e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0070f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00710] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e20] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00711] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e22] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00712] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e24] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00713] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e26] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00714] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e28] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00715] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00716] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00717] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00718] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e30] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00719] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e32] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0071a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e34] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0071b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e36] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0071c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e38] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0071d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0071e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0071f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00720] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e40] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00721] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e42] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00722] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e44] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00723] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e46] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00724] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e48] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00725] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00726] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00727] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00728] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e50] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00729] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e52] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0072a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e54] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0072b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e56] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0072c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e58] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0072d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0072e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0072f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00730] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e60] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00731] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e62] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00732] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e64] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00733] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e66] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00734] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e68] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00735] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00736] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00737] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00738] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e70] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00739] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e72] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0073a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e74] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0073b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e76] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0073c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e78] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0073d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0073e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0073f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00740] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e80] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00741] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e82] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00742] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e84] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00743] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e86] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00744] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e88] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00745] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00746] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00747] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00748] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e90] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00749] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e92] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0074a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e94] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0074b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e96] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0074c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e98] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0074d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0074e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0074f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00750] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00751] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00752] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00753] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00754] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00755] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eaa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00756] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00757] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00758] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00759] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0075a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0075b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0075c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0075d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0075e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0075f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00760] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00761] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00762] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00763] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00764] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00765] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00766] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ecc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00767] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ece] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00768] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00769] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0076a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0076b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0076c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0076d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eda] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0076e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00edc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0076f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ede] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00770] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00771] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00772] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00773] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00774] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00775] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00776] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00777] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00778] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00779] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0077a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0077b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0077c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0077d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0077e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0077f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00780] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f00] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00781] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f02] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00782] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f04] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00783] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f06] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00784] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f08] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00785] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00786] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00787] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00788] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f10] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00789] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f12] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0078a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f14] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0078b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f16] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0078c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f18] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0078d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0078e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0078f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00790] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f20] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00791] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f22] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00792] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f24] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00793] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f26] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00794] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f28] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00795] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00796] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00797] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00798] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f30] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h00799] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f32] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0079a] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f34] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0079b] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f36] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0079c] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f38] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0079d] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0079e] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h0079f] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f40] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f42] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f44] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f46] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f48] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f50] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007a9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f52] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007aa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f54] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ab] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f56] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ac] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f58] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ad] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ae] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007af] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f60] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f62] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f64] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f66] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f68] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f70] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007b9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f72] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ba] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f74] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007bb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f76] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007bc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f78] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007bd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007be] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007bf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f80] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f82] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f84] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f86] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f88] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f90] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007c9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f92] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ca] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f94] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007cb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f96] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007cc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f98] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007cd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9a] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ce] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9c] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007cf] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9e] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00faa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fac] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fae] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007d9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007da] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007db] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007dc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007dd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fba] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007de] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007df] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbe] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fca] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fcc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fce] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007e9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ea] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007eb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ec] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ed] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fda] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ee] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fdc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ef] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fde] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f0] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f1] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f2] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f3] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f4] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f5] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fea] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f6] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fec] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f7] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fee] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f8] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff0] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007f9] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff2] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007fa] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff4] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007fb] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff6] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007fc] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff8] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007fd] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffa] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007fe] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffc] ;
//end
//always_comb begin // 
               I38e438ab568822a1c40149a2acc5d876['h007ff] =  I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffe] ;
//end
