 reg  ['h3fff:0] [$clog2('h7000+1)-1:0] I0310077d53ae4ed9904df42e3f81c634 ;
