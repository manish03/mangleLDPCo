//`include "GF2_LDPC_fgallag_0x00011_assign_inc.sv"
//always_comb begin
              I34f69b29975fc71eeee92e6ac4210723['h00000] = 
          (!fgallag_sel['h00011]) ? 
                       I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00000] : //%
                       I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00001] ;
//end
//always_comb begin // 
               I34f69b29975fc71eeee92e6ac4210723['h00001] =  I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00002] ;
//end
