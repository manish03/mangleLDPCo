 reg  ['h1:0] [$clog2('h7000+1)-1:0] I1e92c8d19105281ae50f051d46adab55b63f3805ee886a8045e61a0f72842ab4 ;
