              Ib215a1b985e00121a1c48cf2ddae939a = 
          (!fgallag_sel[2]) ? 
                       I72dd1fc26b57d741390612b9bcffab1d: 
                       I98c43e93e5f943a7b07ef09985f97014;
              I0d9537bea5895773b487fb385690c92c = 
          (!fgallag_sel[2]) ? 
                       I434c16361fa147e26f4d2c4cc6d69150: 
                       I9e87743bade1ee6fbfdd119cbdb0a3cb;
              I287708a4c364df837b06049357518409 = 
          (!fgallag_sel[2]) ? 
                       I1e6255cf954cd5a58c52ff8e6a55bdbc: 
                       I77a73f3832687dababc30666ac62d1af;
              I9e69bf6d258b709d9706052822d9ae16 = 
          (!fgallag_sel[2]) ? 
                       Iacdfa68e9ab161a0e6c7e559b9954640: 
                       Iedc0dfa42eaada48be02e65be4b39615;
              I0d187ebb6dbedda971b33ceebb6f17eb = 
          (!fgallag_sel[2]) ? 
                       Ib4fb78755c536a284004e41f584d99fb: 
                       I5156cd5e3f0fe53ad559b342c818f41a;
              I83ab1426707044dca3ed926493081311 = 
          (!fgallag_sel[2]) ? 
                       I3cf816bf7fd922df289b13766e931e17: 
                       Ibf2a30f91bd9050391913c02be7c8cad;
              Ib402ea81f3ba6d26feac26905f0c5edc = 
          (!fgallag_sel[2]) ? 
                       Iea12e263d5883f93023d784884645969: 
                       I550762460d0217d3c91c5112546b7929;
              I457501e8372fe81287f139beeaad0452 = 
          (!fgallag_sel[2]) ? 
                       I0d8eaf22a03a0102d8bf7a53a7737943: 
                       I8017a4f092179605074076e8b5690842;
              I6f3ecf6c401215c1242c6d31cb4158d7 = 
          (!fgallag_sel[2]) ? 
                       I57160990c295512e2d98c301632c5120: 
                       Id9f3f35bc6917416d6826d471f8ea441;
              Ia439d59ddaa34c9a8dec425ac4f7aca1 = 
          (!fgallag_sel[2]) ? 
                       I6c9a443b704a7871ac13f164c1cdc88b: 
                       I76498f1e58ff35dc6153f76999f9f7a5;
              I11a9a93502a123a616205de5969bd5c8 = 
          (!fgallag_sel[2]) ? 
                       I200025a860f318f6ff9aaf89b146d16f: 
                       I107ae84d631e3a9574b62f4fdfe56140;
              I346c6ffdb07c9d7a5939fcd142871ef8 = 
          (!fgallag_sel[2]) ? 
                       Ief394bcabeb27c95f3dabe3d5c0bd643: 
                       Ibc52ae3742f657ac6abefd988494c8a1;
              I20fa0bb8e0dc75902328a349f0dca139 = 
          (!fgallag_sel[2]) ? 
                       I969ac5f2b8a9d6778300e3a91968ae4b: 
                       I3172be9cafebc7121994917ff35b25fb;
              Idb4bf6de8f078619ea6dcb51d8f7d329 = 
          (!fgallag_sel[2]) ? 
                       I388e0d1c3f421d7522d6c0521538693e: 
                       I0fa0bdc864c6173b380c763cf3e794ba;
              I8d2f1e18f0064f50176caa84061bf7ec = 
          (!fgallag_sel[2]) ? 
                       I9d6dc129ad747412224b487c4973db3a: 
                       Ic1c5ee07ecd5c9fc9c2c1f9c33cdca08;
              Ic48ab17819fe5de2326e4fcb0a1e84c2 = 
          (!fgallag_sel[2]) ? 
                       I1b2ba3544e2d26b40edbfaedf137812b: 
                       Ieb654d27e0306c60cd9eff05f4be76ca;
              If7332a4a9a6924d2fcbd0af70ecc0d1b = 
          (!fgallag_sel[2]) ? 
                       I462601141783fc299a3b081023233a56: 
                       I4e4e1489c822058cf54782c75c8d6996;
              I65a8d4181ad1817636600b816f41158b = 
          (!fgallag_sel[2]) ? 
                       I361a262df08182fcb917b7aa7aa73465: 
                       Ic8092176d020f45ae84ae72da9ea20a8;
              I746285d851cff1339ce0b99930415c2b = 
          (!fgallag_sel[2]) ? 
                       I361a7201d61113929f346f8b22ac01ef: 
                       I616e26bab7d9ada350f152cce0ac3569;
              I3305daafd6c3dc6ceb95673b361f0480 = 
          (!fgallag_sel[2]) ? 
                       I7cb33be246a06045ff19436b47ccfdca: 
                       Ic5aad088ddcc97dd7a3c8244a27a288e;
              I68babd78d3c2b1d6a064b25a3abd690e = 
          (!fgallag_sel[2]) ? 
                       I79c0e02b51ed3b20ca6de475189b6a48: 
                       I059966174241b59374640dc43018c49c;
              I9e7d989a414d752920fd69ac7c23ca38 = 
          (!fgallag_sel[2]) ? 
                       I1b43d5eb392150245e2a303582b9226f: 
                       Icc5e7d899df8ec350f804c1f32b9fe72;
              Ibf1b1639efba4277e759d747abe85e6b = 
          (!fgallag_sel[2]) ? 
                       I2f8fbab2b60878195ae8b2e1c0ff1208: 
                       I30e9a6bb0816599ede1e93a3091a572c;
               If67570ab71fa30823c9fe1277f35c1fe =  I815a192d304aedca5f772d6bd401ad3f ;
               Ia660cf2aa760392654bbc61cb60d9920 =  I83ce7e2b4c276008c33a5703eba16572 ;
              I2bf7c2dabc30d2207f04e0f6970f2287 = 
          (!fgallag_sel[2]) ? 
                       I984e48eb72dcef91797c57289ba1322e: 
                       I8a0f063aab90c7f50f8eff7e3626483d;
              I75c6cf6f3378e1377047d467a7e827f7 = 
          (!fgallag_sel[2]) ? 
                       Ia49e2201160f9da0d475b16d22efcac1: 
                       I59718bd7f0e7a0c9d63a038f2cb9d3eb;
               Ic3dacf077252960c863e8ec1a880f313 =  I7e703dc56c5c5604eb8e7ed32fd6ce78 ;
              I781a85002cfeb3038120fe37047710bc = 
          (!fgallag_sel[2]) ? 
                       If3582b232dccd45a4f3c07514062003c: 
                       I79a9448f1efc66a407e2dcc243638e6f;
               I0e8936dc5acf0e7c165d76a8b58f2765 =  I57fb6daf7238618d7ce10989a7f41025 ;
               I24b498fb5b12c3d4a5c7c9e36be4baf7 =  I629cd82c8226c17eb439cd2ad664a3b7 ;
              Id33f743a90e9f61fd4267c72442a98fa = 
          (!fgallag_sel[2]) ? 
                       Ida422d40a8abb52f4c78b63807f0ef16: 
                       Ic91b7435580f54bb1e3ffa6ea1b21f69;
               I6423dda227b49522f0d8d79fbfe32ecb =  Id1651e9d3e909ddb1f3779b4129713fd ;
               I6d8b1a2ff9d9d4a659ddd018a5ce1ebb =  I81c0a5fad7512ba9d8537018d6df2c23 ;
               I591484046d2f6f71badbd09db2dd16bc =  Ia6503d131655b73ae90b5553d116e92b ;
              Ibd503cf61b9c2e244852302f6ecbfb49 = 
          (!fgallag_sel[2]) ? 
                       I2c197653e4a8776ad3539f95aff27df5: 
                       I0d6cfa3166445e1396871afad62fba40;
               I42c86c7d63e8f622277ad4cd492dd142 =  Ie597ab8c4dd174055b4bda8dbdec0dd3 ;
               I480e64694b2be630cf58cb8d35e978eb =  I9426c6803cf8c7c6dbc422989eef5380 ;
               I0b029a353bcf76708510cbd17e96da2a =  I947d66b22e42c68930e8bf7d1439a376 ;
               I8d0c242b4c0b43f6d1f3796ae1a1be58 =  I22715ee56f34e2c7cfdae2dd409ac653 ;
               I71e27087daf4bc19fb7e5851935a31e9 =  Id2e3d5dfe5c8ec9128f5a719175c0f35 ;
               Ieff0a4b462cd624e967db20434f0452d =  I0f1ace68f720dfcca74605ec277d0067 ;
               I835c19cffb04dfb43ef7c362c7a9cea0 =  Ia10e05a72a5d3c1e16b99510e94f6121 ;
               Ic506210a4fc9ec0b663ed4a364951fbf =  I8b6f4ea7a19f4b359aa01867c4502ccf ;
              I409f55664c78aaefc044bebb7177392a = 
          (!fgallag_sel[2]) ? 
                       I323124e6fcbab5bdda4bd24c7b2a99c1: 
                       Ib943a483749ffc791a5965ed0840bb0f;
               I9477257b731d59c02213efd459153ea3 =  0;
