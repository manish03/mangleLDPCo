parameter n_minus_m = 'd40;
parameter n_int = 'd208;
parameter m_int = 'd168;



parameter z_int = 'd4;



wire Ia754e5a85bf385f490ebf0d576feded059b06ce14d403f7c4089d1580e192a79; 
assign Ia754e5a85bf385f490ebf0d576feded059b06ce14d403f7c4089d1580e192a79 = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[14] ^ 
        y_nr_in[25] ^ 
        y_nr_in[37] ^ 
0; 



wire I3be0bcc6f2bc65a276fdbf66ebeb0e44bed6099c32a0a9139be3255f0fa0bd7f; 
assign I3be0bcc6f2bc65a276fdbf66ebeb0e44bed6099c32a0a9139be3255f0fa0bd7f = 
        y_nr_in[40] ^ 
        y_nr_in[44] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[0] = 
Ia754e5a85bf385f490ebf0d576feded059b06ce14d403f7c4089d1580e192a79 ^ 
I3be0bcc6f2bc65a276fdbf66ebeb0e44bed6099c32a0a9139be3255f0fa0bd7f ^ 
0; 



wire I43eb78046b932ed5dcde60580cefe0936670786312795b57786877d9ff921559; 
assign I43eb78046b932ed5dcde60580cefe0936670786312795b57786877d9ff921559 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[15] ^ 
        y_nr_in[26] ^ 
        y_nr_in[38] ^ 
0; 



wire Ida43fa065b7b213eb3b72000fbea9c5a47a29c9aa05f8b31b014bb1844564354; 
assign Ida43fa065b7b213eb3b72000fbea9c5a47a29c9aa05f8b31b014bb1844564354 = 
        y_nr_in[41] ^ 
        y_nr_in[45] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[1] = 
I43eb78046b932ed5dcde60580cefe0936670786312795b57786877d9ff921559 ^ 
Ida43fa065b7b213eb3b72000fbea9c5a47a29c9aa05f8b31b014bb1844564354 ^ 
0; 



wire I2d365e84eb318249e8c3b26245554f4163f428d85d6a75b2ab7d272e425197b6; 
assign I2d365e84eb318249e8c3b26245554f4163f428d85d6a75b2ab7d272e425197b6 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[12] ^ 
        y_nr_in[27] ^ 
        y_nr_in[39] ^ 
0; 



wire I97671fa85bef5c41f114b83f918078fd41c22e6c035c9977f72a5107a11ceeba; 
assign I97671fa85bef5c41f114b83f918078fd41c22e6c035c9977f72a5107a11ceeba = 
        y_nr_in[42] ^ 
        y_nr_in[46] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[2] = 
I2d365e84eb318249e8c3b26245554f4163f428d85d6a75b2ab7d272e425197b6 ^ 
I97671fa85bef5c41f114b83f918078fd41c22e6c035c9977f72a5107a11ceeba ^ 
0; 



wire I234474e73bd3f6362909548815d18f613ab8f5ded2cd2b548306f95dbb997b58; 
assign I234474e73bd3f6362909548815d18f613ab8f5ded2cd2b548306f95dbb997b58 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[13] ^ 
        y_nr_in[24] ^ 
        y_nr_in[36] ^ 
0; 



wire I57e0c6461a17a491b5ad66423d595a11842358c61edc9f42415b3476b2c8df9a; 
assign I57e0c6461a17a491b5ad66423d595a11842358c61edc9f42415b3476b2c8df9a = 
        y_nr_in[43] ^ 
        y_nr_in[47] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[3] = 
I234474e73bd3f6362909548815d18f613ab8f5ded2cd2b548306f95dbb997b58 ^ 
I57e0c6461a17a491b5ad66423d595a11842358c61edc9f42415b3476b2c8df9a ^ 
0; 



wire I464a66a04ca267b8ad18ecafd37dedb2ea825b06da339aaeb552e3b4f11b213c; 
assign I464a66a04ca267b8ad18ecafd37dedb2ea825b06da339aaeb552e3b4f11b213c = 
        y_nr_in[3] ^ 
        y_nr_in[14] ^ 
        y_nr_in[17] ^ 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
0; 



wire Ia20a88826b86f8b2c06ce04d767e24364184eee021f1e1bc75608b967d4bb2d6; 
assign Ia20a88826b86f8b2c06ce04d767e24364184eee021f1e1bc75608b967d4bb2d6 = 
        y_nr_in[28] ^ 
        y_nr_in[32] ^ 
        y_nr_in[36] ^ 
        y_nr_in[44] ^ 
        y_nr_in[48] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[4] = 
I464a66a04ca267b8ad18ecafd37dedb2ea825b06da339aaeb552e3b4f11b213c ^ 
Ia20a88826b86f8b2c06ce04d767e24364184eee021f1e1bc75608b967d4bb2d6 ^ 
0; 



wire I27a077b80a3e5b8e3ae31d889453301cd92985b3f6aa3b3b83cc147f3fef419e; 
assign I27a077b80a3e5b8e3ae31d889453301cd92985b3f6aa3b3b83cc147f3fef419e = 
        y_nr_in[0] ^ 
        y_nr_in[15] ^ 
        y_nr_in[18] ^ 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
0; 



wire Ib11b9ebf95e1ad7a5170d9141aca75f5119b5d6e51d0caf66f645ca233c0fec3; 
assign Ib11b9ebf95e1ad7a5170d9141aca75f5119b5d6e51d0caf66f645ca233c0fec3 = 
        y_nr_in[29] ^ 
        y_nr_in[33] ^ 
        y_nr_in[37] ^ 
        y_nr_in[45] ^ 
        y_nr_in[49] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[5] = 
I27a077b80a3e5b8e3ae31d889453301cd92985b3f6aa3b3b83cc147f3fef419e ^ 
Ib11b9ebf95e1ad7a5170d9141aca75f5119b5d6e51d0caf66f645ca233c0fec3 ^ 
0; 



wire I7f2aff8cdf25be8cf51631b3d98ffd590dff21fcb0a7696325e448082ecce2e5; 
assign I7f2aff8cdf25be8cf51631b3d98ffd590dff21fcb0a7696325e448082ecce2e5 = 
        y_nr_in[1] ^ 
        y_nr_in[12] ^ 
        y_nr_in[19] ^ 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
0; 



wire Ia208a631318cc08061a6e7060a645efaf2a532420dd44f900c03059ba0666fa7; 
assign Ia208a631318cc08061a6e7060a645efaf2a532420dd44f900c03059ba0666fa7 = 
        y_nr_in[30] ^ 
        y_nr_in[34] ^ 
        y_nr_in[38] ^ 
        y_nr_in[46] ^ 
        y_nr_in[50] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[6] = 
I7f2aff8cdf25be8cf51631b3d98ffd590dff21fcb0a7696325e448082ecce2e5 ^ 
Ia208a631318cc08061a6e7060a645efaf2a532420dd44f900c03059ba0666fa7 ^ 
0; 



wire I1c3e84d05fc731c6c716c6dd83c7eb1bb762db24e5a8546740d8e2379bf5dfce; 
assign I1c3e84d05fc731c6c716c6dd83c7eb1bb762db24e5a8546740d8e2379bf5dfce = 
        y_nr_in[2] ^ 
        y_nr_in[13] ^ 
        y_nr_in[16] ^ 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
0; 



wire Ifde25f01fd269278c9805cf2b5fc58f2c677698ea9b77153c9c899f011259230; 
assign Ifde25f01fd269278c9805cf2b5fc58f2c677698ea9b77153c9c899f011259230 = 
        y_nr_in[31] ^ 
        y_nr_in[35] ^ 
        y_nr_in[39] ^ 
        y_nr_in[47] ^ 
        y_nr_in[51] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[7] = 
I1c3e84d05fc731c6c716c6dd83c7eb1bb762db24e5a8546740d8e2379bf5dfce ^ 
Ifde25f01fd269278c9805cf2b5fc58f2c677698ea9b77153c9c899f011259230 ^ 
0; 



wire If22ec55e24855fe5b350302d7379bcbbd65d25fd1617cc25db73a594340a76e8; 
assign If22ec55e24855fe5b350302d7379bcbbd65d25fd1617cc25db73a594340a76e8 = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[12] ^ 
        y_nr_in[16] ^ 
        y_nr_in[32] ^ 
0; 



wire I66d3686f1cafbd0abebf237dd1a739191a3a36c38cb85e76cf1f0e511920b0cb; 
assign I66d3686f1cafbd0abebf237dd1a739191a3a36c38cb85e76cf1f0e511920b0cb = 
        y_nr_in[41] ^ 
        y_nr_in[48] ^ 
        y_nr_in[52] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[8] = 
If22ec55e24855fe5b350302d7379bcbbd65d25fd1617cc25db73a594340a76e8 ^ 
I66d3686f1cafbd0abebf237dd1a739191a3a36c38cb85e76cf1f0e511920b0cb ^ 
0; 



wire I990b3bb764321c1d509cc0c72b23d030d9b67d1d06c0a89b644d044708534d17; 
assign I990b3bb764321c1d509cc0c72b23d030d9b67d1d06c0a89b644d044708534d17 = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[13] ^ 
        y_nr_in[17] ^ 
        y_nr_in[33] ^ 
0; 



wire Ia2146d2d8404e6c1b15586909b91158aca8d5ba0e988c20929bc43d7b732cfe8; 
assign Ia2146d2d8404e6c1b15586909b91158aca8d5ba0e988c20929bc43d7b732cfe8 = 
        y_nr_in[42] ^ 
        y_nr_in[49] ^ 
        y_nr_in[53] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[9] = 
I990b3bb764321c1d509cc0c72b23d030d9b67d1d06c0a89b644d044708534d17 ^ 
Ia2146d2d8404e6c1b15586909b91158aca8d5ba0e988c20929bc43d7b732cfe8 ^ 
0; 



wire Ifd1816d795539a639bc67803af6786c22106e4fd77f438194b61b8d9bcd7cf63; 
assign Ifd1816d795539a639bc67803af6786c22106e4fd77f438194b61b8d9bcd7cf63 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[14] ^ 
        y_nr_in[18] ^ 
        y_nr_in[34] ^ 
0; 



wire I322acff95ca02447826f9ce862c8f437cd2ec4028205b675fd3f924baa7af076; 
assign I322acff95ca02447826f9ce862c8f437cd2ec4028205b675fd3f924baa7af076 = 
        y_nr_in[43] ^ 
        y_nr_in[50] ^ 
        y_nr_in[54] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[10] = 
Ifd1816d795539a639bc67803af6786c22106e4fd77f438194b61b8d9bcd7cf63 ^ 
I322acff95ca02447826f9ce862c8f437cd2ec4028205b675fd3f924baa7af076 ^ 
0; 



wire Icf82b42a4b0f156400a64d186eb21b5b5b9f55927e68652afc452b0b355bc492; 
assign Icf82b42a4b0f156400a64d186eb21b5b5b9f55927e68652afc452b0b355bc492 = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[15] ^ 
        y_nr_in[19] ^ 
        y_nr_in[35] ^ 
0; 



wire I459874acad7ca256bdfdc44ad913a9e869e5cecf70a57fc7ed14aa87d87720b3; 
assign I459874acad7ca256bdfdc44ad913a9e869e5cecf70a57fc7ed14aa87d87720b3 = 
        y_nr_in[40] ^ 
        y_nr_in[51] ^ 
        y_nr_in[55] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[11] = 
Icf82b42a4b0f156400a64d186eb21b5b5b9f55927e68652afc452b0b355bc492 ^ 
I459874acad7ca256bdfdc44ad913a9e869e5cecf70a57fc7ed14aa87d87720b3 ^ 
0; 



wire I0025fb037fe0328fd006b99bdb62b02be917ae1e32e4740e9358eb2606a63f28; 
assign I0025fb037fe0328fd006b99bdb62b02be917ae1e32e4740e9358eb2606a63f28 = 
        y_nr_in[4] ^ 
        y_nr_in[10] ^ 
        y_nr_in[18] ^ 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
0; 



wire I70cd9e43dc757d9e39bd65b1b08a0542c2d724f18fd2699e304072753ef64d41; 
assign I70cd9e43dc757d9e39bd65b1b08a0542c2d724f18fd2699e304072753ef64d41 = 
        y_nr_in[30] ^ 
        y_nr_in[34] ^ 
        y_nr_in[36] ^ 
        y_nr_in[40] ^ 
        y_nr_in[52] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[12] = 
I0025fb037fe0328fd006b99bdb62b02be917ae1e32e4740e9358eb2606a63f28 ^ 
I70cd9e43dc757d9e39bd65b1b08a0542c2d724f18fd2699e304072753ef64d41 ^ 
0; 



wire I3ed5de6723367de0aa5ce5e8529765dbec20f386853f551e2663231c0bea9b77; 
assign I3ed5de6723367de0aa5ce5e8529765dbec20f386853f551e2663231c0bea9b77 = 
        y_nr_in[5] ^ 
        y_nr_in[11] ^ 
        y_nr_in[19] ^ 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
0; 



wire I1ace09c863e6485120dffa1ee2426188b7bc7a46649748e5cbcbba75c283146d; 
assign I1ace09c863e6485120dffa1ee2426188b7bc7a46649748e5cbcbba75c283146d = 
        y_nr_in[31] ^ 
        y_nr_in[35] ^ 
        y_nr_in[37] ^ 
        y_nr_in[41] ^ 
        y_nr_in[53] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[13] = 
I3ed5de6723367de0aa5ce5e8529765dbec20f386853f551e2663231c0bea9b77 ^ 
I1ace09c863e6485120dffa1ee2426188b7bc7a46649748e5cbcbba75c283146d ^ 
0; 



wire I3b3784bd62023713306693cdf60f43b969345e335321dd179448b141dbc25ca6; 
assign I3b3784bd62023713306693cdf60f43b969345e335321dd179448b141dbc25ca6 = 
        y_nr_in[6] ^ 
        y_nr_in[8] ^ 
        y_nr_in[16] ^ 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
0; 



wire I3342b099665f88eb8886eb01013b7d43cc689a88148819cf07fe3e3844bf1921; 
assign I3342b099665f88eb8886eb01013b7d43cc689a88148819cf07fe3e3844bf1921 = 
        y_nr_in[28] ^ 
        y_nr_in[32] ^ 
        y_nr_in[38] ^ 
        y_nr_in[42] ^ 
        y_nr_in[54] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[14] = 
I3b3784bd62023713306693cdf60f43b969345e335321dd179448b141dbc25ca6 ^ 
I3342b099665f88eb8886eb01013b7d43cc689a88148819cf07fe3e3844bf1921 ^ 
0; 



wire I923cb17b12cd045b6167b98137ae46f48394c83d7864bc1fc5e795525104cef5; 
assign I923cb17b12cd045b6167b98137ae46f48394c83d7864bc1fc5e795525104cef5 = 
        y_nr_in[7] ^ 
        y_nr_in[9] ^ 
        y_nr_in[17] ^ 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
0; 



wire I219446b1d1ace1b2d1ca60901fe5c3c4982db52b01ee4877d78babb63e3c77e7; 
assign I219446b1d1ace1b2d1ca60901fe5c3c4982db52b01ee4877d78babb63e3c77e7 = 
        y_nr_in[29] ^ 
        y_nr_in[33] ^ 
        y_nr_in[39] ^ 
        y_nr_in[43] ^ 
        y_nr_in[55] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[15] = 
I923cb17b12cd045b6167b98137ae46f48394c83d7864bc1fc5e795525104cef5 ^ 
I219446b1d1ace1b2d1ca60901fe5c3c4982db52b01ee4877d78babb63e3c77e7 ^ 
0; 



wire I8dec0a083eb5938cf56f2752f80e9248cb5d7f6964451857436507d148ca5b38; 
assign I8dec0a083eb5938cf56f2752f80e9248cb5d7f6964451857436507d148ca5b38 = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[47] ^ 
        y_nr_in[56] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[16] = 
I8dec0a083eb5938cf56f2752f80e9248cb5d7f6964451857436507d148ca5b38 ^ 
0; 



wire Idd28fae575f06f4648e8061f79b63200ddf252fbe5e25f399b3a111b92e5fb71; 
assign Idd28fae575f06f4648e8061f79b63200ddf252fbe5e25f399b3a111b92e5fb71 = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[44] ^ 
        y_nr_in[57] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[17] = 
Idd28fae575f06f4648e8061f79b63200ddf252fbe5e25f399b3a111b92e5fb71 ^ 
0; 



wire I7eb73a233c8d98da5a99de909bdb6480edf8d999b9093c62f1c956faea0ea933; 
assign I7eb73a233c8d98da5a99de909bdb6480edf8d999b9093c62f1c956faea0ea933 = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[45] ^ 
        y_nr_in[58] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[18] = 
I7eb73a233c8d98da5a99de909bdb6480edf8d999b9093c62f1c956faea0ea933 ^ 
0; 



wire I9d3c7bd7f2dc6b382f3fdf5e73d847f6c410b5d3e0cef2dc49f9ecba7d88a885; 
assign I9d3c7bd7f2dc6b382f3fdf5e73d847f6c410b5d3e0cef2dc49f9ecba7d88a885 = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[46] ^ 
        y_nr_in[59] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[19] = 
I9d3c7bd7f2dc6b382f3fdf5e73d847f6c410b5d3e0cef2dc49f9ecba7d88a885 ^ 
0; 



wire I465831cf3e551297bf4782c528acda2233762f5176c7b0d5674c409b6f22a4c9; 
assign I465831cf3e551297bf4782c528acda2233762f5176c7b0d5674c409b6f22a4c9 = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[47] ^ 
0; 



wire I0e698d845c730cab5871d5f0cd00937e17460acf945a9d50ff1188dafa145142; 
assign I0e698d845c730cab5871d5f0cd00937e17460acf945a9d50ff1188dafa145142 = 
        y_nr_in[60] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[20] = 
I465831cf3e551297bf4782c528acda2233762f5176c7b0d5674c409b6f22a4c9 ^ 
I0e698d845c730cab5871d5f0cd00937e17460acf945a9d50ff1188dafa145142 ^ 
0; 



wire I0f58d8c06829583b44d0dd3808efd6d42dfb535e6bf3aca181dbec2ab36a001e; 
assign I0f58d8c06829583b44d0dd3808efd6d42dfb535e6bf3aca181dbec2ab36a001e = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[44] ^ 
0; 



wire I0da36b1fc93eb32d0a163d9228207db2d0a233a748e8ca70e9b5cd02df118581; 
assign I0da36b1fc93eb32d0a163d9228207db2d0a233a748e8ca70e9b5cd02df118581 = 
        y_nr_in[61] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[21] = 
I0f58d8c06829583b44d0dd3808efd6d42dfb535e6bf3aca181dbec2ab36a001e ^ 
I0da36b1fc93eb32d0a163d9228207db2d0a233a748e8ca70e9b5cd02df118581 ^ 
0; 



wire Idef21594a072095d16deed7ab8e5f3658ddeb8f1a78e6dd4daffddde27dd9aaf; 
assign Idef21594a072095d16deed7ab8e5f3658ddeb8f1a78e6dd4daffddde27dd9aaf = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[45] ^ 
0; 



wire I0fa5be3d161015811a84fe165c4d98646a3af7a95b6a0c31e0a8a6a05c2a0ca7; 
assign I0fa5be3d161015811a84fe165c4d98646a3af7a95b6a0c31e0a8a6a05c2a0ca7 = 
        y_nr_in[62] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[22] = 
Idef21594a072095d16deed7ab8e5f3658ddeb8f1a78e6dd4daffddde27dd9aaf ^ 
I0fa5be3d161015811a84fe165c4d98646a3af7a95b6a0c31e0a8a6a05c2a0ca7 ^ 
0; 



wire Iaf351feee0df3dc4ea65f211033f2fd55674b9811c2ab9ef961935bc460105e2; 
assign Iaf351feee0df3dc4ea65f211033f2fd55674b9811c2ab9ef961935bc460105e2 = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[46] ^ 
0; 



wire Ie6abf919a65099df3d347445f21e4b69fa490b46bdb6b84a8f1a350e41dd8aa5; 
assign Ie6abf919a65099df3d347445f21e4b69fa490b46bdb6b84a8f1a350e41dd8aa5 = 
        y_nr_in[63] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[23] = 
Iaf351feee0df3dc4ea65f211033f2fd55674b9811c2ab9ef961935bc460105e2 ^ 
Ie6abf919a65099df3d347445f21e4b69fa490b46bdb6b84a8f1a350e41dd8aa5 ^ 
0; 



wire I4f8fc161be410cc37bd9fd5a0afb47551fdbcae4134b83e971e9da3a45d213af; 
assign I4f8fc161be410cc37bd9fd5a0afb47551fdbcae4134b83e971e9da3a45d213af = 
        y_nr_in[3] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
0; 



wire Iafd9234450bab42febd01667ab527105103d5177775f4664793f1912e7fe86dd; 
assign Iafd9234450bab42febd01667ab527105103d5177775f4664793f1912e7fe86dd = 
        y_nr_in[64] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[24] = 
I4f8fc161be410cc37bd9fd5a0afb47551fdbcae4134b83e971e9da3a45d213af ^ 
Iafd9234450bab42febd01667ab527105103d5177775f4664793f1912e7fe86dd ^ 
0; 



wire I8829f524a53813761534199990a3f97a98546986b5cd6d986e17fc9b46b42f69; 
assign I8829f524a53813761534199990a3f97a98546986b5cd6d986e17fc9b46b42f69 = 
        y_nr_in[0] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
0; 



wire I10b2088839c749fdb1549aacb4301d2d4fde02c184628ce338488245c70f36a9; 
assign I10b2088839c749fdb1549aacb4301d2d4fde02c184628ce338488245c70f36a9 = 
        y_nr_in[65] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[25] = 
I8829f524a53813761534199990a3f97a98546986b5cd6d986e17fc9b46b42f69 ^ 
I10b2088839c749fdb1549aacb4301d2d4fde02c184628ce338488245c70f36a9 ^ 
0; 



wire I07cdc26d3bcc2abb3a2c1044967c758acf438c8eb603cddaf4e6706cbfaaca76; 
assign I07cdc26d3bcc2abb3a2c1044967c758acf438c8eb603cddaf4e6706cbfaaca76 = 
        y_nr_in[1] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
0; 



wire I5b916e6d8ff79e034ebd7897cbdbc51d8e9551af827b4d49695968ff1e76620e; 
assign I5b916e6d8ff79e034ebd7897cbdbc51d8e9551af827b4d49695968ff1e76620e = 
        y_nr_in[66] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[26] = 
I07cdc26d3bcc2abb3a2c1044967c758acf438c8eb603cddaf4e6706cbfaaca76 ^ 
I5b916e6d8ff79e034ebd7897cbdbc51d8e9551af827b4d49695968ff1e76620e ^ 
0; 



wire I6faac169f65e2558009cd753e7daef5377ce29ca4004633548b4d4258493f6e2; 
assign I6faac169f65e2558009cd753e7daef5377ce29ca4004633548b4d4258493f6e2 = 
        y_nr_in[2] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
0; 



wire I82761f460ae8fff7e20d1c832724e43f81e3b68a2fa868a6db67960c9fe96f08; 
assign I82761f460ae8fff7e20d1c832724e43f81e3b68a2fa868a6db67960c9fe96f08 = 
        y_nr_in[67] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[27] = 
I6faac169f65e2558009cd753e7daef5377ce29ca4004633548b4d4258493f6e2 ^ 
I82761f460ae8fff7e20d1c832724e43f81e3b68a2fa868a6db67960c9fe96f08 ^ 
0; 



wire I39a74d1f0272013a93cac8b11f5843c80c1dde371a39f87475f75074362c9fe6; 
assign I39a74d1f0272013a93cac8b11f5843c80c1dde371a39f87475f75074362c9fe6 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[47] ^ 
        y_nr_in[52] ^ 
0; 



wire I4c06a0d9de5bda0f9a26d71a97008a9ab7ba84cbb5e402fa46c931782d5e2185; 
assign I4c06a0d9de5bda0f9a26d71a97008a9ab7ba84cbb5e402fa46c931782d5e2185 = 
        y_nr_in[68] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[28] = 
I39a74d1f0272013a93cac8b11f5843c80c1dde371a39f87475f75074362c9fe6 ^ 
I4c06a0d9de5bda0f9a26d71a97008a9ab7ba84cbb5e402fa46c931782d5e2185 ^ 
0; 



wire I95dc040aca47aac6019183871fcf94ea461de319fcf026dad03200e646057e79; 
assign I95dc040aca47aac6019183871fcf94ea461de319fcf026dad03200e646057e79 = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[44] ^ 
        y_nr_in[53] ^ 
0; 



wire Ifb0a16cf41977e063e3af64e7523cfd236ba29a1437c3b28e5317926411be138; 
assign Ifb0a16cf41977e063e3af64e7523cfd236ba29a1437c3b28e5317926411be138 = 
        y_nr_in[69] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[29] = 
I95dc040aca47aac6019183871fcf94ea461de319fcf026dad03200e646057e79 ^ 
Ifb0a16cf41977e063e3af64e7523cfd236ba29a1437c3b28e5317926411be138 ^ 
0; 



wire Ic19fb6228809fd624a696e8f80118bad758b8f09a0f9a29d3327c07a386cdf3b; 
assign Ic19fb6228809fd624a696e8f80118bad758b8f09a0f9a29d3327c07a386cdf3b = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[45] ^ 
        y_nr_in[54] ^ 
0; 



wire I51ebfe4eda50ec6c153247b5ffa66b33f2fb3376686d900e210a7ec6d519d72c; 
assign I51ebfe4eda50ec6c153247b5ffa66b33f2fb3376686d900e210a7ec6d519d72c = 
        y_nr_in[70] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[30] = 
Ic19fb6228809fd624a696e8f80118bad758b8f09a0f9a29d3327c07a386cdf3b ^ 
I51ebfe4eda50ec6c153247b5ffa66b33f2fb3376686d900e210a7ec6d519d72c ^ 
0; 



wire I6df3297499ed45f2bf9081d4e38845ba7ccbc93238350c4396e050b316c85c92; 
assign I6df3297499ed45f2bf9081d4e38845ba7ccbc93238350c4396e050b316c85c92 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[46] ^ 
        y_nr_in[55] ^ 
0; 



wire Id22ea28516b2ffff1ce82b04fa3d1e1c1d3c084ba87f5cffc8fa1c1a85f7f3a2; 
assign Id22ea28516b2ffff1ce82b04fa3d1e1c1d3c084ba87f5cffc8fa1c1a85f7f3a2 = 
        y_nr_in[71] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[31] = 
I6df3297499ed45f2bf9081d4e38845ba7ccbc93238350c4396e050b316c85c92 ^ 
Id22ea28516b2ffff1ce82b04fa3d1e1c1d3c084ba87f5cffc8fa1c1a85f7f3a2 ^ 
0; 



wire If8b3c7cf476024de27e03f04c41c46cf30e76c85f88932d37f178ca5c7a7a729; 
assign If8b3c7cf476024de27e03f04c41c46cf30e76c85f88932d37f178ca5c7a7a729 = 
        y_nr_in[2] ^ 
        y_nr_in[6] ^ 
        y_nr_in[50] ^ 
        y_nr_in[72] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[32] = 
If8b3c7cf476024de27e03f04c41c46cf30e76c85f88932d37f178ca5c7a7a729 ^ 
0; 



wire I9ab3812757676189077c2e66b767871e00523eb3c397aa01786ce06be77a46c9; 
assign I9ab3812757676189077c2e66b767871e00523eb3c397aa01786ce06be77a46c9 = 
        y_nr_in[3] ^ 
        y_nr_in[7] ^ 
        y_nr_in[51] ^ 
        y_nr_in[73] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[33] = 
I9ab3812757676189077c2e66b767871e00523eb3c397aa01786ce06be77a46c9 ^ 
0; 



wire Ie516174657b0c601af7358d7239e94070f6f943211e72cbdc52bc3434e6280dc; 
assign Ie516174657b0c601af7358d7239e94070f6f943211e72cbdc52bc3434e6280dc = 
        y_nr_in[0] ^ 
        y_nr_in[4] ^ 
        y_nr_in[48] ^ 
        y_nr_in[74] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[34] = 
Ie516174657b0c601af7358d7239e94070f6f943211e72cbdc52bc3434e6280dc ^ 
0; 



wire I584c4529f6a3af2fa71f6c2d32075ca11c70c4b43633693e93112dfac8fd72b8; 
assign I584c4529f6a3af2fa71f6c2d32075ca11c70c4b43633693e93112dfac8fd72b8 = 
        y_nr_in[1] ^ 
        y_nr_in[5] ^ 
        y_nr_in[49] ^ 
        y_nr_in[75] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[35] = 
I584c4529f6a3af2fa71f6c2d32075ca11c70c4b43633693e93112dfac8fd72b8 ^ 
0; 



wire I4c0a77b0b23f997a538698670497345f1280b0926567b0f918ae5bafc8a6cbd5; 
assign I4c0a77b0b23f997a538698670497345f1280b0926567b0f918ae5bafc8a6cbd5 = 
        y_nr_in[7] ^ 
        y_nr_in[33] ^ 
        y_nr_in[41] ^ 
        y_nr_in[47] ^ 
        y_nr_in[76] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[36] = 
I4c0a77b0b23f997a538698670497345f1280b0926567b0f918ae5bafc8a6cbd5 ^ 
0; 



wire Ic19cf72cd0de43be6152157c21418d3596f8e3ca4596d58147ca49babb30a844; 
assign Ic19cf72cd0de43be6152157c21418d3596f8e3ca4596d58147ca49babb30a844 = 
        y_nr_in[4] ^ 
        y_nr_in[34] ^ 
        y_nr_in[42] ^ 
        y_nr_in[44] ^ 
        y_nr_in[77] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[37] = 
Ic19cf72cd0de43be6152157c21418d3596f8e3ca4596d58147ca49babb30a844 ^ 
0; 



wire Iaa1af060da3a5b8d3e46149acc730ec7497c7018b078c1ba5e043f7380c82b99; 
assign Iaa1af060da3a5b8d3e46149acc730ec7497c7018b078c1ba5e043f7380c82b99 = 
        y_nr_in[5] ^ 
        y_nr_in[35] ^ 
        y_nr_in[43] ^ 
        y_nr_in[45] ^ 
        y_nr_in[78] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[38] = 
Iaa1af060da3a5b8d3e46149acc730ec7497c7018b078c1ba5e043f7380c82b99 ^ 
0; 



wire I3f8a7acd44f94bcf874351893389df2cf027fdb0e863e75fab3eade382c38359; 
assign I3f8a7acd44f94bcf874351893389df2cf027fdb0e863e75fab3eade382c38359 = 
        y_nr_in[6] ^ 
        y_nr_in[32] ^ 
        y_nr_in[40] ^ 
        y_nr_in[46] ^ 
        y_nr_in[79] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[39] = 
I3f8a7acd44f94bcf874351893389df2cf027fdb0e863e75fab3eade382c38359 ^ 
0; 



wire I05c283f93322c34c0e84af2cb01a12f0ee35062970d97fd23ee6b42ebe92cf5f; 
assign I05c283f93322c34c0e84af2cb01a12f0ee35062970d97fd23ee6b42ebe92cf5f = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[24] ^ 
        y_nr_in[29] ^ 
        y_nr_in[80] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[40] = 
I05c283f93322c34c0e84af2cb01a12f0ee35062970d97fd23ee6b42ebe92cf5f ^ 
0; 



wire I5dbc0e51b05c5c3d823e618842b9969236e729360fa86a98bf4ce7cc78b5eeb5; 
assign I5dbc0e51b05c5c3d823e618842b9969236e729360fa86a98bf4ce7cc78b5eeb5 = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[25] ^ 
        y_nr_in[30] ^ 
        y_nr_in[81] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[41] = 
I5dbc0e51b05c5c3d823e618842b9969236e729360fa86a98bf4ce7cc78b5eeb5 ^ 
0; 



wire I0386a557968a59dfcb5e451f17d9ce280ad8a2f8bbe31166d6732e9c5f677ec6; 
assign I0386a557968a59dfcb5e451f17d9ce280ad8a2f8bbe31166d6732e9c5f677ec6 = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[26] ^ 
        y_nr_in[31] ^ 
        y_nr_in[82] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[42] = 
I0386a557968a59dfcb5e451f17d9ce280ad8a2f8bbe31166d6732e9c5f677ec6 ^ 
0; 



wire Ib4d823cb59b99786fca9e5f03504ffa43c9f1cb1387cb092463d1f9bdf141c3e; 
assign Ib4d823cb59b99786fca9e5f03504ffa43c9f1cb1387cb092463d1f9bdf141c3e = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[27] ^ 
        y_nr_in[28] ^ 
        y_nr_in[83] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[43] = 
Ib4d823cb59b99786fca9e5f03504ffa43c9f1cb1387cb092463d1f9bdf141c3e ^ 
0; 



wire I61011f0b1416d657724b0c249ea6daac420b93d98dd3b993980b0edf3c416fe2; 
assign I61011f0b1416d657724b0c249ea6daac420b93d98dd3b993980b0edf3c416fe2 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[38] ^ 
        y_nr_in[52] ^ 
        y_nr_in[84] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[44] = 
I61011f0b1416d657724b0c249ea6daac420b93d98dd3b993980b0edf3c416fe2 ^ 
0; 



wire I30d79dc675d50733335c0411e487183ac122b0adee90342bbdf6b24b367bd50d; 
assign I30d79dc675d50733335c0411e487183ac122b0adee90342bbdf6b24b367bd50d = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[39] ^ 
        y_nr_in[53] ^ 
        y_nr_in[85] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[45] = 
I30d79dc675d50733335c0411e487183ac122b0adee90342bbdf6b24b367bd50d ^ 
0; 



wire I0c281815ff5350e31934a28187719345d95cfc01af21065419880e555a89e18c; 
assign I0c281815ff5350e31934a28187719345d95cfc01af21065419880e555a89e18c = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[36] ^ 
        y_nr_in[54] ^ 
        y_nr_in[86] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[46] = 
I0c281815ff5350e31934a28187719345d95cfc01af21065419880e555a89e18c ^ 
0; 



wire Ia8a1fd0bc936c264f84030aebee2a8cef11a8ca27f206d541bf906d778935075; 
assign Ia8a1fd0bc936c264f84030aebee2a8cef11a8ca27f206d541bf906d778935075 = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[37] ^ 
        y_nr_in[55] ^ 
        y_nr_in[87] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[47] = 
Ia8a1fd0bc936c264f84030aebee2a8cef11a8ca27f206d541bf906d778935075 ^ 
0; 



wire I2965d0c53d0db4fc12bd1b2158c1506b45b6f3dba342aaf35f9f826335927a4f; 
assign I2965d0c53d0db4fc12bd1b2158c1506b45b6f3dba342aaf35f9f826335927a4f = 
        y_nr_in[7] ^ 
        y_nr_in[15] ^ 
        y_nr_in[46] ^ 
        y_nr_in[88] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[48] = 
I2965d0c53d0db4fc12bd1b2158c1506b45b6f3dba342aaf35f9f826335927a4f ^ 
0; 



wire I0e3c5a96f4e9f85270523d54df7163937f6d95f9b24ff4985e81426ec488fc7e; 
assign I0e3c5a96f4e9f85270523d54df7163937f6d95f9b24ff4985e81426ec488fc7e = 
        y_nr_in[4] ^ 
        y_nr_in[12] ^ 
        y_nr_in[47] ^ 
        y_nr_in[89] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[49] = 
I0e3c5a96f4e9f85270523d54df7163937f6d95f9b24ff4985e81426ec488fc7e ^ 
0; 



wire I539e4b9f773ad2804f34f50cdb1511a465ad3ff410d95d0f9e5fc417213f02c1; 
assign I539e4b9f773ad2804f34f50cdb1511a465ad3ff410d95d0f9e5fc417213f02c1 = 
        y_nr_in[5] ^ 
        y_nr_in[13] ^ 
        y_nr_in[44] ^ 
        y_nr_in[90] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[50] = 
I539e4b9f773ad2804f34f50cdb1511a465ad3ff410d95d0f9e5fc417213f02c1 ^ 
0; 



wire I0e7f1e063308ec29231be6dd166e266fee924483693a44e5d1d42429bf900794; 
assign I0e7f1e063308ec29231be6dd166e266fee924483693a44e5d1d42429bf900794 = 
        y_nr_in[6] ^ 
        y_nr_in[14] ^ 
        y_nr_in[45] ^ 
        y_nr_in[91] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[51] = 
I0e7f1e063308ec29231be6dd166e266fee924483693a44e5d1d42429bf900794 ^ 
0; 



wire I1c1ec23b94c8f0835a9f410a0598716b00ca1f5bb1c52aa9f6f03eb7cfdca0aa; 
assign I1c1ec23b94c8f0835a9f410a0598716b00ca1f5bb1c52aa9f6f03eb7cfdca0aa = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[34] ^ 
        y_nr_in[54] ^ 
        y_nr_in[92] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[52] = 
I1c1ec23b94c8f0835a9f410a0598716b00ca1f5bb1c52aa9f6f03eb7cfdca0aa ^ 
0; 



wire I15397ad3270aed0ea90a6a9aedf0a2269cda3b415eaa4b3f79522bc3d0ed209e; 
assign I15397ad3270aed0ea90a6a9aedf0a2269cda3b415eaa4b3f79522bc3d0ed209e = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[35] ^ 
        y_nr_in[55] ^ 
        y_nr_in[93] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[53] = 
I15397ad3270aed0ea90a6a9aedf0a2269cda3b415eaa4b3f79522bc3d0ed209e ^ 
0; 



wire Ia8e65506773efb18623b15c871910b9e506278ad08cdc3d9af85584eb585196d; 
assign Ia8e65506773efb18623b15c871910b9e506278ad08cdc3d9af85584eb585196d = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[32] ^ 
        y_nr_in[52] ^ 
        y_nr_in[94] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[54] = 
Ia8e65506773efb18623b15c871910b9e506278ad08cdc3d9af85584eb585196d ^ 
0; 



wire I9268d3a7b0e4e454dcfb018b47fa0cbb261e1de20c3fc00578cf4338a116de9d; 
assign I9268d3a7b0e4e454dcfb018b47fa0cbb261e1de20c3fc00578cf4338a116de9d = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[33] ^ 
        y_nr_in[53] ^ 
        y_nr_in[95] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[55] = 
I9268d3a7b0e4e454dcfb018b47fa0cbb261e1de20c3fc00578cf4338a116de9d ^ 
0; 



wire Ic948b765801b28252db81a845202ed5bb4c7b88d185735c290b087faf31e54f3; 
assign Ic948b765801b28252db81a845202ed5bb4c7b88d185735c290b087faf31e54f3 = 
        y_nr_in[7] ^ 
        y_nr_in[25] ^ 
        y_nr_in[47] ^ 
        y_nr_in[52] ^ 
        y_nr_in[96] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[56] = 
Ic948b765801b28252db81a845202ed5bb4c7b88d185735c290b087faf31e54f3 ^ 
0; 



wire Ie7fba38c244b4b0063545d270e36e5c6de425f13ee76efbea7f998b1806575d8; 
assign Ie7fba38c244b4b0063545d270e36e5c6de425f13ee76efbea7f998b1806575d8 = 
        y_nr_in[4] ^ 
        y_nr_in[26] ^ 
        y_nr_in[44] ^ 
        y_nr_in[53] ^ 
        y_nr_in[97] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[57] = 
Ie7fba38c244b4b0063545d270e36e5c6de425f13ee76efbea7f998b1806575d8 ^ 
0; 



wire Ic78a37f6dff689a73e3c867b6a1f732d8b87e77e148590359b6808c8f63ba162; 
assign Ic78a37f6dff689a73e3c867b6a1f732d8b87e77e148590359b6808c8f63ba162 = 
        y_nr_in[5] ^ 
        y_nr_in[27] ^ 
        y_nr_in[45] ^ 
        y_nr_in[54] ^ 
        y_nr_in[98] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[58] = 
Ic78a37f6dff689a73e3c867b6a1f732d8b87e77e148590359b6808c8f63ba162 ^ 
0; 



wire I6b93a394f20c2016695ccb4f7b85a006dc392fa36957b0a32a681c889a3d7b9f; 
assign I6b93a394f20c2016695ccb4f7b85a006dc392fa36957b0a32a681c889a3d7b9f = 
        y_nr_in[6] ^ 
        y_nr_in[24] ^ 
        y_nr_in[46] ^ 
        y_nr_in[55] ^ 
        y_nr_in[99] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[59] = 
I6b93a394f20c2016695ccb4f7b85a006dc392fa36957b0a32a681c889a3d7b9f ^ 
0; 



wire I007726f15ab00032d1871542c0e2231f004a3dbf62ec3feeeeb5173645e9c865; 
assign I007726f15ab00032d1871542c0e2231f004a3dbf62ec3feeeeb5173645e9c865 = 
        y_nr_in[3] ^ 
        y_nr_in[43] ^ 
        y_nr_in[45] ^ 
        y_nr_in[100] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[60] = 
I007726f15ab00032d1871542c0e2231f004a3dbf62ec3feeeeb5173645e9c865 ^ 
0; 



wire I10b3e9eaae0279c310f37ccd71904c84928328ed0e0295c3570662e302fa970a; 
assign I10b3e9eaae0279c310f37ccd71904c84928328ed0e0295c3570662e302fa970a = 
        y_nr_in[0] ^ 
        y_nr_in[40] ^ 
        y_nr_in[46] ^ 
        y_nr_in[101] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[61] = 
I10b3e9eaae0279c310f37ccd71904c84928328ed0e0295c3570662e302fa970a ^ 
0; 



wire I87613384bb8a7868c938a170f77b161f54493631a78fe81a7a7b04acc9e32b78; 
assign I87613384bb8a7868c938a170f77b161f54493631a78fe81a7a7b04acc9e32b78 = 
        y_nr_in[1] ^ 
        y_nr_in[41] ^ 
        y_nr_in[47] ^ 
        y_nr_in[102] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[62] = 
I87613384bb8a7868c938a170f77b161f54493631a78fe81a7a7b04acc9e32b78 ^ 
0; 



wire I894dd1817650b7f2bd2193783393fa9c2261579e5002d007926d5fbc0b910046; 
assign I894dd1817650b7f2bd2193783393fa9c2261579e5002d007926d5fbc0b910046 = 
        y_nr_in[2] ^ 
        y_nr_in[42] ^ 
        y_nr_in[44] ^ 
        y_nr_in[103] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[63] = 
I894dd1817650b7f2bd2193783393fa9c2261579e5002d007926d5fbc0b910046 ^ 
0; 



wire I65a0c6df5ad822e458be8380dd3471ff79fcab89a4f67fc5660d895af1733783; 
assign I65a0c6df5ad822e458be8380dd3471ff79fcab89a4f67fc5660d895af1733783 = 
        y_nr_in[7] ^ 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
        y_nr_in[50] ^ 
        y_nr_in[104] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[64] = 
I65a0c6df5ad822e458be8380dd3471ff79fcab89a4f67fc5660d895af1733783 ^ 
0; 



wire Icff0e6943b82a3293ff9dec141aacf6ee3e21c67458206a952738748c8e39ef1; 
assign Icff0e6943b82a3293ff9dec141aacf6ee3e21c67458206a952738748c8e39ef1 = 
        y_nr_in[4] ^ 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
        y_nr_in[51] ^ 
        y_nr_in[105] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[65] = 
Icff0e6943b82a3293ff9dec141aacf6ee3e21c67458206a952738748c8e39ef1 ^ 
0; 



wire I896c0703d30b5b2c87bc9c0d3ef81aeb24ed2bd11a232c442aba62d61b26172d; 
assign I896c0703d30b5b2c87bc9c0d3ef81aeb24ed2bd11a232c442aba62d61b26172d = 
        y_nr_in[5] ^ 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
        y_nr_in[48] ^ 
        y_nr_in[106] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[66] = 
I896c0703d30b5b2c87bc9c0d3ef81aeb24ed2bd11a232c442aba62d61b26172d ^ 
0; 



wire I81949e45ff6df2d131be75edd099ce3ec8942af4b5a1edc98fe909f342a92f37; 
assign I81949e45ff6df2d131be75edd099ce3ec8942af4b5a1edc98fe909f342a92f37 = 
        y_nr_in[6] ^ 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
        y_nr_in[49] ^ 
        y_nr_in[107] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[67] = 
I81949e45ff6df2d131be75edd099ce3ec8942af4b5a1edc98fe909f342a92f37 ^ 
0; 



wire If9ba3bf083697edc1ad40c606f53666a4ffdc23f68e26f82e6d283cea2fb4e01; 
assign If9ba3bf083697edc1ad40c606f53666a4ffdc23f68e26f82e6d283cea2fb4e01 = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[46] ^ 
        y_nr_in[48] ^ 
        y_nr_in[108] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[68] = 
If9ba3bf083697edc1ad40c606f53666a4ffdc23f68e26f82e6d283cea2fb4e01 ^ 
0; 



wire I1e63b71c64c10c264bf211563596fbc4ea9077598c159461bcb60cdc8e3b0ee4; 
assign I1e63b71c64c10c264bf211563596fbc4ea9077598c159461bcb60cdc8e3b0ee4 = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[47] ^ 
        y_nr_in[49] ^ 
        y_nr_in[109] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[69] = 
I1e63b71c64c10c264bf211563596fbc4ea9077598c159461bcb60cdc8e3b0ee4 ^ 
0; 



wire I23506b6c3d31e69452a3dcd4cbc892909c621f67a05c17901116f07116e77ab6; 
assign I23506b6c3d31e69452a3dcd4cbc892909c621f67a05c17901116f07116e77ab6 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[44] ^ 
        y_nr_in[50] ^ 
        y_nr_in[110] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[70] = 
I23506b6c3d31e69452a3dcd4cbc892909c621f67a05c17901116f07116e77ab6 ^ 
0; 



wire Iba05f3c0c354ff1968ab792f9724617bd9e01c802df4fc7c143df3b11e865a1b; 
assign Iba05f3c0c354ff1968ab792f9724617bd9e01c802df4fc7c143df3b11e865a1b = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[45] ^ 
        y_nr_in[51] ^ 
        y_nr_in[111] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[71] = 
Iba05f3c0c354ff1968ab792f9724617bd9e01c802df4fc7c143df3b11e865a1b ^ 
0; 



wire I226987acce4f66cc93d4f1f184b1081306f28001528a0db24d5a57bb4aeb28b6; 
assign I226987acce4f66cc93d4f1f184b1081306f28001528a0db24d5a57bb4aeb28b6 = 
        y_nr_in[0] ^ 
        y_nr_in[26] ^ 
        y_nr_in[30] ^ 
        y_nr_in[112] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[72] = 
I226987acce4f66cc93d4f1f184b1081306f28001528a0db24d5a57bb4aeb28b6 ^ 
0; 



wire Ib441bd8d21dc9f52b7e6b034aaa811ee40802e92c5241db91eebf50ae50a58dc; 
assign Ib441bd8d21dc9f52b7e6b034aaa811ee40802e92c5241db91eebf50ae50a58dc = 
        y_nr_in[1] ^ 
        y_nr_in[27] ^ 
        y_nr_in[31] ^ 
        y_nr_in[113] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[73] = 
Ib441bd8d21dc9f52b7e6b034aaa811ee40802e92c5241db91eebf50ae50a58dc ^ 
0; 



wire I97bb7b93e1c49d40c0ed8c3f09a0120028b65877d30e418e99ddb7140a6f7f43; 
assign I97bb7b93e1c49d40c0ed8c3f09a0120028b65877d30e418e99ddb7140a6f7f43 = 
        y_nr_in[2] ^ 
        y_nr_in[24] ^ 
        y_nr_in[28] ^ 
        y_nr_in[114] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[74] = 
I97bb7b93e1c49d40c0ed8c3f09a0120028b65877d30e418e99ddb7140a6f7f43 ^ 
0; 



wire I1c870b52db1059eb26e38f2e16bff0743a5d35b2771339689e244c0f31fe2abe; 
assign I1c870b52db1059eb26e38f2e16bff0743a5d35b2771339689e244c0f31fe2abe = 
        y_nr_in[3] ^ 
        y_nr_in[25] ^ 
        y_nr_in[29] ^ 
        y_nr_in[115] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[75] = 
I1c870b52db1059eb26e38f2e16bff0743a5d35b2771339689e244c0f31fe2abe ^ 
0; 



wire Ie6bb8d210bacc308c2f64785de6697a550b4d5158fb4b2d1903a4b1cfda09f82; 
assign Ie6bb8d210bacc308c2f64785de6697a550b4d5158fb4b2d1903a4b1cfda09f82 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[41] ^ 
        y_nr_in[116] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[76] = 
Ie6bb8d210bacc308c2f64785de6697a550b4d5158fb4b2d1903a4b1cfda09f82 ^ 
0; 



wire I0aabeae0f04a070f5c5a0630dd54ad72ab6b729cf47554d3228bbb154ae64deb; 
assign I0aabeae0f04a070f5c5a0630dd54ad72ab6b729cf47554d3228bbb154ae64deb = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[42] ^ 
        y_nr_in[117] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[77] = 
I0aabeae0f04a070f5c5a0630dd54ad72ab6b729cf47554d3228bbb154ae64deb ^ 
0; 



wire Ie0011cc23ee1152177360e4f99d5b7f5544a8e376aeca83eefb6d7a768e187a7; 
assign Ie0011cc23ee1152177360e4f99d5b7f5544a8e376aeca83eefb6d7a768e187a7 = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[43] ^ 
        y_nr_in[118] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[78] = 
Ie0011cc23ee1152177360e4f99d5b7f5544a8e376aeca83eefb6d7a768e187a7 ^ 
0; 



wire Id3f138b278c9fb85d20ad3e79ae7571bdd214a2a4739d72916ea106442b280ab; 
assign Id3f138b278c9fb85d20ad3e79ae7571bdd214a2a4739d72916ea106442b280ab = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[40] ^ 
        y_nr_in[119] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[79] = 
Id3f138b278c9fb85d20ad3e79ae7571bdd214a2a4739d72916ea106442b280ab ^ 
0; 



wire I817d2bad756252a5d8a6a15f128d70d9a21980c4709b4c17542219c339120a40; 
assign I817d2bad756252a5d8a6a15f128d70d9a21980c4709b4c17542219c339120a40 = 
        y_nr_in[6] ^ 
        y_nr_in[17] ^ 
        y_nr_in[45] ^ 
        y_nr_in[120] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[80] = 
I817d2bad756252a5d8a6a15f128d70d9a21980c4709b4c17542219c339120a40 ^ 
0; 



wire Ia4c380315cff761b2fdd6dc9aa4fff5462d27d3037dce146a45875a7a5bb4df8; 
assign Ia4c380315cff761b2fdd6dc9aa4fff5462d27d3037dce146a45875a7a5bb4df8 = 
        y_nr_in[7] ^ 
        y_nr_in[18] ^ 
        y_nr_in[46] ^ 
        y_nr_in[121] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[81] = 
Ia4c380315cff761b2fdd6dc9aa4fff5462d27d3037dce146a45875a7a5bb4df8 ^ 
0; 



wire If271fdce69f8cacb9e600fc90b61ab1511716fcb86913ba38f665cacabb50fe8; 
assign If271fdce69f8cacb9e600fc90b61ab1511716fcb86913ba38f665cacabb50fe8 = 
        y_nr_in[4] ^ 
        y_nr_in[19] ^ 
        y_nr_in[47] ^ 
        y_nr_in[122] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[82] = 
If271fdce69f8cacb9e600fc90b61ab1511716fcb86913ba38f665cacabb50fe8 ^ 
0; 



wire Iaac030fe8d7fe878e27fbda3fb868dcfa515c6e7513dc98d3a8d0bbe6d57675e; 
assign Iaac030fe8d7fe878e27fbda3fb868dcfa515c6e7513dc98d3a8d0bbe6d57675e = 
        y_nr_in[5] ^ 
        y_nr_in[16] ^ 
        y_nr_in[44] ^ 
        y_nr_in[123] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[83] = 
Iaac030fe8d7fe878e27fbda3fb868dcfa515c6e7513dc98d3a8d0bbe6d57675e ^ 
0; 



wire Ia96fb479d1d6c02b5c3e481de6867e9d0513243d2170cb49c08d90fb41839250; 
assign Ia96fb479d1d6c02b5c3e481de6867e9d0513243d2170cb49c08d90fb41839250 = 
        y_nr_in[0] ^ 
        y_nr_in[34] ^ 
        y_nr_in[54] ^ 
        y_nr_in[124] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[84] = 
Ia96fb479d1d6c02b5c3e481de6867e9d0513243d2170cb49c08d90fb41839250 ^ 
0; 



wire I88f12ff1bcc190c53bb7c2b6c96dbe7afbd7c7e25b870e14082445f1c8cc5d2b; 
assign I88f12ff1bcc190c53bb7c2b6c96dbe7afbd7c7e25b870e14082445f1c8cc5d2b = 
        y_nr_in[1] ^ 
        y_nr_in[35] ^ 
        y_nr_in[55] ^ 
        y_nr_in[125] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[85] = 
I88f12ff1bcc190c53bb7c2b6c96dbe7afbd7c7e25b870e14082445f1c8cc5d2b ^ 
0; 



wire Ia51c100452ac1527679780a2666be18950106bb42c6022fe02e67de531fb38bd; 
assign Ia51c100452ac1527679780a2666be18950106bb42c6022fe02e67de531fb38bd = 
        y_nr_in[2] ^ 
        y_nr_in[32] ^ 
        y_nr_in[52] ^ 
        y_nr_in[126] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[86] = 
Ia51c100452ac1527679780a2666be18950106bb42c6022fe02e67de531fb38bd ^ 
0; 



wire I6d52676190fa65365e3cddf27f40aa2d08ce8920bf4163237fb93a1909697597; 
assign I6d52676190fa65365e3cddf27f40aa2d08ce8920bf4163237fb93a1909697597 = 
        y_nr_in[3] ^ 
        y_nr_in[33] ^ 
        y_nr_in[53] ^ 
        y_nr_in[127] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[87] = 
I6d52676190fa65365e3cddf27f40aa2d08ce8920bf4163237fb93a1909697597 ^ 
0; 



wire I6bd5e8ab0c792d1d26fd6a07d8654383129caf127128980988d5425b66dea09f; 
assign I6bd5e8ab0c792d1d26fd6a07d8654383129caf127128980988d5425b66dea09f = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
        y_nr_in[128] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[88] = 
I6bd5e8ab0c792d1d26fd6a07d8654383129caf127128980988d5425b66dea09f ^ 
0; 



wire I835d5175e5bf4d6fe594d11a7e468458124ad49d7ece381e64eea258d0334700; 
assign I835d5175e5bf4d6fe594d11a7e468458124ad49d7ece381e64eea258d0334700 = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
        y_nr_in[129] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[89] = 
I835d5175e5bf4d6fe594d11a7e468458124ad49d7ece381e64eea258d0334700 ^ 
0; 



wire I27acd5f33c9d37311573644c4981723ce95a321acf13c6129616189d024cc6cf; 
assign I27acd5f33c9d37311573644c4981723ce95a321acf13c6129616189d024cc6cf = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
        y_nr_in[130] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[90] = 
I27acd5f33c9d37311573644c4981723ce95a321acf13c6129616189d024cc6cf ^ 
0; 



wire I11e423c1cee3dfc6efb69311d7010c2c96b708fdf40870e28d5b0845404d9e4f; 
assign I11e423c1cee3dfc6efb69311d7010c2c96b708fdf40870e28d5b0845404d9e4f = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
        y_nr_in[131] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[91] = 
I11e423c1cee3dfc6efb69311d7010c2c96b708fdf40870e28d5b0845404d9e4f ^ 
0; 



wire I3d2e1897d88ee4b73834010cfa6b8cd7dbd688988e9ac4df1335d9d37069a945; 
assign I3d2e1897d88ee4b73834010cfa6b8cd7dbd688988e9ac4df1335d9d37069a945 = 
        y_nr_in[3] ^ 
        y_nr_in[15] ^ 
        y_nr_in[22] ^ 
        y_nr_in[132] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[92] = 
I3d2e1897d88ee4b73834010cfa6b8cd7dbd688988e9ac4df1335d9d37069a945 ^ 
0; 



wire Iac36bda63af4630e9a6c0c775807c887b2a5ca0dd73b74e44add776990f98d95; 
assign Iac36bda63af4630e9a6c0c775807c887b2a5ca0dd73b74e44add776990f98d95 = 
        y_nr_in[0] ^ 
        y_nr_in[12] ^ 
        y_nr_in[23] ^ 
        y_nr_in[133] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[93] = 
Iac36bda63af4630e9a6c0c775807c887b2a5ca0dd73b74e44add776990f98d95 ^ 
0; 



wire I62caa4186011831a856349b528e7960392ea47b5251d440b34cb851a3d1dc110; 
assign I62caa4186011831a856349b528e7960392ea47b5251d440b34cb851a3d1dc110 = 
        y_nr_in[1] ^ 
        y_nr_in[13] ^ 
        y_nr_in[20] ^ 
        y_nr_in[134] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[94] = 
I62caa4186011831a856349b528e7960392ea47b5251d440b34cb851a3d1dc110 ^ 
0; 



wire Icb2398e1bedbaec03b084b301cafc1a27801836e82376f7b60f52844aecfbb8c; 
assign Icb2398e1bedbaec03b084b301cafc1a27801836e82376f7b60f52844aecfbb8c = 
        y_nr_in[2] ^ 
        y_nr_in[14] ^ 
        y_nr_in[21] ^ 
        y_nr_in[135] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[95] = 
Icb2398e1bedbaec03b084b301cafc1a27801836e82376f7b60f52844aecfbb8c ^ 
0; 



wire If8eadc7cfcc71a24af45cc9d48724d2abf589bd1318ff67a395bf55783660f0c; 
assign If8eadc7cfcc71a24af45cc9d48724d2abf589bd1318ff67a395bf55783660f0c = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
        y_nr_in[36] ^ 
        y_nr_in[136] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[96] = 
If8eadc7cfcc71a24af45cc9d48724d2abf589bd1318ff67a395bf55783660f0c ^ 
0; 



wire I2d0933613217d268e25a1aac304f4aee5638748fef3951272c2b91efecd93bdb; 
assign I2d0933613217d268e25a1aac304f4aee5638748fef3951272c2b91efecd93bdb = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
        y_nr_in[37] ^ 
        y_nr_in[137] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[97] = 
I2d0933613217d268e25a1aac304f4aee5638748fef3951272c2b91efecd93bdb ^ 
0; 



wire I41629d3151ecea09c2d44e6fc04f48f4a4f18fffd7c4810de0f4b7fa4f53dfd4; 
assign I41629d3151ecea09c2d44e6fc04f48f4a4f18fffd7c4810de0f4b7fa4f53dfd4 = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
        y_nr_in[38] ^ 
        y_nr_in[138] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[98] = 
I41629d3151ecea09c2d44e6fc04f48f4a4f18fffd7c4810de0f4b7fa4f53dfd4 ^ 
0; 



wire Id30b3770b2e8a6c5e42a801d5c6713fff3ae0c9d2390c2bffec9ee45be1e87ba; 
assign Id30b3770b2e8a6c5e42a801d5c6713fff3ae0c9d2390c2bffec9ee45be1e87ba = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
        y_nr_in[39] ^ 
        y_nr_in[139] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[99] = 
Id30b3770b2e8a6c5e42a801d5c6713fff3ae0c9d2390c2bffec9ee45be1e87ba ^ 
0; 



wire I635529633fb5c781ff2eb732acb4eee465bb9e4b6d4183f39b4865ba4eb31b4b; 
assign I635529633fb5c781ff2eb732acb4eee465bb9e4b6d4183f39b4865ba4eb31b4b = 
        y_nr_in[0] ^ 
        y_nr_in[20] ^ 
        y_nr_in[140] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[100] = 
I635529633fb5c781ff2eb732acb4eee465bb9e4b6d4183f39b4865ba4eb31b4b ^ 
0; 



wire Ib43f498373d2604355dda197f261dc55aced0df6271d3a9deccb273e9b367ded; 
assign Ib43f498373d2604355dda197f261dc55aced0df6271d3a9deccb273e9b367ded = 
        y_nr_in[1] ^ 
        y_nr_in[21] ^ 
        y_nr_in[141] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[101] = 
Ib43f498373d2604355dda197f261dc55aced0df6271d3a9deccb273e9b367ded ^ 
0; 



wire I4be9db8469c22ef12ff4969ebf88b2a0a3e325555b340a91c0f2ecfcac19aa65; 
assign I4be9db8469c22ef12ff4969ebf88b2a0a3e325555b340a91c0f2ecfcac19aa65 = 
        y_nr_in[2] ^ 
        y_nr_in[22] ^ 
        y_nr_in[142] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[102] = 
I4be9db8469c22ef12ff4969ebf88b2a0a3e325555b340a91c0f2ecfcac19aa65 ^ 
0; 



wire Ia6e8d5c54e6e3484c792ea4fb20d5fcee3237194f07ec815e34d99a3e9cfd93b; 
assign Ia6e8d5c54e6e3484c792ea4fb20d5fcee3237194f07ec815e34d99a3e9cfd93b = 
        y_nr_in[3] ^ 
        y_nr_in[23] ^ 
        y_nr_in[143] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[103] = 
Ia6e8d5c54e6e3484c792ea4fb20d5fcee3237194f07ec815e34d99a3e9cfd93b ^ 
0; 



wire I9d1526550d0b0bfc7e7e25788aa16598e9cbeaaf8102db6f6df1374d4c8a3e20; 
assign I9d1526550d0b0bfc7e7e25788aa16598e9cbeaaf8102db6f6df1374d4c8a3e20 = 
        y_nr_in[9] ^ 
        y_nr_in[31] ^ 
        y_nr_in[48] ^ 
        y_nr_in[54] ^ 
        y_nr_in[144] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[104] = 
I9d1526550d0b0bfc7e7e25788aa16598e9cbeaaf8102db6f6df1374d4c8a3e20 ^ 
0; 



wire Icf0fa899a5eaa151abe226aa3c4898a14f6ccfb446cc37c6938972da56c7b6be; 
assign Icf0fa899a5eaa151abe226aa3c4898a14f6ccfb446cc37c6938972da56c7b6be = 
        y_nr_in[10] ^ 
        y_nr_in[28] ^ 
        y_nr_in[49] ^ 
        y_nr_in[55] ^ 
        y_nr_in[145] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[105] = 
Icf0fa899a5eaa151abe226aa3c4898a14f6ccfb446cc37c6938972da56c7b6be ^ 
0; 



wire I8ff28927e344f2a273e2babaab16ab8f79e26d11708a05f6afdba223b716fe36; 
assign I8ff28927e344f2a273e2babaab16ab8f79e26d11708a05f6afdba223b716fe36 = 
        y_nr_in[11] ^ 
        y_nr_in[29] ^ 
        y_nr_in[50] ^ 
        y_nr_in[52] ^ 
        y_nr_in[146] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[106] = 
I8ff28927e344f2a273e2babaab16ab8f79e26d11708a05f6afdba223b716fe36 ^ 
0; 



wire I829f2f6aa47f6700a660b0d559837b3a5d7d208f0a86238bea5ac0ccc900e446; 
assign I829f2f6aa47f6700a660b0d559837b3a5d7d208f0a86238bea5ac0ccc900e446 = 
        y_nr_in[8] ^ 
        y_nr_in[30] ^ 
        y_nr_in[51] ^ 
        y_nr_in[53] ^ 
        y_nr_in[147] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[107] = 
I829f2f6aa47f6700a660b0d559837b3a5d7d208f0a86238bea5ac0ccc900e446 ^ 
0; 



wire Ibc34c5299448c47acb4b03b7250f319573b1c05abbb8c2b3458cb0a34facbaf9; 
assign Ibc34c5299448c47acb4b03b7250f319573b1c05abbb8c2b3458cb0a34facbaf9 = 
        y_nr_in[0] ^ 
        y_nr_in[27] ^ 
        y_nr_in[148] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[108] = 
Ibc34c5299448c47acb4b03b7250f319573b1c05abbb8c2b3458cb0a34facbaf9 ^ 
0; 



wire I53c2782b0c8ab82eaf6d3c901b1a704d8face020eff60bab85ac16d20cacfc89; 
assign I53c2782b0c8ab82eaf6d3c901b1a704d8face020eff60bab85ac16d20cacfc89 = 
        y_nr_in[1] ^ 
        y_nr_in[24] ^ 
        y_nr_in[149] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[109] = 
I53c2782b0c8ab82eaf6d3c901b1a704d8face020eff60bab85ac16d20cacfc89 ^ 
0; 



wire I012dd64060af6bba3f9980b2a8bba98e058138b704cabfe32080d48ef5a699c0; 
assign I012dd64060af6bba3f9980b2a8bba98e058138b704cabfe32080d48ef5a699c0 = 
        y_nr_in[2] ^ 
        y_nr_in[25] ^ 
        y_nr_in[150] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[110] = 
I012dd64060af6bba3f9980b2a8bba98e058138b704cabfe32080d48ef5a699c0 ^ 
0; 



wire I09f86a8aee66c743be462b26e4bf264d1b5e7d9371d02f27ec876c1c023b410c; 
assign I09f86a8aee66c743be462b26e4bf264d1b5e7d9371d02f27ec876c1c023b410c = 
        y_nr_in[3] ^ 
        y_nr_in[26] ^ 
        y_nr_in[151] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[111] = 
I09f86a8aee66c743be462b26e4bf264d1b5e7d9371d02f27ec876c1c023b410c ^ 
0; 



wire I183c80ed9f4376e550fe169249a2e349d8e1c99c457ba08be8025586e75a0e23; 
assign I183c80ed9f4376e550fe169249a2e349d8e1c99c457ba08be8025586e75a0e23 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[23] ^ 
        y_nr_in[152] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[112] = 
I183c80ed9f4376e550fe169249a2e349d8e1c99c457ba08be8025586e75a0e23 ^ 
0; 



wire Ibe5ca11f38b74b767d5092156093fa3e335a2af04e5b1a74ac6b7dea73f21c93; 
assign Ibe5ca11f38b74b767d5092156093fa3e335a2af04e5b1a74ac6b7dea73f21c93 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[20] ^ 
        y_nr_in[153] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[113] = 
Ibe5ca11f38b74b767d5092156093fa3e335a2af04e5b1a74ac6b7dea73f21c93 ^ 
0; 



wire I586fb4b534c740086576f7412ab9956c8b7aecef364c087673f5f61e77f82a1a; 
assign I586fb4b534c740086576f7412ab9956c8b7aecef364c087673f5f61e77f82a1a = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[21] ^ 
        y_nr_in[154] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[114] = 
I586fb4b534c740086576f7412ab9956c8b7aecef364c087673f5f61e77f82a1a ^ 
0; 



wire I7561f10d84b41620a8ef4f2d92d36edb02cd2281977f91a2291be0d65ccfb4ea; 
assign I7561f10d84b41620a8ef4f2d92d36edb02cd2281977f91a2291be0d65ccfb4ea = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[22] ^ 
        y_nr_in[155] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[115] = 
I7561f10d84b41620a8ef4f2d92d36edb02cd2281977f91a2291be0d65ccfb4ea ^ 
0; 



wire Iba7e7ff6d4d2eceb97e52d11e1af99bc8711b2358bc90f941b1d5b7054d8f022; 
assign Iba7e7ff6d4d2eceb97e52d11e1af99bc8711b2358bc90f941b1d5b7054d8f022 = 
        y_nr_in[2] ^ 
        y_nr_in[16] ^ 
        y_nr_in[156] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[116] = 
Iba7e7ff6d4d2eceb97e52d11e1af99bc8711b2358bc90f941b1d5b7054d8f022 ^ 
0; 



wire I548677fe1e30d06ab0c5e3791db2e34537fbf6b1f484265913c3f2bf1fbc1b1d; 
assign I548677fe1e30d06ab0c5e3791db2e34537fbf6b1f484265913c3f2bf1fbc1b1d = 
        y_nr_in[3] ^ 
        y_nr_in[17] ^ 
        y_nr_in[157] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[117] = 
I548677fe1e30d06ab0c5e3791db2e34537fbf6b1f484265913c3f2bf1fbc1b1d ^ 
0; 



wire I740598afb66f316809fb1627c7594236da13cf4bf6fe3034b45247a0bad3d868; 
assign I740598afb66f316809fb1627c7594236da13cf4bf6fe3034b45247a0bad3d868 = 
        y_nr_in[0] ^ 
        y_nr_in[18] ^ 
        y_nr_in[158] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[118] = 
I740598afb66f316809fb1627c7594236da13cf4bf6fe3034b45247a0bad3d868 ^ 
0; 



wire I8866602383e779b8e52b8889527675ab62a90b2a636768b5ec48321720412ad5; 
assign I8866602383e779b8e52b8889527675ab62a90b2a636768b5ec48321720412ad5 = 
        y_nr_in[1] ^ 
        y_nr_in[19] ^ 
        y_nr_in[159] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[119] = 
I8866602383e779b8e52b8889527675ab62a90b2a636768b5ec48321720412ad5 ^ 
0; 



wire I1e88a0a859a6e0f4a59680a9fc99c809f5f6ccffbd5f2cd0aa90ba328f643dc5; 
assign I1e88a0a859a6e0f4a59680a9fc99c809f5f6ccffbd5f2cd0aa90ba328f643dc5 = 
        y_nr_in[11] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[36] ^ 
        y_nr_in[160] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[120] = 
I1e88a0a859a6e0f4a59680a9fc99c809f5f6ccffbd5f2cd0aa90ba328f643dc5 ^ 
0; 



wire I548f4fbc1ec7695988dab22516f9c93ea264c7834ff89f5f52c11a551b874743; 
assign I548f4fbc1ec7695988dab22516f9c93ea264c7834ff89f5f52c11a551b874743 = 
        y_nr_in[8] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[37] ^ 
        y_nr_in[161] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[121] = 
I548f4fbc1ec7695988dab22516f9c93ea264c7834ff89f5f52c11a551b874743 ^ 
0; 



wire I124bf7f050a4d1f64408c9f7a1a111d04d6d59047d613ee06daaeb9d0614b57b; 
assign I124bf7f050a4d1f64408c9f7a1a111d04d6d59047d613ee06daaeb9d0614b57b = 
        y_nr_in[9] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[38] ^ 
        y_nr_in[162] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[122] = 
I124bf7f050a4d1f64408c9f7a1a111d04d6d59047d613ee06daaeb9d0614b57b ^ 
0; 



wire Ie460ea553c65465e294fbbe9f3021a8627d8243fc684ebeb2ba2e2bb77f577e0; 
assign Ie460ea553c65465e294fbbe9f3021a8627d8243fc684ebeb2ba2e2bb77f577e0 = 
        y_nr_in[10] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[39] ^ 
        y_nr_in[163] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[123] = 
Ie460ea553c65465e294fbbe9f3021a8627d8243fc684ebeb2ba2e2bb77f577e0 ^ 
0; 



wire I1a8e72beb7b2012de2b4e70c32e7c75928ab55c82aa3e4a54e81c3d15e070f27; 
assign I1a8e72beb7b2012de2b4e70c32e7c75928ab55c82aa3e4a54e81c3d15e070f27 = 
        y_nr_in[6] ^ 
        y_nr_in[53] ^ 
        y_nr_in[164] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[124] = 
I1a8e72beb7b2012de2b4e70c32e7c75928ab55c82aa3e4a54e81c3d15e070f27 ^ 
0; 



wire I9ec4d26cfe02337527e90e8741619742f322b87851a948babfa910f6e2e06d62; 
assign I9ec4d26cfe02337527e90e8741619742f322b87851a948babfa910f6e2e06d62 = 
        y_nr_in[7] ^ 
        y_nr_in[54] ^ 
        y_nr_in[165] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[125] = 
I9ec4d26cfe02337527e90e8741619742f322b87851a948babfa910f6e2e06d62 ^ 
0; 



wire I98f3cc475aa7cb3ef452e91ee8b36f0ad3a084ebaebdeee42f50ed322b765904; 
assign I98f3cc475aa7cb3ef452e91ee8b36f0ad3a084ebaebdeee42f50ed322b765904 = 
        y_nr_in[4] ^ 
        y_nr_in[55] ^ 
        y_nr_in[166] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[126] = 
I98f3cc475aa7cb3ef452e91ee8b36f0ad3a084ebaebdeee42f50ed322b765904 ^ 
0; 



wire Ic1da980412da922b348d1cf919be86a04e135bb552ab3f9a83888a600287ed9c; 
assign Ic1da980412da922b348d1cf919be86a04e135bb552ab3f9a83888a600287ed9c = 
        y_nr_in[5] ^ 
        y_nr_in[52] ^ 
        y_nr_in[167] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[127] = 
Ic1da980412da922b348d1cf919be86a04e135bb552ab3f9a83888a600287ed9c ^ 
0; 



wire Ief5434fcb978b538c56cd1e62bd39737afe99c3591661313922e534867485c3e; 
assign Ief5434fcb978b538c56cd1e62bd39737afe99c3591661313922e534867485c3e = 
        y_nr_in[2] ^ 
        y_nr_in[20] ^ 
        y_nr_in[50] ^ 
        y_nr_in[168] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[128] = 
Ief5434fcb978b538c56cd1e62bd39737afe99c3591661313922e534867485c3e ^ 
0; 



wire Ic923aca9c0e123e8526c516dfbaf9e12fe628ed7956a9245266d0c05e72ad072; 
assign Ic923aca9c0e123e8526c516dfbaf9e12fe628ed7956a9245266d0c05e72ad072 = 
        y_nr_in[3] ^ 
        y_nr_in[21] ^ 
        y_nr_in[51] ^ 
        y_nr_in[169] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[129] = 
Ic923aca9c0e123e8526c516dfbaf9e12fe628ed7956a9245266d0c05e72ad072 ^ 
0; 



wire Ied046dccaee2d2f5abceafb984589a6cbc250bf754e8c88cb4139eaa8e05a673; 
assign Ied046dccaee2d2f5abceafb984589a6cbc250bf754e8c88cb4139eaa8e05a673 = 
        y_nr_in[0] ^ 
        y_nr_in[22] ^ 
        y_nr_in[48] ^ 
        y_nr_in[170] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[130] = 
Ied046dccaee2d2f5abceafb984589a6cbc250bf754e8c88cb4139eaa8e05a673 ^ 
0; 



wire Id460401256d461c8446008f1a2a79aaadd0f52dc60b2409f50eb54f08a48165e; 
assign Id460401256d461c8446008f1a2a79aaadd0f52dc60b2409f50eb54f08a48165e = 
        y_nr_in[1] ^ 
        y_nr_in[23] ^ 
        y_nr_in[49] ^ 
        y_nr_in[171] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[131] = 
Id460401256d461c8446008f1a2a79aaadd0f52dc60b2409f50eb54f08a48165e ^ 
0; 



wire Id213bf07258b38900e6c46f518300c22d9fd5f18908a15092025c6cb84abfdd9; 
assign Id213bf07258b38900e6c46f518300c22d9fd5f18908a15092025c6cb84abfdd9 = 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
        y_nr_in[43] ^ 
        y_nr_in[172] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[132] = 
Id213bf07258b38900e6c46f518300c22d9fd5f18908a15092025c6cb84abfdd9 ^ 
0; 



wire I56684935e34c7f6d27c30daef8a0bef4f6bae679825dfaeaf7d9037915c85452; 
assign I56684935e34c7f6d27c30daef8a0bef4f6bae679825dfaeaf7d9037915c85452 = 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
        y_nr_in[40] ^ 
        y_nr_in[173] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[133] = 
I56684935e34c7f6d27c30daef8a0bef4f6bae679825dfaeaf7d9037915c85452 ^ 
0; 



wire I2c4d0b067fcb722018c8b55411adb913f75fe00b277ef1e0fd58d6903d8cdebf; 
assign I2c4d0b067fcb722018c8b55411adb913f75fe00b277ef1e0fd58d6903d8cdebf = 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
        y_nr_in[41] ^ 
        y_nr_in[174] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[134] = 
I2c4d0b067fcb722018c8b55411adb913f75fe00b277ef1e0fd58d6903d8cdebf ^ 
0; 



wire I25f169675f7b2c40d508a415966d827bc294d4c3895aa04d0a5100d473803c14; 
assign I25f169675f7b2c40d508a415966d827bc294d4c3895aa04d0a5100d473803c14 = 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
        y_nr_in[42] ^ 
        y_nr_in[175] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[135] = 
I25f169675f7b2c40d508a415966d827bc294d4c3895aa04d0a5100d473803c14 ^ 
0; 



wire I13e087bef67c2ce5927101c6c6e0090a15f05e93a0507d9014ea3401f480745e; 
assign I13e087bef67c2ce5927101c6c6e0090a15f05e93a0507d9014ea3401f480745e = 
        y_nr_in[3] ^ 
        y_nr_in[49] ^ 
        y_nr_in[52] ^ 
        y_nr_in[176] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[136] = 
I13e087bef67c2ce5927101c6c6e0090a15f05e93a0507d9014ea3401f480745e ^ 
0; 



wire Ifa999747365603ce92391d8e4d9394c0601d78531c3e1235d7141bdd1bb171ed; 
assign Ifa999747365603ce92391d8e4d9394c0601d78531c3e1235d7141bdd1bb171ed = 
        y_nr_in[0] ^ 
        y_nr_in[50] ^ 
        y_nr_in[53] ^ 
        y_nr_in[177] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[137] = 
Ifa999747365603ce92391d8e4d9394c0601d78531c3e1235d7141bdd1bb171ed ^ 
0; 



wire Idfec1ceb40ed0b911611f7f7e0c63c84f9109f367ab0af1988674965fbc3ca34; 
assign Idfec1ceb40ed0b911611f7f7e0c63c84f9109f367ab0af1988674965fbc3ca34 = 
        y_nr_in[1] ^ 
        y_nr_in[51] ^ 
        y_nr_in[54] ^ 
        y_nr_in[178] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[138] = 
Idfec1ceb40ed0b911611f7f7e0c63c84f9109f367ab0af1988674965fbc3ca34 ^ 
0; 



wire I2b19017cda532c473e23616c17d73afb77e4b0158e97e2f9ee9f9450e88c5108; 
assign I2b19017cda532c473e23616c17d73afb77e4b0158e97e2f9ee9f9450e88c5108 = 
        y_nr_in[2] ^ 
        y_nr_in[48] ^ 
        y_nr_in[55] ^ 
        y_nr_in[179] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[139] = 
I2b19017cda532c473e23616c17d73afb77e4b0158e97e2f9ee9f9450e88c5108 ^ 
0; 



wire I168e76ede86e369ea0fe70cc239c2ce829312bb2c81901b99e5b486f95332b2f; 
assign I168e76ede86e369ea0fe70cc239c2ce829312bb2c81901b99e5b486f95332b2f = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[47] ^ 
        y_nr_in[180] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[140] = 
I168e76ede86e369ea0fe70cc239c2ce829312bb2c81901b99e5b486f95332b2f ^ 
0; 



wire I8ab8ceb7257501f392c27a1cdcbd45cace80e3f4fc4285b9615c86b24856be35; 
assign I8ab8ceb7257501f392c27a1cdcbd45cace80e3f4fc4285b9615c86b24856be35 = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[44] ^ 
        y_nr_in[181] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[141] = 
I8ab8ceb7257501f392c27a1cdcbd45cace80e3f4fc4285b9615c86b24856be35 ^ 
0; 



wire I33292c0e118bd99d4c823ba2af97c7289c3776d62194b209a1421d1c14976d38; 
assign I33292c0e118bd99d4c823ba2af97c7289c3776d62194b209a1421d1c14976d38 = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[45] ^ 
        y_nr_in[182] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[142] = 
I33292c0e118bd99d4c823ba2af97c7289c3776d62194b209a1421d1c14976d38 ^ 
0; 



wire I34ba1272a20f37beb381565247934ca6e2e1de666d6a0feb586333de63380b59; 
assign I34ba1272a20f37beb381565247934ca6e2e1de666d6a0feb586333de63380b59 = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[46] ^ 
        y_nr_in[183] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[143] = 
I34ba1272a20f37beb381565247934ca6e2e1de666d6a0feb586333de63380b59 ^ 
0; 



wire I1e362f85d7d0b8b3bed640dcc5c7e1f1703141e53866ec0825ccff1ba18297f6; 
assign I1e362f85d7d0b8b3bed640dcc5c7e1f1703141e53866ec0825ccff1ba18297f6 = 
        y_nr_in[0] ^ 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
        y_nr_in[184] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[144] = 
I1e362f85d7d0b8b3bed640dcc5c7e1f1703141e53866ec0825ccff1ba18297f6 ^ 
0; 



wire I1c0c28df19037241029ddaaed1878c81c288207f4c296c5168e6378156b5f52c; 
assign I1c0c28df19037241029ddaaed1878c81c288207f4c296c5168e6378156b5f52c = 
        y_nr_in[1] ^ 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
        y_nr_in[185] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[145] = 
I1c0c28df19037241029ddaaed1878c81c288207f4c296c5168e6378156b5f52c ^ 
0; 



wire I589b23237566079f86870b64d1bb0cf663cb2e781e79e07115b9c9bdfbbcfb5f; 
assign I589b23237566079f86870b64d1bb0cf663cb2e781e79e07115b9c9bdfbbcfb5f = 
        y_nr_in[2] ^ 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
        y_nr_in[186] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[146] = 
I589b23237566079f86870b64d1bb0cf663cb2e781e79e07115b9c9bdfbbcfb5f ^ 
0; 



wire I59f36cddab524833c92b6f591130a898f93c2719d190e4ed77766788d65a84ab; 
assign I59f36cddab524833c92b6f591130a898f93c2719d190e4ed77766788d65a84ab = 
        y_nr_in[3] ^ 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
        y_nr_in[187] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[147] = 
I59f36cddab524833c92b6f591130a898f93c2719d190e4ed77766788d65a84ab ^ 
0; 



wire I068bbcde5f56c740277c9e5c7d69881d9bbf9f676864b0c31445340d7002f058; 
assign I068bbcde5f56c740277c9e5c7d69881d9bbf9f676864b0c31445340d7002f058 = 
        y_nr_in[43] ^ 
        y_nr_in[55] ^ 
        y_nr_in[188] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[148] = 
I068bbcde5f56c740277c9e5c7d69881d9bbf9f676864b0c31445340d7002f058 ^ 
0; 



wire I8be6e7b03ec56774494eb385f84ff747765133dedf7435da0720b8a4af27d09e; 
assign I8be6e7b03ec56774494eb385f84ff747765133dedf7435da0720b8a4af27d09e = 
        y_nr_in[40] ^ 
        y_nr_in[52] ^ 
        y_nr_in[189] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[149] = 
I8be6e7b03ec56774494eb385f84ff747765133dedf7435da0720b8a4af27d09e ^ 
0; 



wire Ibc32b9d6e7ce9601f2ed8dcd86dcbaf8a79f60859b8716968216007c0cee2443; 
assign Ibc32b9d6e7ce9601f2ed8dcd86dcbaf8a79f60859b8716968216007c0cee2443 = 
        y_nr_in[41] ^ 
        y_nr_in[53] ^ 
        y_nr_in[190] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[150] = 
Ibc32b9d6e7ce9601f2ed8dcd86dcbaf8a79f60859b8716968216007c0cee2443 ^ 
0; 



wire Idc954068278ec51e4f799a9374617c371b489938ccb49199457f36321c36258b; 
assign Idc954068278ec51e4f799a9374617c371b489938ccb49199457f36321c36258b = 
        y_nr_in[42] ^ 
        y_nr_in[54] ^ 
        y_nr_in[191] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[151] = 
Idc954068278ec51e4f799a9374617c371b489938ccb49199457f36321c36258b ^ 
0; 



wire I42a6e56d6b386e7e8141dc70e9e1a5ac7b6296794ad8e3c2d72a7d51a16efdca; 
assign I42a6e56d6b386e7e8141dc70e9e1a5ac7b6296794ad8e3c2d72a7d51a16efdca = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[46] ^ 
        y_nr_in[192] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[152] = 
I42a6e56d6b386e7e8141dc70e9e1a5ac7b6296794ad8e3c2d72a7d51a16efdca ^ 
0; 



wire I6465aad3fd136b121662710a7cbffb17792c48b3af2c14cd67ecc457c62310e4; 
assign I6465aad3fd136b121662710a7cbffb17792c48b3af2c14cd67ecc457c62310e4 = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[47] ^ 
        y_nr_in[193] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[153] = 
I6465aad3fd136b121662710a7cbffb17792c48b3af2c14cd67ecc457c62310e4 ^ 
0; 



wire I33e30920b3c5020dd3a6662ec05427a67059725e65f9668470eec1755a59f97e; 
assign I33e30920b3c5020dd3a6662ec05427a67059725e65f9668470eec1755a59f97e = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[44] ^ 
        y_nr_in[194] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[154] = 
I33e30920b3c5020dd3a6662ec05427a67059725e65f9668470eec1755a59f97e ^ 
0; 



wire I9d482d4edb12871b7fa8f4f251d84d19080ffa35272ae8d5d071a610b1972401; 
assign I9d482d4edb12871b7fa8f4f251d84d19080ffa35272ae8d5d071a610b1972401 = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[45] ^ 
        y_nr_in[195] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[155] = 
I9d482d4edb12871b7fa8f4f251d84d19080ffa35272ae8d5d071a610b1972401 ^ 
0; 



wire Ifda034d14f43980bfdec0086c9f215c2314c27b4b2e33ce828bb6f3553c9cdd9; 
assign Ifda034d14f43980bfdec0086c9f215c2314c27b4b2e33ce828bb6f3553c9cdd9 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[50] ^ 
        y_nr_in[196] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[156] = 
Ifda034d14f43980bfdec0086c9f215c2314c27b4b2e33ce828bb6f3553c9cdd9 ^ 
0; 



wire Id06a5ffbb0da9c3435179445b5cd9bd7b3276f5fec240e8e5ce9b0efa6d11cec; 
assign Id06a5ffbb0da9c3435179445b5cd9bd7b3276f5fec240e8e5ce9b0efa6d11cec = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[51] ^ 
        y_nr_in[197] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[157] = 
Id06a5ffbb0da9c3435179445b5cd9bd7b3276f5fec240e8e5ce9b0efa6d11cec ^ 
0; 



wire I04d7d839b0414897f0841839595d97d904afdd78b99e29be0a3e5f119851a8e5; 
assign I04d7d839b0414897f0841839595d97d904afdd78b99e29be0a3e5f119851a8e5 = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[48] ^ 
        y_nr_in[198] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[158] = 
I04d7d839b0414897f0841839595d97d904afdd78b99e29be0a3e5f119851a8e5 ^ 
0; 



wire I5daec9e5796bbd6fc33ca6b136cc0ebe23d741899c9dff1c7c42383012ced787; 
assign I5daec9e5796bbd6fc33ca6b136cc0ebe23d741899c9dff1c7c42383012ced787 = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[49] ^ 
        y_nr_in[199] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[159] = 
I5daec9e5796bbd6fc33ca6b136cc0ebe23d741899c9dff1c7c42383012ced787 ^ 
0; 



wire Id0771405707f40d21e97c9e476aebaaaa07e735d255a8b179fdaa8d7f11a716f; 
assign Id0771405707f40d21e97c9e476aebaaaa07e735d255a8b179fdaa8d7f11a716f = 
        y_nr_in[8] ^ 
        y_nr_in[43] ^ 
        y_nr_in[52] ^ 
        y_nr_in[200] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[160] = 
Id0771405707f40d21e97c9e476aebaaaa07e735d255a8b179fdaa8d7f11a716f ^ 
0; 



wire I7865c37819b58e5fda240d7f8992e42f295e4eca78b03a08f367fafe8c15fbbf; 
assign I7865c37819b58e5fda240d7f8992e42f295e4eca78b03a08f367fafe8c15fbbf = 
        y_nr_in[9] ^ 
        y_nr_in[40] ^ 
        y_nr_in[53] ^ 
        y_nr_in[201] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[161] = 
I7865c37819b58e5fda240d7f8992e42f295e4eca78b03a08f367fafe8c15fbbf ^ 
0; 



wire I96d0cd2ffcd997637e4aeac0e9598224187594760d9f54cf9e3a7a927792259c; 
assign I96d0cd2ffcd997637e4aeac0e9598224187594760d9f54cf9e3a7a927792259c = 
        y_nr_in[10] ^ 
        y_nr_in[41] ^ 
        y_nr_in[54] ^ 
        y_nr_in[202] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[162] = 
I96d0cd2ffcd997637e4aeac0e9598224187594760d9f54cf9e3a7a927792259c ^ 
0; 



wire Ic6a319304fd7fca920679069affbc8e184db6d362f387151a038db8b0ae57fe8; 
assign Ic6a319304fd7fca920679069affbc8e184db6d362f387151a038db8b0ae57fe8 = 
        y_nr_in[11] ^ 
        y_nr_in[42] ^ 
        y_nr_in[55] ^ 
        y_nr_in[203] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[163] = 
Ic6a319304fd7fca920679069affbc8e184db6d362f387151a038db8b0ae57fe8 ^ 
0; 



wire Ic315c229c5b58969dc552d7ac12986ca4bd140b2c2b6c3f1817a51f14b64ca4d; 
assign Ic315c229c5b58969dc552d7ac12986ca4bd140b2c2b6c3f1817a51f14b64ca4d = 
        y_nr_in[5] ^ 
        y_nr_in[21] ^ 
        y_nr_in[46] ^ 
        y_nr_in[204] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[164] = 
Ic315c229c5b58969dc552d7ac12986ca4bd140b2c2b6c3f1817a51f14b64ca4d ^ 
0; 



wire Idc653a6631b1430ba54f080f7c7d682bbf5ff462d871d1b8b8b2bc2e5ce2cb3a; 
assign Idc653a6631b1430ba54f080f7c7d682bbf5ff462d871d1b8b8b2bc2e5ce2cb3a = 
        y_nr_in[6] ^ 
        y_nr_in[22] ^ 
        y_nr_in[47] ^ 
        y_nr_in[205] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[165] = 
Idc653a6631b1430ba54f080f7c7d682bbf5ff462d871d1b8b8b2bc2e5ce2cb3a ^ 
0; 



wire I57fb4eebb0b52139d167f65b01752de6f072e9bfa51811a4e24a432640a4bac0; 
assign I57fb4eebb0b52139d167f65b01752de6f072e9bfa51811a4e24a432640a4bac0 = 
        y_nr_in[7] ^ 
        y_nr_in[23] ^ 
        y_nr_in[44] ^ 
        y_nr_in[206] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[166] = 
I57fb4eebb0b52139d167f65b01752de6f072e9bfa51811a4e24a432640a4bac0 ^ 
0; 



wire I3f556e466d879253b69c492c9b2b198cfd9c440cd598ceb8fa8284cde0ad3df0; 
assign I3f556e466d879253b69c492c9b2b198cfd9c440cd598ceb8fa8284cde0ad3df0 = 
        y_nr_in[4] ^ 
        y_nr_in[20] ^ 
        y_nr_in[45] ^ 
        y_nr_in[207] ^ 
0; 



assign I800f06299ed1c747ea99ba7e3d3514c2a6f018f998f100e828eff738a229aeb9[167] = 
I3f556e466d879253b69c492c9b2b198cfd9c440cd598ceb8fa8284cde0ad3df0 ^ 
0; 



