 reg  ['h1ffff:0] [$clog2('h7000+1)-1:0] I7ed8af01513aac613cc7f755746bce57 ;
