parameter n_minus_m = 'd40;
parameter n_int = 'd208;
parameter m_int = 'd168;



parameter z_int = 'd4;



wire [m_int-1:0] Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c; 
wire Ic03b2bba447638cf5ba15e511366289ff81c1b93d193a0538489ba2565296f0a;
assign Ic03b2bba447638cf5ba15e511366289ff81c1b93d193a0538489ba2565296f0a = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[14] ^ 
0; 



wire Iedd82dd94c389d4a476e5bb200b072f312af7202cbf32d65d7540e16bdf47035;
assign Iedd82dd94c389d4a476e5bb200b072f312af7202cbf32d65d7540e16bdf47035 = 
        y_nr_in[25] ^ 
        y_nr_in[37] ^ 
        y_nr_in[3] ^ 
0; 



wire Iacf9f0469ca978b08f5e278f94ee91a38d34cd1e73f172817c5442772535c61e;
assign Iacf9f0469ca978b08f5e278f94ee91a38d34cd1e73f172817c5442772535c61e = 
        y_nr_in[14] ^ 
        y_nr_in[17] ^ 
        y_nr_in[21] ^ 
0; 



wire I0992ec582a0556b79da864b679dbcf57f71ff5458bca91375e0829b6504d1032;
assign I0992ec582a0556b79da864b679dbcf57f71ff5458bca91375e0829b6504d1032 = 
        y_nr_in[26] ^ 
        y_nr_in[28] ^ 
        y_nr_in[32] ^ 
0; 



wire I47af3c7c5a7f4ab7b0fa73849e3eed0ad8251b62621cf07ed4b835d813ba1dbe;
assign I47af3c7c5a7f4ab7b0fa73849e3eed0ad8251b62621cf07ed4b835d813ba1dbe = 
        y_nr_in[36] ^ 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
0; 



wire Ib47a7459aef485060f49a417b8619cb078deb77bf7094c6a2b94a762211dcbdd;
assign Ib47a7459aef485060f49a417b8619cb078deb77bf7094c6a2b94a762211dcbdd = 
        y_nr_in[12] ^ 
        y_nr_in[16] ^ 
        y_nr_in[32] ^ 
0; 



wire Ia3174d0d2a2a5245e247f4d63e0bfb149961032d8797887d3b7c0611b8408fe8;
assign Ia3174d0d2a2a5245e247f4d63e0bfb149961032d8797887d3b7c0611b8408fe8 = 
        y_nr_in[4] ^ 
        y_nr_in[10] ^ 
        y_nr_in[18] ^ 
0; 



wire Ibddf4c3f19e99f47a435f4cf6dbd1ad1703e9534daf2edac08b153e0136279a4;
assign Ibddf4c3f19e99f47a435f4cf6dbd1ad1703e9534daf2edac08b153e0136279a4 = 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
        y_nr_in[30] ^ 
0; 



wire Ie62630445e48b8650666cb06a196cbe8fb464502c91319068e9b9c1c15bbf93e;
assign Ie62630445e48b8650666cb06a196cbe8fb464502c91319068e9b9c1c15bbf93e = 
        y_nr_in[34] ^ 
        y_nr_in[36] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[167] = 
Ic03b2bba447638cf5ba15e511366289ff81c1b93d193a0538489ba2565296f0a ^ 
Iedd82dd94c389d4a476e5bb200b072f312af7202cbf32d65d7540e16bdf47035 ^ 
Iacf9f0469ca978b08f5e278f94ee91a38d34cd1e73f172817c5442772535c61e ^ 
I0992ec582a0556b79da864b679dbcf57f71ff5458bca91375e0829b6504d1032 ^ 
I47af3c7c5a7f4ab7b0fa73849e3eed0ad8251b62621cf07ed4b835d813ba1dbe ^ 
Ib47a7459aef485060f49a417b8619cb078deb77bf7094c6a2b94a762211dcbdd ^ 
Ia3174d0d2a2a5245e247f4d63e0bfb149961032d8797887d3b7c0611b8408fe8 ^ 
Ibddf4c3f19e99f47a435f4cf6dbd1ad1703e9534daf2edac08b153e0136279a4 ^ 
Ie62630445e48b8650666cb06a196cbe8fb464502c91319068e9b9c1c15bbf93e ^ 
0; 



wire Iac791f5d19a7c542254f5d4b9b0fa6eef7eeb9b06f8a9916a3dc9da1bbda42ba;
assign Iac791f5d19a7c542254f5d4b9b0fa6eef7eeb9b06f8a9916a3dc9da1bbda42ba = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[15] ^ 
0; 



wire Ie88a242b25c2fbf1d9f5800d92b3fae86edf8b29993930dd06e7ecdcffacf212;
assign Ie88a242b25c2fbf1d9f5800d92b3fae86edf8b29993930dd06e7ecdcffacf212 = 
        y_nr_in[26] ^ 
        y_nr_in[38] ^ 
        y_nr_in[0] ^ 
0; 



wire I766ae41e1b152fe6af0be4a78b9e7ba001ff2936caefb0a89a2e11b1cf91164e;
assign I766ae41e1b152fe6af0be4a78b9e7ba001ff2936caefb0a89a2e11b1cf91164e = 
        y_nr_in[15] ^ 
        y_nr_in[18] ^ 
        y_nr_in[22] ^ 
0; 



wire I911547b3d7cbd99015ec8e23a3a6e6b06c4ddd5caaa2028dff9e2b255d80e5fb;
assign I911547b3d7cbd99015ec8e23a3a6e6b06c4ddd5caaa2028dff9e2b255d80e5fb = 
        y_nr_in[27] ^ 
        y_nr_in[29] ^ 
        y_nr_in[33] ^ 
0; 



wire Ia1648355a668c98d3e56d22e8820c317ba6743a0872fc63d27abe88bb38baba6;
assign Ia1648355a668c98d3e56d22e8820c317ba6743a0872fc63d27abe88bb38baba6 = 
        y_nr_in[37] ^ 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
0; 



wire Ic4e8b9cc64bed9afb08f97c676d674c833beee78ab59c6fc96068c46bbf2cafc;
assign Ic4e8b9cc64bed9afb08f97c676d674c833beee78ab59c6fc96068c46bbf2cafc = 
        y_nr_in[13] ^ 
        y_nr_in[17] ^ 
        y_nr_in[33] ^ 
0; 



wire Ic88c1bc4702c8cebbc502460e20db86b9b99a15a34413f84468bd6da387369e7;
assign Ic88c1bc4702c8cebbc502460e20db86b9b99a15a34413f84468bd6da387369e7 = 
        y_nr_in[5] ^ 
        y_nr_in[11] ^ 
        y_nr_in[19] ^ 
0; 



wire Iec133d23e39923dfbc21a1414e142bbe841a5f151d6fde6d9916a908ca75374a;
assign Iec133d23e39923dfbc21a1414e142bbe841a5f151d6fde6d9916a908ca75374a = 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
        y_nr_in[31] ^ 
0; 



wire Ic3878a882e9c8548378475efc42a603d8af9be1ab6319a5af2907c71bd255aea;
assign Ic3878a882e9c8548378475efc42a603d8af9be1ab6319a5af2907c71bd255aea = 
        y_nr_in[35] ^ 
        y_nr_in[37] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[166] = 
Iac791f5d19a7c542254f5d4b9b0fa6eef7eeb9b06f8a9916a3dc9da1bbda42ba ^ 
Ie88a242b25c2fbf1d9f5800d92b3fae86edf8b29993930dd06e7ecdcffacf212 ^ 
I766ae41e1b152fe6af0be4a78b9e7ba001ff2936caefb0a89a2e11b1cf91164e ^ 
I911547b3d7cbd99015ec8e23a3a6e6b06c4ddd5caaa2028dff9e2b255d80e5fb ^ 
Ia1648355a668c98d3e56d22e8820c317ba6743a0872fc63d27abe88bb38baba6 ^ 
Ic4e8b9cc64bed9afb08f97c676d674c833beee78ab59c6fc96068c46bbf2cafc ^ 
Ic88c1bc4702c8cebbc502460e20db86b9b99a15a34413f84468bd6da387369e7 ^ 
Iec133d23e39923dfbc21a1414e142bbe841a5f151d6fde6d9916a908ca75374a ^ 
Ic3878a882e9c8548378475efc42a603d8af9be1ab6319a5af2907c71bd255aea ^ 
0; 



wire If1ee4ad64aeb58b31a2d63964b9e7d9ed3262b98d14da43b315d4fe70ed9f413;
assign If1ee4ad64aeb58b31a2d63964b9e7d9ed3262b98d14da43b315d4fe70ed9f413 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[12] ^ 
0; 



wire I729ab5e0f24be138808d0f0fb1a85c34068d17c0444ed6e7ec150b8cf2321902;
assign I729ab5e0f24be138808d0f0fb1a85c34068d17c0444ed6e7ec150b8cf2321902 = 
        y_nr_in[27] ^ 
        y_nr_in[39] ^ 
        y_nr_in[1] ^ 
0; 



wire I84aebfe4105a92659656af779927dd1c1d6b1319e04926a29a8c5bfb6efdf6c6;
assign I84aebfe4105a92659656af779927dd1c1d6b1319e04926a29a8c5bfb6efdf6c6 = 
        y_nr_in[12] ^ 
        y_nr_in[19] ^ 
        y_nr_in[23] ^ 
0; 



wire I5ac9293e51815e81a2ea43e6c0c2f4584e8aa92468263844f22dd277bf20fb02;
assign I5ac9293e51815e81a2ea43e6c0c2f4584e8aa92468263844f22dd277bf20fb02 = 
        y_nr_in[24] ^ 
        y_nr_in[30] ^ 
        y_nr_in[34] ^ 
0; 



wire I4a19e53822fe615bcf1cc74ecac7740aa492ed3d3ff52c57c9919d1732b2de48;
assign I4a19e53822fe615bcf1cc74ecac7740aa492ed3d3ff52c57c9919d1732b2de48 = 
        y_nr_in[38] ^ 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
0; 



wire I16df24cc348fcf594db15ecd1a08146f675c8eb4df138cfaf07c25ff158d742b;
assign I16df24cc348fcf594db15ecd1a08146f675c8eb4df138cfaf07c25ff158d742b = 
        y_nr_in[14] ^ 
        y_nr_in[18] ^ 
        y_nr_in[34] ^ 
0; 



wire Ib03c7e791e07d151d6a84b1c5be1df0998d5506c3eb948da9b640e4afccce94a;
assign Ib03c7e791e07d151d6a84b1c5be1df0998d5506c3eb948da9b640e4afccce94a = 
        y_nr_in[6] ^ 
        y_nr_in[8] ^ 
        y_nr_in[16] ^ 
0; 



wire I8dbaa75663c0e825b23f8c64b580d645b8aafc883c4720b64ac8da7213433578;
assign I8dbaa75663c0e825b23f8c64b580d645b8aafc883c4720b64ac8da7213433578 = 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
        y_nr_in[28] ^ 
0; 



wire I813485e1705cedefbbb872d49c8c3f55c6d0c6440e0b31444f6b9e5e8a0b720b;
assign I813485e1705cedefbbb872d49c8c3f55c6d0c6440e0b31444f6b9e5e8a0b720b = 
        y_nr_in[32] ^ 
        y_nr_in[38] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[165] = 
If1ee4ad64aeb58b31a2d63964b9e7d9ed3262b98d14da43b315d4fe70ed9f413 ^ 
I729ab5e0f24be138808d0f0fb1a85c34068d17c0444ed6e7ec150b8cf2321902 ^ 
I84aebfe4105a92659656af779927dd1c1d6b1319e04926a29a8c5bfb6efdf6c6 ^ 
I5ac9293e51815e81a2ea43e6c0c2f4584e8aa92468263844f22dd277bf20fb02 ^ 
I4a19e53822fe615bcf1cc74ecac7740aa492ed3d3ff52c57c9919d1732b2de48 ^ 
I16df24cc348fcf594db15ecd1a08146f675c8eb4df138cfaf07c25ff158d742b ^ 
Ib03c7e791e07d151d6a84b1c5be1df0998d5506c3eb948da9b640e4afccce94a ^ 
I8dbaa75663c0e825b23f8c64b580d645b8aafc883c4720b64ac8da7213433578 ^ 
I813485e1705cedefbbb872d49c8c3f55c6d0c6440e0b31444f6b9e5e8a0b720b ^ 
0; 



wire I2b7edf8e0a2ea23cfc68797e318e75ad0d62c5279dcdd15f1f16f72c4f231745;
assign I2b7edf8e0a2ea23cfc68797e318e75ad0d62c5279dcdd15f1f16f72c4f231745 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[13] ^ 
0; 



wire I6b654dceb4abb2d4f4117292e4abb82ad4736884245d9359716dd64171ce075c;
assign I6b654dceb4abb2d4f4117292e4abb82ad4736884245d9359716dd64171ce075c = 
        y_nr_in[24] ^ 
        y_nr_in[36] ^ 
        y_nr_in[2] ^ 
0; 



wire Ic9e20741342ac8d9e0b5c8064d33d674dc1830a2133c46972aba04b17f31e762;
assign Ic9e20741342ac8d9e0b5c8064d33d674dc1830a2133c46972aba04b17f31e762 = 
        y_nr_in[13] ^ 
        y_nr_in[16] ^ 
        y_nr_in[20] ^ 
0; 



wire Ia6bd1e117f94aabde2317aaf6edf0b629665320453de800a6e09c5ca6f21728d;
assign Ia6bd1e117f94aabde2317aaf6edf0b629665320453de800a6e09c5ca6f21728d = 
        y_nr_in[25] ^ 
        y_nr_in[31] ^ 
        y_nr_in[35] ^ 
0; 



wire I2b498074090142494a2e0080a3bb631d5a04e85a75d56ce1cef04a4afbb139e0;
assign I2b498074090142494a2e0080a3bb631d5a04e85a75d56ce1cef04a4afbb139e0 = 
        y_nr_in[39] ^ 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
0; 



wire I9ed7ab2137031f54c9e57d9615a4f20cb8f09375f8b6a469ff0fc872ca300220;
assign I9ed7ab2137031f54c9e57d9615a4f20cb8f09375f8b6a469ff0fc872ca300220 = 
        y_nr_in[15] ^ 
        y_nr_in[19] ^ 
        y_nr_in[35] ^ 
0; 



wire Ie3e896f4aed44b3afadc325f55877e9d622c081545cf83aa93163b110ce8577a;
assign Ie3e896f4aed44b3afadc325f55877e9d622c081545cf83aa93163b110ce8577a = 
        y_nr_in[7] ^ 
        y_nr_in[9] ^ 
        y_nr_in[17] ^ 
0; 



wire Ie0011f08acb9bb4b4ee59ee1acb2c4e9de4a0be5e1be53c6b0af1c6b197abee2;
assign Ie0011f08acb9bb4b4ee59ee1acb2c4e9de4a0be5e1be53c6b0af1c6b197abee2 = 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
        y_nr_in[29] ^ 
0; 



wire I98f1b83559e42ab63f837f32ba11ed46b81066a22308a8858013a2e14066d38a;
assign I98f1b83559e42ab63f837f32ba11ed46b81066a22308a8858013a2e14066d38a = 
        y_nr_in[33] ^ 
        y_nr_in[39] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[164] = 
I2b7edf8e0a2ea23cfc68797e318e75ad0d62c5279dcdd15f1f16f72c4f231745 ^ 
I6b654dceb4abb2d4f4117292e4abb82ad4736884245d9359716dd64171ce075c ^ 
Ic9e20741342ac8d9e0b5c8064d33d674dc1830a2133c46972aba04b17f31e762 ^ 
Ia6bd1e117f94aabde2317aaf6edf0b629665320453de800a6e09c5ca6f21728d ^ 
I2b498074090142494a2e0080a3bb631d5a04e85a75d56ce1cef04a4afbb139e0 ^ 
I9ed7ab2137031f54c9e57d9615a4f20cb8f09375f8b6a469ff0fc872ca300220 ^ 
Ie3e896f4aed44b3afadc325f55877e9d622c081545cf83aa93163b110ce8577a ^ 
Ie0011f08acb9bb4b4ee59ee1acb2c4e9de4a0be5e1be53c6b0af1c6b197abee2 ^ 
I98f1b83559e42ab63f837f32ba11ed46b81066a22308a8858013a2e14066d38a ^ 
0; 



wire I66114ebf49758b85fa88173cde89be4e76b7d35cadcea53c73018b32c968928e;
assign I66114ebf49758b85fa88173cde89be4e76b7d35cadcea53c73018b32c968928e = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[14] ^ 
0; 



wire I09ab146dcfc299eb45c496708ef501ae7adaddb3366bc9346fe2d0787a2462ad;
assign I09ab146dcfc299eb45c496708ef501ae7adaddb3366bc9346fe2d0787a2462ad = 
        y_nr_in[25] ^ 
        y_nr_in[37] ^ 
        y_nr_in[40] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[163] = 
I66114ebf49758b85fa88173cde89be4e76b7d35cadcea53c73018b32c968928e ^ 
I09ab146dcfc299eb45c496708ef501ae7adaddb3366bc9346fe2d0787a2462ad ^ 
0; 



wire I85d19610152535540624bce37e88a0212ea10e49076fa932cf011349f6047bf0;
assign I85d19610152535540624bce37e88a0212ea10e49076fa932cf011349f6047bf0 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[15] ^ 
0; 



wire I64791be3ad9109e626afa75a98c8d0d792149c1d54016881809da5af04a0e384;
assign I64791be3ad9109e626afa75a98c8d0d792149c1d54016881809da5af04a0e384 = 
        y_nr_in[26] ^ 
        y_nr_in[38] ^ 
        y_nr_in[41] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[162] = 
I85d19610152535540624bce37e88a0212ea10e49076fa932cf011349f6047bf0 ^ 
I64791be3ad9109e626afa75a98c8d0d792149c1d54016881809da5af04a0e384 ^ 
0; 



wire Ib1b3643dc8b0921d548e81b347057dc6dd4d5ad184fc51c67819bfe36308f9c3;
assign Ib1b3643dc8b0921d548e81b347057dc6dd4d5ad184fc51c67819bfe36308f9c3 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[12] ^ 
0; 



wire I3f46b46cdea70163ead954ce7cddb9426ca8af6c4ba1cd67fb81b25318dd1a51;
assign I3f46b46cdea70163ead954ce7cddb9426ca8af6c4ba1cd67fb81b25318dd1a51 = 
        y_nr_in[27] ^ 
        y_nr_in[39] ^ 
        y_nr_in[42] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[161] = 
Ib1b3643dc8b0921d548e81b347057dc6dd4d5ad184fc51c67819bfe36308f9c3 ^ 
I3f46b46cdea70163ead954ce7cddb9426ca8af6c4ba1cd67fb81b25318dd1a51 ^ 
0; 



wire I98abd59ea45c34049379ee6f12c587b30a1da4de32d3070f7e69adc0f9fc4f4c;
assign I98abd59ea45c34049379ee6f12c587b30a1da4de32d3070f7e69adc0f9fc4f4c = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[13] ^ 
0; 



wire I575f70d8cdf578436f1c4a28df7193c167c3afad67d511e7a50ea08ee201328e;
assign I575f70d8cdf578436f1c4a28df7193c167c3afad67d511e7a50ea08ee201328e = 
        y_nr_in[24] ^ 
        y_nr_in[36] ^ 
        y_nr_in[43] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[160] = 
I98abd59ea45c34049379ee6f12c587b30a1da4de32d3070f7e69adc0f9fc4f4c ^ 
I575f70d8cdf578436f1c4a28df7193c167c3afad67d511e7a50ea08ee201328e ^ 
0; 



wire I9e6675aa0733abe263e12611ab91432a8c0c8845b2cc6470c0892e4bf592b952;
assign I9e6675aa0733abe263e12611ab91432a8c0c8845b2cc6470c0892e4bf592b952 = 
        y_nr_in[3] ^ 
        y_nr_in[14] ^ 
        y_nr_in[17] ^ 
0; 



wire Ic08db7865858b018e4d903e6cede7fa6fdfc2835c63b14879defaec28ca05954;
assign Ic08db7865858b018e4d903e6cede7fa6fdfc2835c63b14879defaec28ca05954 = 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
        y_nr_in[28] ^ 
0; 



wire If08bdc3b48c23f2a579be4139c5a8720039e7d9b87d1ea781c9ab522b92465cd;
assign If08bdc3b48c23f2a579be4139c5a8720039e7d9b87d1ea781c9ab522b92465cd = 
        y_nr_in[32] ^ 
        y_nr_in[36] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[159] = 
I9e6675aa0733abe263e12611ab91432a8c0c8845b2cc6470c0892e4bf592b952 ^ 
Ic08db7865858b018e4d903e6cede7fa6fdfc2835c63b14879defaec28ca05954 ^ 
If08bdc3b48c23f2a579be4139c5a8720039e7d9b87d1ea781c9ab522b92465cd ^ 
0; 



wire I6de6fe4c522d22a10ebba344a52da5f9938ab78ea1170471deda3bda1568dee4;
assign I6de6fe4c522d22a10ebba344a52da5f9938ab78ea1170471deda3bda1568dee4 = 
        y_nr_in[0] ^ 
        y_nr_in[15] ^ 
        y_nr_in[18] ^ 
0; 



wire Ie18ab9008e399fd861af074e7dcf889c783cbbf155b7e26bcc291d5e450ec47c;
assign Ie18ab9008e399fd861af074e7dcf889c783cbbf155b7e26bcc291d5e450ec47c = 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
        y_nr_in[29] ^ 
0; 



wire Ic6cd571ce4830c9b73cb3817606c2f0c642a40e0120a852b51ce8fd84a460976;
assign Ic6cd571ce4830c9b73cb3817606c2f0c642a40e0120a852b51ce8fd84a460976 = 
        y_nr_in[33] ^ 
        y_nr_in[37] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[158] = 
I6de6fe4c522d22a10ebba344a52da5f9938ab78ea1170471deda3bda1568dee4 ^ 
Ie18ab9008e399fd861af074e7dcf889c783cbbf155b7e26bcc291d5e450ec47c ^ 
Ic6cd571ce4830c9b73cb3817606c2f0c642a40e0120a852b51ce8fd84a460976 ^ 
0; 



wire Ic0dedd09d29bc666a177c4f8f1aac7e081134411a025698ffe952de1a47cd4ea;
assign Ic0dedd09d29bc666a177c4f8f1aac7e081134411a025698ffe952de1a47cd4ea = 
        y_nr_in[1] ^ 
        y_nr_in[12] ^ 
        y_nr_in[19] ^ 
0; 



wire I7033877127d107f386702d703bbf5d09944327b54c344a2183ab59432f1dd38b;
assign I7033877127d107f386702d703bbf5d09944327b54c344a2183ab59432f1dd38b = 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
        y_nr_in[30] ^ 
0; 



wire I83847df0ccc11aee3bcc85c5799fe02fc69b9b11d418093ba0e48edf0ca638c9;
assign I83847df0ccc11aee3bcc85c5799fe02fc69b9b11d418093ba0e48edf0ca638c9 = 
        y_nr_in[34] ^ 
        y_nr_in[38] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[157] = 
Ic0dedd09d29bc666a177c4f8f1aac7e081134411a025698ffe952de1a47cd4ea ^ 
I7033877127d107f386702d703bbf5d09944327b54c344a2183ab59432f1dd38b ^ 
I83847df0ccc11aee3bcc85c5799fe02fc69b9b11d418093ba0e48edf0ca638c9 ^ 
0; 



wire Ifc905cf9062222c11f5bd5d42856c5cd90aef46202ad17cac28de6a4c79188a0;
assign Ifc905cf9062222c11f5bd5d42856c5cd90aef46202ad17cac28de6a4c79188a0 = 
        y_nr_in[2] ^ 
        y_nr_in[13] ^ 
        y_nr_in[16] ^ 
0; 



wire Iabcae1466aca23a97807b870802432b1a9133e9c5b1107af1d17fa29ae2349fa;
assign Iabcae1466aca23a97807b870802432b1a9133e9c5b1107af1d17fa29ae2349fa = 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
        y_nr_in[31] ^ 
0; 



wire I38cfc35692114c0f78eb7e848455037e75419c4d94f9ae7b0bd34be92148d822;
assign I38cfc35692114c0f78eb7e848455037e75419c4d94f9ae7b0bd34be92148d822 = 
        y_nr_in[35] ^ 
        y_nr_in[39] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[156] = 
Ifc905cf9062222c11f5bd5d42856c5cd90aef46202ad17cac28de6a4c79188a0 ^ 
Iabcae1466aca23a97807b870802432b1a9133e9c5b1107af1d17fa29ae2349fa ^ 
I38cfc35692114c0f78eb7e848455037e75419c4d94f9ae7b0bd34be92148d822 ^ 
0; 



wire I39b9e146b624c47c64074bc132b83b1c4753edc20128f1b570ce586aa990a361;
assign I39b9e146b624c47c64074bc132b83b1c4753edc20128f1b570ce586aa990a361 = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[12] ^ 
0; 



wire If4782b9a6f137d441f49270c1f5792c3c82aa0b4181f102fd829d34e92908a18;
assign If4782b9a6f137d441f49270c1f5792c3c82aa0b4181f102fd829d34e92908a18 = 
        y_nr_in[16] ^ 
        y_nr_in[32] ^ 
        y_nr_in[41] ^ 
0; 



wire Ic9ac5fae78e4edf3f4386d3b9e6413586e877b674b4bd58b0901afe2bcd4fad1;
assign Ic9ac5fae78e4edf3f4386d3b9e6413586e877b674b4bd58b0901afe2bcd4fad1 = 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[155] = 
I39b9e146b624c47c64074bc132b83b1c4753edc20128f1b570ce586aa990a361 ^ 
If4782b9a6f137d441f49270c1f5792c3c82aa0b4181f102fd829d34e92908a18 ^ 
Ic9ac5fae78e4edf3f4386d3b9e6413586e877b674b4bd58b0901afe2bcd4fad1 ^ 
0; 



wire I8c2a7cade24a98f62797ff246db0618e2031ec48015c9fbfdf2d6559c0536377;
assign I8c2a7cade24a98f62797ff246db0618e2031ec48015c9fbfdf2d6559c0536377 = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[13] ^ 
0; 



wire Ic69d76766fb488361fb56fd190a88a81f06803c8d1716f0253c485b72feaac53;
assign Ic69d76766fb488361fb56fd190a88a81f06803c8d1716f0253c485b72feaac53 = 
        y_nr_in[17] ^ 
        y_nr_in[33] ^ 
        y_nr_in[42] ^ 
0; 



wire I1e2311c30ff9a73dc61dec199bf6b3ab33c14e1f7f8c10019ce05e5e3b0ee413;
assign I1e2311c30ff9a73dc61dec199bf6b3ab33c14e1f7f8c10019ce05e5e3b0ee413 = 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[154] = 
I8c2a7cade24a98f62797ff246db0618e2031ec48015c9fbfdf2d6559c0536377 ^ 
Ic69d76766fb488361fb56fd190a88a81f06803c8d1716f0253c485b72feaac53 ^ 
I1e2311c30ff9a73dc61dec199bf6b3ab33c14e1f7f8c10019ce05e5e3b0ee413 ^ 
0; 



wire I76ce9b3a35c82ecffdcbed87005640a6ffdf4cbb54e8d0280fe0fe1a47ec4153;
assign I76ce9b3a35c82ecffdcbed87005640a6ffdf4cbb54e8d0280fe0fe1a47ec4153 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[14] ^ 
0; 



wire I4708468f8391617733b308fac7685318e53210aa0cb4c54f84eae68f5df5a979;
assign I4708468f8391617733b308fac7685318e53210aa0cb4c54f84eae68f5df5a979 = 
        y_nr_in[18] ^ 
        y_nr_in[34] ^ 
        y_nr_in[43] ^ 
0; 



wire I559b8de6e88c7999fd1658a92374e26f146bc56347af825b373e8c3c3c94bfe6;
assign I559b8de6e88c7999fd1658a92374e26f146bc56347af825b373e8c3c3c94bfe6 = 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[153] = 
I76ce9b3a35c82ecffdcbed87005640a6ffdf4cbb54e8d0280fe0fe1a47ec4153 ^ 
I4708468f8391617733b308fac7685318e53210aa0cb4c54f84eae68f5df5a979 ^ 
I559b8de6e88c7999fd1658a92374e26f146bc56347af825b373e8c3c3c94bfe6 ^ 
0; 



wire Icec9f82ed5458da4eeaed077c58e91d3501f3067dda84ffba55bf76aee5404cd;
assign Icec9f82ed5458da4eeaed077c58e91d3501f3067dda84ffba55bf76aee5404cd = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[15] ^ 
0; 



wire I8f0d9addae8d828d43015c922d7333c89906db27ab32fca73f81c54315c9bfde;
assign I8f0d9addae8d828d43015c922d7333c89906db27ab32fca73f81c54315c9bfde = 
        y_nr_in[19] ^ 
        y_nr_in[35] ^ 
        y_nr_in[40] ^ 
0; 



wire I040fabcf8c64dc85058af7c3ac6037167e279bb0f1bbc4885341f854d85a7b7f;
assign I040fabcf8c64dc85058af7c3ac6037167e279bb0f1bbc4885341f854d85a7b7f = 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[152] = 
Icec9f82ed5458da4eeaed077c58e91d3501f3067dda84ffba55bf76aee5404cd ^ 
I8f0d9addae8d828d43015c922d7333c89906db27ab32fca73f81c54315c9bfde ^ 
I040fabcf8c64dc85058af7c3ac6037167e279bb0f1bbc4885341f854d85a7b7f ^ 
0; 



wire Ica3e70c51fbbb23af567352e4d10f1931a92bbfe1e3ea9d9888a9fd29b207813;
assign Ica3e70c51fbbb23af567352e4d10f1931a92bbfe1e3ea9d9888a9fd29b207813 = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[151] = 
Ica3e70c51fbbb23af567352e4d10f1931a92bbfe1e3ea9d9888a9fd29b207813 ^ 
0; 



wire Ifa3c0791921cff838fa1d35eed6744fd64727fc362c31d54baa6fc3d8cff13d2;
assign Ifa3c0791921cff838fa1d35eed6744fd64727fc362c31d54baa6fc3d8cff13d2 = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[150] = 
Ifa3c0791921cff838fa1d35eed6744fd64727fc362c31d54baa6fc3d8cff13d2 ^ 
0; 



wire Idc56dcfa439c82ce544cec043fbb3f4b4ff644879ce68c071c6247ea236e1071;
assign Idc56dcfa439c82ce544cec043fbb3f4b4ff644879ce68c071c6247ea236e1071 = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[149] = 
Idc56dcfa439c82ce544cec043fbb3f4b4ff644879ce68c071c6247ea236e1071 ^ 
0; 



wire I1e29ad7126c9994135a12ef7507fa4d7988055cc266445a55effbf6de0a0bf1a;
assign I1e29ad7126c9994135a12ef7507fa4d7988055cc266445a55effbf6de0a0bf1a = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[148] = 
I1e29ad7126c9994135a12ef7507fa4d7988055cc266445a55effbf6de0a0bf1a ^ 
0; 



wire Ic80cfcf328cef7e9932b182f78996b4571cd505fce91f1bc6e1558c98751dc19;
assign Ic80cfcf328cef7e9932b182f78996b4571cd505fce91f1bc6e1558c98751dc19 = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[22] ^ 
0; 



wire Ib32fbf2ce5ebae1700f9ed1264dc6ccec4d49d411a6d0333aea050ce8139b610;
assign Ib32fbf2ce5ebae1700f9ed1264dc6ccec4d49d411a6d0333aea050ce8139b610 = 
        y_nr_in[31] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[147] = 
Ic80cfcf328cef7e9932b182f78996b4571cd505fce91f1bc6e1558c98751dc19 ^ 
Ib32fbf2ce5ebae1700f9ed1264dc6ccec4d49d411a6d0333aea050ce8139b610 ^ 
0; 



wire I4537c147914b240750383c57700b9c4687a349f441c6fda2c8ab80aa93ec8272;
assign I4537c147914b240750383c57700b9c4687a349f441c6fda2c8ab80aa93ec8272 = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[23] ^ 
0; 



wire Ic358968cbf334449efb91fe3a98a6228903c5c0bef6f2e81cfca8cd8735984d0;
assign Ic358968cbf334449efb91fe3a98a6228903c5c0bef6f2e81cfca8cd8735984d0 = 
        y_nr_in[28] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[146] = 
I4537c147914b240750383c57700b9c4687a349f441c6fda2c8ab80aa93ec8272 ^ 
Ic358968cbf334449efb91fe3a98a6228903c5c0bef6f2e81cfca8cd8735984d0 ^ 
0; 



wire Ie32b6bd5e13ab6e0255cfa736314da54c7eb2ed64454f351be4fc653cc73ad3d;
assign Ie32b6bd5e13ab6e0255cfa736314da54c7eb2ed64454f351be4fc653cc73ad3d = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[20] ^ 
0; 



wire If4991a5d7d21efa79dc59a917034abd85e727ca8e4d68922a3ba80b6dafeed93;
assign If4991a5d7d21efa79dc59a917034abd85e727ca8e4d68922a3ba80b6dafeed93 = 
        y_nr_in[29] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[145] = 
Ie32b6bd5e13ab6e0255cfa736314da54c7eb2ed64454f351be4fc653cc73ad3d ^ 
If4991a5d7d21efa79dc59a917034abd85e727ca8e4d68922a3ba80b6dafeed93 ^ 
0; 



wire Ie2e2b08e080a117ff65e7040ffa15e72db6c1310243629d972c7139b0f5a3c05;
assign Ie2e2b08e080a117ff65e7040ffa15e72db6c1310243629d972c7139b0f5a3c05 = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[21] ^ 
0; 



wire I684fc51d495fedfd9bdafe94485a2cd8688ee121e5c2978bab87f9fd4e37d80b;
assign I684fc51d495fedfd9bdafe94485a2cd8688ee121e5c2978bab87f9fd4e37d80b = 
        y_nr_in[30] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[144] = 
Ie2e2b08e080a117ff65e7040ffa15e72db6c1310243629d972c7139b0f5a3c05 ^ 
I684fc51d495fedfd9bdafe94485a2cd8688ee121e5c2978bab87f9fd4e37d80b ^ 
0; 



wire Icd559c515beaeb5e638188f70e32299ef43943b0ce1d19e80f29eba0679bee12;
assign Icd559c515beaeb5e638188f70e32299ef43943b0ce1d19e80f29eba0679bee12 = 
        y_nr_in[3] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
0; 



wire I9b85a437b6ccee7b3eb0bb207780c3ac9d23084c0717639c860e0eede8ceb424;
assign I9b85a437b6ccee7b3eb0bb207780c3ac9d23084c0717639c860e0eede8ceb424 = 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[143] = 
Icd559c515beaeb5e638188f70e32299ef43943b0ce1d19e80f29eba0679bee12 ^ 
I9b85a437b6ccee7b3eb0bb207780c3ac9d23084c0717639c860e0eede8ceb424 ^ 
0; 



wire Ieffbeb4c9fb0242ffc90388bc5d16c0c78b4062ddbdfbb930493030a31fbc952;
assign Ieffbeb4c9fb0242ffc90388bc5d16c0c78b4062ddbdfbb930493030a31fbc952 = 
        y_nr_in[0] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
0; 



wire I432a5b3a6f7b766c46f38fa8352f92193958b9b99b3303b9de56ca31d1e02cac;
assign I432a5b3a6f7b766c46f38fa8352f92193958b9b99b3303b9de56ca31d1e02cac = 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[142] = 
Ieffbeb4c9fb0242ffc90388bc5d16c0c78b4062ddbdfbb930493030a31fbc952 ^ 
I432a5b3a6f7b766c46f38fa8352f92193958b9b99b3303b9de56ca31d1e02cac ^ 
0; 



wire I92b68e093194b90a895bbcb5099de8d29c6794a60a577d4eed46d76e9b32c771;
assign I92b68e093194b90a895bbcb5099de8d29c6794a60a577d4eed46d76e9b32c771 = 
        y_nr_in[1] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
0; 



wire I8e6aa109e626ccf41e30d5be046926ea4911a5c96c395439be996defe16abedd;
assign I8e6aa109e626ccf41e30d5be046926ea4911a5c96c395439be996defe16abedd = 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[141] = 
I92b68e093194b90a895bbcb5099de8d29c6794a60a577d4eed46d76e9b32c771 ^ 
I8e6aa109e626ccf41e30d5be046926ea4911a5c96c395439be996defe16abedd ^ 
0; 



wire Ib76ac2efd49415c33cd7fcdf86117582203844469bef6fb1aa6f18900ca60a5c;
assign Ib76ac2efd49415c33cd7fcdf86117582203844469bef6fb1aa6f18900ca60a5c = 
        y_nr_in[2] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
0; 



wire I03b405c1cc83c255c00b4083014452478f0a29d2c8627b935765fd2a2aacb8c7;
assign I03b405c1cc83c255c00b4083014452478f0a29d2c8627b935765fd2a2aacb8c7 = 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[140] = 
Ib76ac2efd49415c33cd7fcdf86117582203844469bef6fb1aa6f18900ca60a5c ^ 
I03b405c1cc83c255c00b4083014452478f0a29d2c8627b935765fd2a2aacb8c7 ^ 
0; 



wire If0fdcc606689de54b4d5c073b32361cd4e2dd18918d442f8ba79f91104fdb8d1;
assign If0fdcc606689de54b4d5c073b32361cd4e2dd18918d442f8ba79f91104fdb8d1 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
0; 



wire I0ae1486b18345160a62ea7f5aae0f08023802f01b5e5a8c25a66341390f7e985;
assign I0ae1486b18345160a62ea7f5aae0f08023802f01b5e5a8c25a66341390f7e985 = 
        y_nr_in[47] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[139] = 
If0fdcc606689de54b4d5c073b32361cd4e2dd18918d442f8ba79f91104fdb8d1 ^ 
I0ae1486b18345160a62ea7f5aae0f08023802f01b5e5a8c25a66341390f7e985 ^ 
0; 



wire Ia304d4a11073812e03c60d974ce8263b191a6a8e0e607016cb97e203e1ce574c;
assign Ia304d4a11073812e03c60d974ce8263b191a6a8e0e607016cb97e203e1ce574c = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
0; 



wire Ifd4d0c5293adb43eef92c64f186765fd3f7e65fbc89c2eb7d8cc142bb6fc133a;
assign Ifd4d0c5293adb43eef92c64f186765fd3f7e65fbc89c2eb7d8cc142bb6fc133a = 
        y_nr_in[44] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[138] = 
Ia304d4a11073812e03c60d974ce8263b191a6a8e0e607016cb97e203e1ce574c ^ 
Ifd4d0c5293adb43eef92c64f186765fd3f7e65fbc89c2eb7d8cc142bb6fc133a ^ 
0; 



wire I5a2c723ed8fd3c3a348a0c101a5dc19af4119ed12bf2e21b4a99534a0f4c685b;
assign I5a2c723ed8fd3c3a348a0c101a5dc19af4119ed12bf2e21b4a99534a0f4c685b = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
0; 



wire I55b033f99a170527e217f660dfcaf4f9161f15bae2cdb4a559a487ff4677528a;
assign I55b033f99a170527e217f660dfcaf4f9161f15bae2cdb4a559a487ff4677528a = 
        y_nr_in[45] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[137] = 
I5a2c723ed8fd3c3a348a0c101a5dc19af4119ed12bf2e21b4a99534a0f4c685b ^ 
I55b033f99a170527e217f660dfcaf4f9161f15bae2cdb4a559a487ff4677528a ^ 
0; 



wire I68abd03f6b7e831232b1811637b67182a1547f4b49ce74bf3c64be5d8c92a353;
assign I68abd03f6b7e831232b1811637b67182a1547f4b49ce74bf3c64be5d8c92a353 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
0; 



wire I21b5c839087fd1584cd5e0c684d1e6f8c5e191e24144d1f5ed36d1354863d459;
assign I21b5c839087fd1584cd5e0c684d1e6f8c5e191e24144d1f5ed36d1354863d459 = 
        y_nr_in[46] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[136] = 
I68abd03f6b7e831232b1811637b67182a1547f4b49ce74bf3c64be5d8c92a353 ^ 
I21b5c839087fd1584cd5e0c684d1e6f8c5e191e24144d1f5ed36d1354863d459 ^ 
0; 



wire I9036d79d85649603ba008bee293e9a61721de8dfb3ea0c780caf8befb8c59da2;
assign I9036d79d85649603ba008bee293e9a61721de8dfb3ea0c780caf8befb8c59da2 = 
        y_nr_in[2] ^ 
        y_nr_in[6] ^ 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[135] = 
I9036d79d85649603ba008bee293e9a61721de8dfb3ea0c780caf8befb8c59da2 ^ 
0; 



wire I8723d833aaa6375f50399022729689f26a214a6d3386577cbe76e43bfaead2f9;
assign I8723d833aaa6375f50399022729689f26a214a6d3386577cbe76e43bfaead2f9 = 
        y_nr_in[3] ^ 
        y_nr_in[7] ^ 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[134] = 
I8723d833aaa6375f50399022729689f26a214a6d3386577cbe76e43bfaead2f9 ^ 
0; 



wire I6b6989abe368b02139bf779aa6bd0ea63a67a493bf3a170d2fe37b0f62462b7b;
assign I6b6989abe368b02139bf779aa6bd0ea63a67a493bf3a170d2fe37b0f62462b7b = 
        y_nr_in[0] ^ 
        y_nr_in[4] ^ 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[133] = 
I6b6989abe368b02139bf779aa6bd0ea63a67a493bf3a170d2fe37b0f62462b7b ^ 
0; 



wire I0808f3f511663abe7288885dd511c482c1b6b7f8bff3b15b4a791e9004c78b75;
assign I0808f3f511663abe7288885dd511c482c1b6b7f8bff3b15b4a791e9004c78b75 = 
        y_nr_in[1] ^ 
        y_nr_in[5] ^ 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[132] = 
I0808f3f511663abe7288885dd511c482c1b6b7f8bff3b15b4a791e9004c78b75 ^ 
0; 



wire I54b1cfe31e5bd3dbbd4fa7c0e7800e1690c59de900c6dc0fe6045bff598d6972;
assign I54b1cfe31e5bd3dbbd4fa7c0e7800e1690c59de900c6dc0fe6045bff598d6972 = 
        y_nr_in[7] ^ 
        y_nr_in[33] ^ 
        y_nr_in[41] ^ 
0; 



wire Ib251b7951905b6876a85ea96e1feae5cb5a86a410589c43796edba5db8616ad8;
assign Ib251b7951905b6876a85ea96e1feae5cb5a86a410589c43796edba5db8616ad8 = 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[131] = 
I54b1cfe31e5bd3dbbd4fa7c0e7800e1690c59de900c6dc0fe6045bff598d6972 ^ 
Ib251b7951905b6876a85ea96e1feae5cb5a86a410589c43796edba5db8616ad8 ^ 
0; 



wire Ifdeff48f8f63ae1b707c6d44f01b027e2fb439655b8f09b37027edd781ee975e;
assign Ifdeff48f8f63ae1b707c6d44f01b027e2fb439655b8f09b37027edd781ee975e = 
        y_nr_in[4] ^ 
        y_nr_in[34] ^ 
        y_nr_in[42] ^ 
0; 



wire I6a0b1d89dfcab30226aac89e1ed7c5d7da6d77a210e41e38a0d234369f386366;
assign I6a0b1d89dfcab30226aac89e1ed7c5d7da6d77a210e41e38a0d234369f386366 = 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[130] = 
Ifdeff48f8f63ae1b707c6d44f01b027e2fb439655b8f09b37027edd781ee975e ^ 
I6a0b1d89dfcab30226aac89e1ed7c5d7da6d77a210e41e38a0d234369f386366 ^ 
0; 



wire Iee83a9c6af510d609d531cafcc69628ca25af630d1b1c423885d4bbac737161f;
assign Iee83a9c6af510d609d531cafcc69628ca25af630d1b1c423885d4bbac737161f = 
        y_nr_in[5] ^ 
        y_nr_in[35] ^ 
        y_nr_in[43] ^ 
0; 



wire I924238012e56f966e02a2105a9fcb7acca5f7597114881270cd74a6aca4a3aca;
assign I924238012e56f966e02a2105a9fcb7acca5f7597114881270cd74a6aca4a3aca = 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[129] = 
Iee83a9c6af510d609d531cafcc69628ca25af630d1b1c423885d4bbac737161f ^ 
I924238012e56f966e02a2105a9fcb7acca5f7597114881270cd74a6aca4a3aca ^ 
0; 



wire I04e612eeeb21a866edeba1827f31fa3cfc5da5103261c5ff87c84c10b29e377d;
assign I04e612eeeb21a866edeba1827f31fa3cfc5da5103261c5ff87c84c10b29e377d = 
        y_nr_in[6] ^ 
        y_nr_in[32] ^ 
        y_nr_in[40] ^ 
0; 



wire Ifaed497c88df5e21d2c16270af29e46b6f0268d94489a891476049befca20a5a;
assign Ifaed497c88df5e21d2c16270af29e46b6f0268d94489a891476049befca20a5a = 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[128] = 
I04e612eeeb21a866edeba1827f31fa3cfc5da5103261c5ff87c84c10b29e377d ^ 
Ifaed497c88df5e21d2c16270af29e46b6f0268d94489a891476049befca20a5a ^ 
0; 



wire I0e0ac64caea92a1d75ed5a9ff960681180e0d9a0b5a7e7522163cd406b908016;
assign I0e0ac64caea92a1d75ed5a9ff960681180e0d9a0b5a7e7522163cd406b908016 = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[24] ^ 
0; 



wire I13329cf585ce2adddb84617f67bbccd866e1895fce56c3d3f606320150d64d2b;
assign I13329cf585ce2adddb84617f67bbccd866e1895fce56c3d3f606320150d64d2b = 
        y_nr_in[29] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[127] = 
I0e0ac64caea92a1d75ed5a9ff960681180e0d9a0b5a7e7522163cd406b908016 ^ 
I13329cf585ce2adddb84617f67bbccd866e1895fce56c3d3f606320150d64d2b ^ 
0; 



wire I6ae1ea820cf145f6e4643d41e39249c25380a19ccaa261f4cb5bc84ca04d1269;
assign I6ae1ea820cf145f6e4643d41e39249c25380a19ccaa261f4cb5bc84ca04d1269 = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[25] ^ 
0; 



wire I01c985d7b21c3404f2869130530caada54505fdd35e9f77a7f659b9401eb839b;
assign I01c985d7b21c3404f2869130530caada54505fdd35e9f77a7f659b9401eb839b = 
        y_nr_in[30] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[126] = 
I6ae1ea820cf145f6e4643d41e39249c25380a19ccaa261f4cb5bc84ca04d1269 ^ 
I01c985d7b21c3404f2869130530caada54505fdd35e9f77a7f659b9401eb839b ^ 
0; 



wire Icb2b0bd16431524939cdded20f245161f930c9c47942f8120e64560b9bc36d7b;
assign Icb2b0bd16431524939cdded20f245161f930c9c47942f8120e64560b9bc36d7b = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[26] ^ 
0; 



wire I6dc5f8037a6203884ca1d472f4228937785b19ab4c3a5bca62b0bbb44f4db717;
assign I6dc5f8037a6203884ca1d472f4228937785b19ab4c3a5bca62b0bbb44f4db717 = 
        y_nr_in[31] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[125] = 
Icb2b0bd16431524939cdded20f245161f930c9c47942f8120e64560b9bc36d7b ^ 
I6dc5f8037a6203884ca1d472f4228937785b19ab4c3a5bca62b0bbb44f4db717 ^ 
0; 



wire I09dd53def80e325c7ea5c3c8e2f064b02ebfe59c3b761e79a215a689b5e7cc40;
assign I09dd53def80e325c7ea5c3c8e2f064b02ebfe59c3b761e79a215a689b5e7cc40 = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[27] ^ 
0; 



wire Ic4ee10cf7e9ac1639974ed5497d880be058a326ee49d22970f95ada0e17981bd;
assign Ic4ee10cf7e9ac1639974ed5497d880be058a326ee49d22970f95ada0e17981bd = 
        y_nr_in[28] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[124] = 
I09dd53def80e325c7ea5c3c8e2f064b02ebfe59c3b761e79a215a689b5e7cc40 ^ 
Ic4ee10cf7e9ac1639974ed5497d880be058a326ee49d22970f95ada0e17981bd ^ 
0; 



wire I8a013efc26787c6ce8f85e42c73d78841020ba2c76844a4dae33aeece25c5357;
assign I8a013efc26787c6ce8f85e42c73d78841020ba2c76844a4dae33aeece25c5357 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[38] ^ 
0; 



wire If146f5cbb87aa733d3670aa11cd2d473c0210e93b491076f9b0cb47897cb6de4;
assign If146f5cbb87aa733d3670aa11cd2d473c0210e93b491076f9b0cb47897cb6de4 = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[123] = 
I8a013efc26787c6ce8f85e42c73d78841020ba2c76844a4dae33aeece25c5357 ^ 
If146f5cbb87aa733d3670aa11cd2d473c0210e93b491076f9b0cb47897cb6de4 ^ 
0; 



wire Ie3eb10e9c58d1d3a6b6508f0e4e6f01474249cb13ffb479b1f5413308fb904d5;
assign Ie3eb10e9c58d1d3a6b6508f0e4e6f01474249cb13ffb479b1f5413308fb904d5 = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[39] ^ 
0; 



wire I48a86dd4562ad1ee7cb983fa5ec48fe22a062ac29f56d39e0c2a22c62f35ddd1;
assign I48a86dd4562ad1ee7cb983fa5ec48fe22a062ac29f56d39e0c2a22c62f35ddd1 = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[122] = 
Ie3eb10e9c58d1d3a6b6508f0e4e6f01474249cb13ffb479b1f5413308fb904d5 ^ 
I48a86dd4562ad1ee7cb983fa5ec48fe22a062ac29f56d39e0c2a22c62f35ddd1 ^ 
0; 



wire I198acfe9869520864d1e204df0f6f9c2de50b8e2d495153b89eed1618a9aa245;
assign I198acfe9869520864d1e204df0f6f9c2de50b8e2d495153b89eed1618a9aa245 = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[36] ^ 
0; 



wire I3495bb31e6b02c8c5f2618d5ecfd6abcd4a1245c4eed492511e8901b6bad3fc3;
assign I3495bb31e6b02c8c5f2618d5ecfd6abcd4a1245c4eed492511e8901b6bad3fc3 = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[121] = 
I198acfe9869520864d1e204df0f6f9c2de50b8e2d495153b89eed1618a9aa245 ^ 
I3495bb31e6b02c8c5f2618d5ecfd6abcd4a1245c4eed492511e8901b6bad3fc3 ^ 
0; 



wire I73018bcf124b97c0bc6e72cd6ea93dbfa91414b23010be5b621483f62f3a4578;
assign I73018bcf124b97c0bc6e72cd6ea93dbfa91414b23010be5b621483f62f3a4578 = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[37] ^ 
0; 



wire I9903aa61767059cb2cf1c8df7e5de26f980377650fb9e885ebfe1518e9cca7c2;
assign I9903aa61767059cb2cf1c8df7e5de26f980377650fb9e885ebfe1518e9cca7c2 = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[120] = 
I73018bcf124b97c0bc6e72cd6ea93dbfa91414b23010be5b621483f62f3a4578 ^ 
I9903aa61767059cb2cf1c8df7e5de26f980377650fb9e885ebfe1518e9cca7c2 ^ 
0; 



wire I6f6357d36e2e7908a0040f12e0e72e8fbee173fa530262abf4fd5ca4d98f4668;
assign I6f6357d36e2e7908a0040f12e0e72e8fbee173fa530262abf4fd5ca4d98f4668 = 
        y_nr_in[7] ^ 
        y_nr_in[15] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[119] = 
I6f6357d36e2e7908a0040f12e0e72e8fbee173fa530262abf4fd5ca4d98f4668 ^ 
0; 



wire I0016f92178cc6d08a0bf61e8ace71cb46a555e6d5691390e2e8d68f36cf884f1;
assign I0016f92178cc6d08a0bf61e8ace71cb46a555e6d5691390e2e8d68f36cf884f1 = 
        y_nr_in[4] ^ 
        y_nr_in[12] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[118] = 
I0016f92178cc6d08a0bf61e8ace71cb46a555e6d5691390e2e8d68f36cf884f1 ^ 
0; 



wire I828edcf234bef402fe2316bb47470ed601da0d7c8873c5a08924ed7d7b8acc13;
assign I828edcf234bef402fe2316bb47470ed601da0d7c8873c5a08924ed7d7b8acc13 = 
        y_nr_in[5] ^ 
        y_nr_in[13] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[117] = 
I828edcf234bef402fe2316bb47470ed601da0d7c8873c5a08924ed7d7b8acc13 ^ 
0; 



wire If9954bea361542b75caef106626c8c70a82af99e72e42bb3ef82bcdce6812c14;
assign If9954bea361542b75caef106626c8c70a82af99e72e42bb3ef82bcdce6812c14 = 
        y_nr_in[6] ^ 
        y_nr_in[14] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[116] = 
If9954bea361542b75caef106626c8c70a82af99e72e42bb3ef82bcdce6812c14 ^ 
0; 



wire I0e74277dc013daff01c991b662f603636c49561ddcdcce2a615c6e436223375e;
assign I0e74277dc013daff01c991b662f603636c49561ddcdcce2a615c6e436223375e = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[34] ^ 
0; 



wire Ic970d99e98ba5644a886ece2cddf97502187fec5ec54399b862f39a4a2df007a;
assign Ic970d99e98ba5644a886ece2cddf97502187fec5ec54399b862f39a4a2df007a = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[115] = 
I0e74277dc013daff01c991b662f603636c49561ddcdcce2a615c6e436223375e ^ 
Ic970d99e98ba5644a886ece2cddf97502187fec5ec54399b862f39a4a2df007a ^ 
0; 



wire I8270680f0bdef107e425e370941e7551c61b94445426e1d05ae82ebccd640a31;
assign I8270680f0bdef107e425e370941e7551c61b94445426e1d05ae82ebccd640a31 = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[35] ^ 
0; 



wire I0fde1f6cd5768c0db88db6fe4787f0666b60526f54dbb03b20e7140016de2d6d;
assign I0fde1f6cd5768c0db88db6fe4787f0666b60526f54dbb03b20e7140016de2d6d = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[114] = 
I8270680f0bdef107e425e370941e7551c61b94445426e1d05ae82ebccd640a31 ^ 
I0fde1f6cd5768c0db88db6fe4787f0666b60526f54dbb03b20e7140016de2d6d ^ 
0; 



wire If4b9e7140e7d54fc9a5edf7419466cc3b1ffafae193e57955ab6ba0126935612;
assign If4b9e7140e7d54fc9a5edf7419466cc3b1ffafae193e57955ab6ba0126935612 = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[32] ^ 
0; 



wire Iafc7a22c3b9522c120eab1986d620ab111ef19085a4d93c555cb29508320258a;
assign Iafc7a22c3b9522c120eab1986d620ab111ef19085a4d93c555cb29508320258a = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[113] = 
If4b9e7140e7d54fc9a5edf7419466cc3b1ffafae193e57955ab6ba0126935612 ^ 
Iafc7a22c3b9522c120eab1986d620ab111ef19085a4d93c555cb29508320258a ^ 
0; 



wire I11a3fb05b63d83c01200575b62acae3aadc314ce9aab3cfc712ad953e8c6be0d;
assign I11a3fb05b63d83c01200575b62acae3aadc314ce9aab3cfc712ad953e8c6be0d = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[33] ^ 
0; 



wire I661dbdae6a06dfb663e0eab81a4eeea0bf32d10fddee29ca17dfc8892fa0c1fd;
assign I661dbdae6a06dfb663e0eab81a4eeea0bf32d10fddee29ca17dfc8892fa0c1fd = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[112] = 
I11a3fb05b63d83c01200575b62acae3aadc314ce9aab3cfc712ad953e8c6be0d ^ 
I661dbdae6a06dfb663e0eab81a4eeea0bf32d10fddee29ca17dfc8892fa0c1fd ^ 
0; 



wire Idf28e7e65f6083f41b0e07b8e973799209c760d5847f4455789ca23d090e95a4;
assign Idf28e7e65f6083f41b0e07b8e973799209c760d5847f4455789ca23d090e95a4 = 
        y_nr_in[7] ^ 
        y_nr_in[25] ^ 
        y_nr_in[47] ^ 
0; 



wire If137b1c6ddff5cbc91b835e9e6a58bf730fe508bf743278acc77bcfc08055740;
assign If137b1c6ddff5cbc91b835e9e6a58bf730fe508bf743278acc77bcfc08055740 = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[111] = 
Idf28e7e65f6083f41b0e07b8e973799209c760d5847f4455789ca23d090e95a4 ^ 
If137b1c6ddff5cbc91b835e9e6a58bf730fe508bf743278acc77bcfc08055740 ^ 
0; 



wire I568ed6b5eb066fb08f700df101440b08ab685ae80d50bbe9001d0631786bb568;
assign I568ed6b5eb066fb08f700df101440b08ab685ae80d50bbe9001d0631786bb568 = 
        y_nr_in[4] ^ 
        y_nr_in[26] ^ 
        y_nr_in[44] ^ 
0; 



wire I6526732e56e3f5dcd1535b6ecb28529241fe7a4f5edfc8e98552d7809b71a2f3;
assign I6526732e56e3f5dcd1535b6ecb28529241fe7a4f5edfc8e98552d7809b71a2f3 = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[110] = 
I568ed6b5eb066fb08f700df101440b08ab685ae80d50bbe9001d0631786bb568 ^ 
I6526732e56e3f5dcd1535b6ecb28529241fe7a4f5edfc8e98552d7809b71a2f3 ^ 
0; 



wire I0e482967ea7d57374d6f59e40de6353c393a3d4a2a00d2ba78e8771b2fc70c49;
assign I0e482967ea7d57374d6f59e40de6353c393a3d4a2a00d2ba78e8771b2fc70c49 = 
        y_nr_in[5] ^ 
        y_nr_in[27] ^ 
        y_nr_in[45] ^ 
0; 



wire I1d2c7f473b80536c78739cb61fe4b82f212f19bf96e30a8c767456f7395e5b57;
assign I1d2c7f473b80536c78739cb61fe4b82f212f19bf96e30a8c767456f7395e5b57 = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[109] = 
I0e482967ea7d57374d6f59e40de6353c393a3d4a2a00d2ba78e8771b2fc70c49 ^ 
I1d2c7f473b80536c78739cb61fe4b82f212f19bf96e30a8c767456f7395e5b57 ^ 
0; 



wire Icdf9ac94d836cad93dfa839c9a62b7e868031f7668df7c94ef1697e802dcc877;
assign Icdf9ac94d836cad93dfa839c9a62b7e868031f7668df7c94ef1697e802dcc877 = 
        y_nr_in[6] ^ 
        y_nr_in[24] ^ 
        y_nr_in[46] ^ 
0; 



wire I61fd8679995a76dfae8612070cc2f5076c5f927d6a74c74e20594c0204e582a8;
assign I61fd8679995a76dfae8612070cc2f5076c5f927d6a74c74e20594c0204e582a8 = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[108] = 
Icdf9ac94d836cad93dfa839c9a62b7e868031f7668df7c94ef1697e802dcc877 ^ 
I61fd8679995a76dfae8612070cc2f5076c5f927d6a74c74e20594c0204e582a8 ^ 
0; 



wire I460fa50de867246cdbafbb2ed7c1ecd55ded8d3aedcfdb817d6ccf8db5871d23;
assign I460fa50de867246cdbafbb2ed7c1ecd55ded8d3aedcfdb817d6ccf8db5871d23 = 
        y_nr_in[3] ^ 
        y_nr_in[43] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[107] = 
I460fa50de867246cdbafbb2ed7c1ecd55ded8d3aedcfdb817d6ccf8db5871d23 ^ 
0; 



wire I9b1e08a0ca00dc7e8f7daf895fda5497cbe70eaa656ac4ff277551e97018fefb;
assign I9b1e08a0ca00dc7e8f7daf895fda5497cbe70eaa656ac4ff277551e97018fefb = 
        y_nr_in[0] ^ 
        y_nr_in[40] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[106] = 
I9b1e08a0ca00dc7e8f7daf895fda5497cbe70eaa656ac4ff277551e97018fefb ^ 
0; 



wire Ibbe4b59beb321340409af03246b06a8e9a4d456aa02b0997ebc46f152fa802a8;
assign Ibbe4b59beb321340409af03246b06a8e9a4d456aa02b0997ebc46f152fa802a8 = 
        y_nr_in[1] ^ 
        y_nr_in[41] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[105] = 
Ibbe4b59beb321340409af03246b06a8e9a4d456aa02b0997ebc46f152fa802a8 ^ 
0; 



wire Ibc45c4ef0bbb3d113baea1e18c7f8d3f6f96e321f2ab4ebe81f846bf69777242;
assign Ibc45c4ef0bbb3d113baea1e18c7f8d3f6f96e321f2ab4ebe81f846bf69777242 = 
        y_nr_in[2] ^ 
        y_nr_in[42] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[104] = 
Ibc45c4ef0bbb3d113baea1e18c7f8d3f6f96e321f2ab4ebe81f846bf69777242 ^ 
0; 



wire Ie0f8f4f7109da8084b2b8eca4bc4215906cfc7e6edd880b1aa29939559202701;
assign Ie0f8f4f7109da8084b2b8eca4bc4215906cfc7e6edd880b1aa29939559202701 = 
        y_nr_in[7] ^ 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
0; 



wire I4a034e140ff6704507718dc662e31d17937378bf7f4fcf2e3c7c5893e82f1446;
assign I4a034e140ff6704507718dc662e31d17937378bf7f4fcf2e3c7c5893e82f1446 = 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[103] = 
Ie0f8f4f7109da8084b2b8eca4bc4215906cfc7e6edd880b1aa29939559202701 ^ 
I4a034e140ff6704507718dc662e31d17937378bf7f4fcf2e3c7c5893e82f1446 ^ 
0; 



wire I57c8dc6535a07e9500c1d69fb47ae667fe2f17d2582a74d8353a783a62c45a8a;
assign I57c8dc6535a07e9500c1d69fb47ae667fe2f17d2582a74d8353a783a62c45a8a = 
        y_nr_in[4] ^ 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
0; 



wire I04638b9702944c928ffa6af39c16d2b2459bafb08c217632829160b6e59bf366;
assign I04638b9702944c928ffa6af39c16d2b2459bafb08c217632829160b6e59bf366 = 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[102] = 
I57c8dc6535a07e9500c1d69fb47ae667fe2f17d2582a74d8353a783a62c45a8a ^ 
I04638b9702944c928ffa6af39c16d2b2459bafb08c217632829160b6e59bf366 ^ 
0; 



wire Ide2a61371c25d75c6fe8b6f961d9d61ffa5a571c624df6eca6606b9ec20d1bba;
assign Ide2a61371c25d75c6fe8b6f961d9d61ffa5a571c624df6eca6606b9ec20d1bba = 
        y_nr_in[5] ^ 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
0; 



wire Idbfb2cc978510c1c9dcf503b4116b3df6f85be5bdb63340fe67fb22281e4c3d5;
assign Idbfb2cc978510c1c9dcf503b4116b3df6f85be5bdb63340fe67fb22281e4c3d5 = 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[101] = 
Ide2a61371c25d75c6fe8b6f961d9d61ffa5a571c624df6eca6606b9ec20d1bba ^ 
Idbfb2cc978510c1c9dcf503b4116b3df6f85be5bdb63340fe67fb22281e4c3d5 ^ 
0; 



wire Ice55a85f2415b4c7279ede14afed095c630a5bc515e04d114b4b0d51cd3799d6;
assign Ice55a85f2415b4c7279ede14afed095c630a5bc515e04d114b4b0d51cd3799d6 = 
        y_nr_in[6] ^ 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
0; 



wire Ic528b972a32ef56e743cd2588508ea3ce39cb9a3eb1ac6ff5290b9eb3db01728;
assign Ic528b972a32ef56e743cd2588508ea3ce39cb9a3eb1ac6ff5290b9eb3db01728 = 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[100] = 
Ice55a85f2415b4c7279ede14afed095c630a5bc515e04d114b4b0d51cd3799d6 ^ 
Ic528b972a32ef56e743cd2588508ea3ce39cb9a3eb1ac6ff5290b9eb3db01728 ^ 
0; 



wire Ic815e6831394d6bd3233a3e4459d1bf98d212c4e76047397ea19d092b25e36df;
assign Ic815e6831394d6bd3233a3e4459d1bf98d212c4e76047397ea19d092b25e36df = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[46] ^ 
0; 



wire I187ae6c92c5db73f13c20c8c99a5d179a56b9cb61b478de1310032a0fd4ff666;
assign I187ae6c92c5db73f13c20c8c99a5d179a56b9cb61b478de1310032a0fd4ff666 = 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[99] = 
Ic815e6831394d6bd3233a3e4459d1bf98d212c4e76047397ea19d092b25e36df ^ 
I187ae6c92c5db73f13c20c8c99a5d179a56b9cb61b478de1310032a0fd4ff666 ^ 
0; 



wire I6a680c4155beebef7694e7ee0792fae3bda79332e666cf11255339a2c8d7058b;
assign I6a680c4155beebef7694e7ee0792fae3bda79332e666cf11255339a2c8d7058b = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[47] ^ 
0; 



wire Ib069571649c5c887e2cbd7a4d0338ab559f7c4dd886046a2d09167a46334c555;
assign Ib069571649c5c887e2cbd7a4d0338ab559f7c4dd886046a2d09167a46334c555 = 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[98] = 
I6a680c4155beebef7694e7ee0792fae3bda79332e666cf11255339a2c8d7058b ^ 
Ib069571649c5c887e2cbd7a4d0338ab559f7c4dd886046a2d09167a46334c555 ^ 
0; 



wire I6e417d3a471a9e0d9f5d49dea659fcf95546c65bf8a89b4ff8236b99e60f164f;
assign I6e417d3a471a9e0d9f5d49dea659fcf95546c65bf8a89b4ff8236b99e60f164f = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[44] ^ 
0; 



wire I491c60a528bfdd4cb94bf33383eeef5c85a5278bac31ed0f7b506350ac7f36f9;
assign I491c60a528bfdd4cb94bf33383eeef5c85a5278bac31ed0f7b506350ac7f36f9 = 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[97] = 
I6e417d3a471a9e0d9f5d49dea659fcf95546c65bf8a89b4ff8236b99e60f164f ^ 
I491c60a528bfdd4cb94bf33383eeef5c85a5278bac31ed0f7b506350ac7f36f9 ^ 
0; 



wire I91641d702f8e03b4ac11a95d171c335003dc9432f89e8c5b2de0b1a15af20f83;
assign I91641d702f8e03b4ac11a95d171c335003dc9432f89e8c5b2de0b1a15af20f83 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[45] ^ 
0; 



wire Ifc3aef378b28c216a4af8fb5f7dcdf89cf548b2e36f0bf0c77ad0b11d82eddce;
assign Ifc3aef378b28c216a4af8fb5f7dcdf89cf548b2e36f0bf0c77ad0b11d82eddce = 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[96] = 
I91641d702f8e03b4ac11a95d171c335003dc9432f89e8c5b2de0b1a15af20f83 ^ 
Ifc3aef378b28c216a4af8fb5f7dcdf89cf548b2e36f0bf0c77ad0b11d82eddce ^ 
0; 



wire Ie2b96c7554f57d93f81837f59c7f9a2c8f6cb907e2338b0c70294da7d0127afb;
assign Ie2b96c7554f57d93f81837f59c7f9a2c8f6cb907e2338b0c70294da7d0127afb = 
        y_nr_in[0] ^ 
        y_nr_in[26] ^ 
        y_nr_in[30] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[95] = 
Ie2b96c7554f57d93f81837f59c7f9a2c8f6cb907e2338b0c70294da7d0127afb ^ 
0; 



wire I17884245955f22f700a4465acc6df8ea9a629629dbfa7317da5b1639d55d1328;
assign I17884245955f22f700a4465acc6df8ea9a629629dbfa7317da5b1639d55d1328 = 
        y_nr_in[1] ^ 
        y_nr_in[27] ^ 
        y_nr_in[31] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[94] = 
I17884245955f22f700a4465acc6df8ea9a629629dbfa7317da5b1639d55d1328 ^ 
0; 



wire I856ef2bb3dc89e261fcfd023d50ce1779036a51c8abccb8eff03feadeb2136c1;
assign I856ef2bb3dc89e261fcfd023d50ce1779036a51c8abccb8eff03feadeb2136c1 = 
        y_nr_in[2] ^ 
        y_nr_in[24] ^ 
        y_nr_in[28] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[93] = 
I856ef2bb3dc89e261fcfd023d50ce1779036a51c8abccb8eff03feadeb2136c1 ^ 
0; 



wire Ic3a6500f0db687d0d51af6fbdb08f18912f269e77726fdfa48dd416825b289f9;
assign Ic3a6500f0db687d0d51af6fbdb08f18912f269e77726fdfa48dd416825b289f9 = 
        y_nr_in[3] ^ 
        y_nr_in[25] ^ 
        y_nr_in[29] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[92] = 
Ic3a6500f0db687d0d51af6fbdb08f18912f269e77726fdfa48dd416825b289f9 ^ 
0; 



wire Ib27dc99958ae9b7eb461d6d0c638490563f842df99914da2d3b080bdd6ca8cf4;
assign Ib27dc99958ae9b7eb461d6d0c638490563f842df99914da2d3b080bdd6ca8cf4 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[41] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[91] = 
Ib27dc99958ae9b7eb461d6d0c638490563f842df99914da2d3b080bdd6ca8cf4 ^ 
0; 



wire Ia864fdd01430b3da092a9470cf806a86a8c8a8af5ea75238dde57eb4dc0152dc;
assign Ia864fdd01430b3da092a9470cf806a86a8c8a8af5ea75238dde57eb4dc0152dc = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[42] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[90] = 
Ia864fdd01430b3da092a9470cf806a86a8c8a8af5ea75238dde57eb4dc0152dc ^ 
0; 



wire If40b9c212bd0e0de6f44f266a1bdc600f3aacc50aa5bde4a4d88f3edd1bf545c;
assign If40b9c212bd0e0de6f44f266a1bdc600f3aacc50aa5bde4a4d88f3edd1bf545c = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[43] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[89] = 
If40b9c212bd0e0de6f44f266a1bdc600f3aacc50aa5bde4a4d88f3edd1bf545c ^ 
0; 



wire Icd8eb0102066b27b8a486a88894c9df50f922063098ef993825f3ac1b4924686;
assign Icd8eb0102066b27b8a486a88894c9df50f922063098ef993825f3ac1b4924686 = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[40] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[88] = 
Icd8eb0102066b27b8a486a88894c9df50f922063098ef993825f3ac1b4924686 ^ 
0; 



wire I3493fe8f496c669528edad1b2638d9849cd91fe9aaad26300f8fed57aa5af16b;
assign I3493fe8f496c669528edad1b2638d9849cd91fe9aaad26300f8fed57aa5af16b = 
        y_nr_in[6] ^ 
        y_nr_in[17] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[87] = 
I3493fe8f496c669528edad1b2638d9849cd91fe9aaad26300f8fed57aa5af16b ^ 
0; 



wire Iee6d3f0d039c72da19a800305f1b5ae80057a2366ab53fb37bcbbf6fe541da47;
assign Iee6d3f0d039c72da19a800305f1b5ae80057a2366ab53fb37bcbbf6fe541da47 = 
        y_nr_in[7] ^ 
        y_nr_in[18] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[86] = 
Iee6d3f0d039c72da19a800305f1b5ae80057a2366ab53fb37bcbbf6fe541da47 ^ 
0; 



wire Ie287803eacbc0f4a71a1a0ac982c3ee7fa386e67f8660465bb0753e8222a6eb0;
assign Ie287803eacbc0f4a71a1a0ac982c3ee7fa386e67f8660465bb0753e8222a6eb0 = 
        y_nr_in[4] ^ 
        y_nr_in[19] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[85] = 
Ie287803eacbc0f4a71a1a0ac982c3ee7fa386e67f8660465bb0753e8222a6eb0 ^ 
0; 



wire I47715d5589693a211add4325635d4f400f10ff3764c88053c43945b8987786a0;
assign I47715d5589693a211add4325635d4f400f10ff3764c88053c43945b8987786a0 = 
        y_nr_in[5] ^ 
        y_nr_in[16] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[84] = 
I47715d5589693a211add4325635d4f400f10ff3764c88053c43945b8987786a0 ^ 
0; 



wire Id67bcba60edfed75aaccd2da1f874ebc0f9f0724c9e4e6eb7de598640c2fd1ee;
assign Id67bcba60edfed75aaccd2da1f874ebc0f9f0724c9e4e6eb7de598640c2fd1ee = 
        y_nr_in[0] ^ 
        y_nr_in[34] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[83] = 
Id67bcba60edfed75aaccd2da1f874ebc0f9f0724c9e4e6eb7de598640c2fd1ee ^ 
0; 



wire I8508ddaab52430f316f9f16f378014ffc6a953fc4c4925dc22b3f01fab1e04ec;
assign I8508ddaab52430f316f9f16f378014ffc6a953fc4c4925dc22b3f01fab1e04ec = 
        y_nr_in[1] ^ 
        y_nr_in[35] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[82] = 
I8508ddaab52430f316f9f16f378014ffc6a953fc4c4925dc22b3f01fab1e04ec ^ 
0; 



wire I3588f0f60c6328afd0bfe1581a303b8f31e2ae540c44f66b3d384abaa24adfa1;
assign I3588f0f60c6328afd0bfe1581a303b8f31e2ae540c44f66b3d384abaa24adfa1 = 
        y_nr_in[2] ^ 
        y_nr_in[32] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[81] = 
I3588f0f60c6328afd0bfe1581a303b8f31e2ae540c44f66b3d384abaa24adfa1 ^ 
0; 



wire Ie24702beb392c5cd6079ed852052c54b3c86e2f10600e0dca3b8da0b62173a37;
assign Ie24702beb392c5cd6079ed852052c54b3c86e2f10600e0dca3b8da0b62173a37 = 
        y_nr_in[3] ^ 
        y_nr_in[33] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[80] = 
Ie24702beb392c5cd6079ed852052c54b3c86e2f10600e0dca3b8da0b62173a37 ^ 
0; 



wire I34b0ed27c72aebdc29f3e3cc6a170d2b86346de7b312ffebc3590537e8c36dda;
assign I34b0ed27c72aebdc29f3e3cc6a170d2b86346de7b312ffebc3590537e8c36dda = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[79] = 
I34b0ed27c72aebdc29f3e3cc6a170d2b86346de7b312ffebc3590537e8c36dda ^ 
0; 



wire I6eb66d4ad80b754c798d8c65f508f306cb534e3e6f249c4b0fa2ee249edd48b4;
assign I6eb66d4ad80b754c798d8c65f508f306cb534e3e6f249c4b0fa2ee249edd48b4 = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[78] = 
I6eb66d4ad80b754c798d8c65f508f306cb534e3e6f249c4b0fa2ee249edd48b4 ^ 
0; 



wire I4c5fd7f7ce5884fa78166d52d40761ae321ea77b9af18883e25457e5b8669979;
assign I4c5fd7f7ce5884fa78166d52d40761ae321ea77b9af18883e25457e5b8669979 = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[77] = 
I4c5fd7f7ce5884fa78166d52d40761ae321ea77b9af18883e25457e5b8669979 ^ 
0; 



wire I749df42857ecb08093aee2c6644a8d7ae85aacfbdd2223f385356c9c6d9debf2;
assign I749df42857ecb08093aee2c6644a8d7ae85aacfbdd2223f385356c9c6d9debf2 = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[76] = 
I749df42857ecb08093aee2c6644a8d7ae85aacfbdd2223f385356c9c6d9debf2 ^ 
0; 



wire I53dc58bcb983b221b7a34972e449bc96837c8331da3c4766e2b8f7dadfbe1df5;
assign I53dc58bcb983b221b7a34972e449bc96837c8331da3c4766e2b8f7dadfbe1df5 = 
        y_nr_in[3] ^ 
        y_nr_in[15] ^ 
        y_nr_in[22] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[75] = 
I53dc58bcb983b221b7a34972e449bc96837c8331da3c4766e2b8f7dadfbe1df5 ^ 
0; 



wire I713925d1fb7388f25956294817f33209972f03f18c8aacec62e323d73ce4d899;
assign I713925d1fb7388f25956294817f33209972f03f18c8aacec62e323d73ce4d899 = 
        y_nr_in[0] ^ 
        y_nr_in[12] ^ 
        y_nr_in[23] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[74] = 
I713925d1fb7388f25956294817f33209972f03f18c8aacec62e323d73ce4d899 ^ 
0; 



wire Id591d53cae95d78d56e6790d8d48fdb1fccd924a3d74702da7da5906959360e3;
assign Id591d53cae95d78d56e6790d8d48fdb1fccd924a3d74702da7da5906959360e3 = 
        y_nr_in[1] ^ 
        y_nr_in[13] ^ 
        y_nr_in[20] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[73] = 
Id591d53cae95d78d56e6790d8d48fdb1fccd924a3d74702da7da5906959360e3 ^ 
0; 



wire I73435e48db187904fd803883a02dbb1dd75475a4acafef77a92b97309c741547;
assign I73435e48db187904fd803883a02dbb1dd75475a4acafef77a92b97309c741547 = 
        y_nr_in[2] ^ 
        y_nr_in[14] ^ 
        y_nr_in[21] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[72] = 
I73435e48db187904fd803883a02dbb1dd75475a4acafef77a92b97309c741547 ^ 
0; 



wire I49252a481f98d44f48d620df37f7d2d75e8a81d0cfab91bb4eb7916b02e723f1;
assign I49252a481f98d44f48d620df37f7d2d75e8a81d0cfab91bb4eb7916b02e723f1 = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
        y_nr_in[36] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[71] = 
I49252a481f98d44f48d620df37f7d2d75e8a81d0cfab91bb4eb7916b02e723f1 ^ 
0; 



wire I5080b7960640e21fb77dc33352d27bf9decc8acbed5287cfa78f7c86f5185b67;
assign I5080b7960640e21fb77dc33352d27bf9decc8acbed5287cfa78f7c86f5185b67 = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
        y_nr_in[37] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[70] = 
I5080b7960640e21fb77dc33352d27bf9decc8acbed5287cfa78f7c86f5185b67 ^ 
0; 



wire I517f12ae677e7d31fe721b16e3d659791b88c96a49f102fc4f8f784fab4e16cf;
assign I517f12ae677e7d31fe721b16e3d659791b88c96a49f102fc4f8f784fab4e16cf = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
        y_nr_in[38] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[69] = 
I517f12ae677e7d31fe721b16e3d659791b88c96a49f102fc4f8f784fab4e16cf ^ 
0; 



wire I8af4fe02e31ae2c79e572080447a2006f2c54deee1e3f370e18aa76d8e6e8009;
assign I8af4fe02e31ae2c79e572080447a2006f2c54deee1e3f370e18aa76d8e6e8009 = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
        y_nr_in[39] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[68] = 
I8af4fe02e31ae2c79e572080447a2006f2c54deee1e3f370e18aa76d8e6e8009 ^ 
0; 



wire I1ab665c6065ef3648ba7c3f60490950063786ffa51ecfe072b7b742287e40e08;
assign I1ab665c6065ef3648ba7c3f60490950063786ffa51ecfe072b7b742287e40e08 = 
        y_nr_in[0] ^ 
        y_nr_in[20] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[67] = 
I1ab665c6065ef3648ba7c3f60490950063786ffa51ecfe072b7b742287e40e08 ^ 
0; 



wire I596474d97feb75010bbe35074c3d27ab53abab03c5f847dde9ed7e12c18a06b3;
assign I596474d97feb75010bbe35074c3d27ab53abab03c5f847dde9ed7e12c18a06b3 = 
        y_nr_in[1] ^ 
        y_nr_in[21] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[66] = 
I596474d97feb75010bbe35074c3d27ab53abab03c5f847dde9ed7e12c18a06b3 ^ 
0; 



wire Ib8ca8cb082f23a8576f5be9d860e817e4b4b743a50e7acb71d670fd34eb3a757;
assign Ib8ca8cb082f23a8576f5be9d860e817e4b4b743a50e7acb71d670fd34eb3a757 = 
        y_nr_in[2] ^ 
        y_nr_in[22] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[65] = 
Ib8ca8cb082f23a8576f5be9d860e817e4b4b743a50e7acb71d670fd34eb3a757 ^ 
0; 



wire I36f163a586d548d9b2289c99f0ee152ce6af33124f04fdc15b7934eb27e80e57;
assign I36f163a586d548d9b2289c99f0ee152ce6af33124f04fdc15b7934eb27e80e57 = 
        y_nr_in[3] ^ 
        y_nr_in[23] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[64] = 
I36f163a586d548d9b2289c99f0ee152ce6af33124f04fdc15b7934eb27e80e57 ^ 
0; 



wire Ie80a6a85ea5a89ff4d07c8d0f73db32f967fae4ce8c4d7d08a0588ea9f1f8690;
assign Ie80a6a85ea5a89ff4d07c8d0f73db32f967fae4ce8c4d7d08a0588ea9f1f8690 = 
        y_nr_in[9] ^ 
        y_nr_in[31] ^ 
        y_nr_in[48] ^ 
0; 



wire I2ba5ef033b7b82351761dff13dfefd872c97b8685a5d1bc784b4bf02d6c87d39;
assign I2ba5ef033b7b82351761dff13dfefd872c97b8685a5d1bc784b4bf02d6c87d39 = 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[63] = 
Ie80a6a85ea5a89ff4d07c8d0f73db32f967fae4ce8c4d7d08a0588ea9f1f8690 ^ 
I2ba5ef033b7b82351761dff13dfefd872c97b8685a5d1bc784b4bf02d6c87d39 ^ 
0; 



wire Icbbd64503e6a0d82ec8627bebd70e7b3d0781e378b46fe8deefc4aae0f552c1c;
assign Icbbd64503e6a0d82ec8627bebd70e7b3d0781e378b46fe8deefc4aae0f552c1c = 
        y_nr_in[10] ^ 
        y_nr_in[28] ^ 
        y_nr_in[49] ^ 
0; 



wire I286072f35d8290d6c8e9e3def951d8acd165dee25d8e779a61db19f19f669b1d;
assign I286072f35d8290d6c8e9e3def951d8acd165dee25d8e779a61db19f19f669b1d = 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[62] = 
Icbbd64503e6a0d82ec8627bebd70e7b3d0781e378b46fe8deefc4aae0f552c1c ^ 
I286072f35d8290d6c8e9e3def951d8acd165dee25d8e779a61db19f19f669b1d ^ 
0; 



wire I53fbf7ceacac2cb4382d381d1397bf17070108bbca2a2a7f6c5c74ea262c0efd;
assign I53fbf7ceacac2cb4382d381d1397bf17070108bbca2a2a7f6c5c74ea262c0efd = 
        y_nr_in[11] ^ 
        y_nr_in[29] ^ 
        y_nr_in[50] ^ 
0; 



wire Iee963cac29e88334eec5d027674ef03159de83d4deed1fde3debd840e986cdb2;
assign Iee963cac29e88334eec5d027674ef03159de83d4deed1fde3debd840e986cdb2 = 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[61] = 
I53fbf7ceacac2cb4382d381d1397bf17070108bbca2a2a7f6c5c74ea262c0efd ^ 
Iee963cac29e88334eec5d027674ef03159de83d4deed1fde3debd840e986cdb2 ^ 
0; 



wire I57ae842a4001d14a9ead5fbdda7ed281087e3d9c6a838e9f23d583e7b9580d3e;
assign I57ae842a4001d14a9ead5fbdda7ed281087e3d9c6a838e9f23d583e7b9580d3e = 
        y_nr_in[8] ^ 
        y_nr_in[30] ^ 
        y_nr_in[51] ^ 
0; 



wire I2372eae8be20255d9196b8eaca424420614b1fcb506174c9dbaf33d47fcc0584;
assign I2372eae8be20255d9196b8eaca424420614b1fcb506174c9dbaf33d47fcc0584 = 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[60] = 
I57ae842a4001d14a9ead5fbdda7ed281087e3d9c6a838e9f23d583e7b9580d3e ^ 
I2372eae8be20255d9196b8eaca424420614b1fcb506174c9dbaf33d47fcc0584 ^ 
0; 



wire Ie77f954a2c57942bfa06d607d78ea178a615bf38c160431bff53683987a1fed5;
assign Ie77f954a2c57942bfa06d607d78ea178a615bf38c160431bff53683987a1fed5 = 
        y_nr_in[0] ^ 
        y_nr_in[27] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[59] = 
Ie77f954a2c57942bfa06d607d78ea178a615bf38c160431bff53683987a1fed5 ^ 
0; 



wire Ie963a8840cb2771f615bd29bc69d572a2992b1ae6391979fff65625d8a31cc8f;
assign Ie963a8840cb2771f615bd29bc69d572a2992b1ae6391979fff65625d8a31cc8f = 
        y_nr_in[1] ^ 
        y_nr_in[24] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[58] = 
Ie963a8840cb2771f615bd29bc69d572a2992b1ae6391979fff65625d8a31cc8f ^ 
0; 



wire I615148ffa13066e02286c8fe3cb5e02104938f716f63286ea03a31309b5ef87d;
assign I615148ffa13066e02286c8fe3cb5e02104938f716f63286ea03a31309b5ef87d = 
        y_nr_in[2] ^ 
        y_nr_in[25] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[57] = 
I615148ffa13066e02286c8fe3cb5e02104938f716f63286ea03a31309b5ef87d ^ 
0; 



wire Ia89469f2c045394fd67fc5894edf5a18e01cec8b06d2330030b2650a1ac75095;
assign Ia89469f2c045394fd67fc5894edf5a18e01cec8b06d2330030b2650a1ac75095 = 
        y_nr_in[3] ^ 
        y_nr_in[26] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[56] = 
Ia89469f2c045394fd67fc5894edf5a18e01cec8b06d2330030b2650a1ac75095 ^ 
0; 



wire Ib6f4d9266a6f14fc6caf20815aa51585d46b9bb64cbc3583614a9f47a04aedc5;
assign Ib6f4d9266a6f14fc6caf20815aa51585d46b9bb64cbc3583614a9f47a04aedc5 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[23] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[55] = 
Ib6f4d9266a6f14fc6caf20815aa51585d46b9bb64cbc3583614a9f47a04aedc5 ^ 
0; 



wire I3e60785d78abce1e17afa451061f2c16cf218fde5959c5b8c3773cdfefb00357;
assign I3e60785d78abce1e17afa451061f2c16cf218fde5959c5b8c3773cdfefb00357 = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[20] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[54] = 
I3e60785d78abce1e17afa451061f2c16cf218fde5959c5b8c3773cdfefb00357 ^ 
0; 



wire I85e3a5446ecf87fa69161582b8d2570fffbf6166b18f3e3fb7dab2b3934173c6;
assign I85e3a5446ecf87fa69161582b8d2570fffbf6166b18f3e3fb7dab2b3934173c6 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[21] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[53] = 
I85e3a5446ecf87fa69161582b8d2570fffbf6166b18f3e3fb7dab2b3934173c6 ^ 
0; 



wire Ifbe4a51ca6a0ff79d51706849ccac91d91013bf1d4c10860f9c09fec7d7acaf8;
assign Ifbe4a51ca6a0ff79d51706849ccac91d91013bf1d4c10860f9c09fec7d7acaf8 = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[22] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[52] = 
Ifbe4a51ca6a0ff79d51706849ccac91d91013bf1d4c10860f9c09fec7d7acaf8 ^ 
0; 



wire Iaa7fcac337b655b01c8c08546d9e383ead46575b522ed4a4355628ba67ca4fb1;
assign Iaa7fcac337b655b01c8c08546d9e383ead46575b522ed4a4355628ba67ca4fb1 = 
        y_nr_in[2] ^ 
        y_nr_in[16] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[51] = 
Iaa7fcac337b655b01c8c08546d9e383ead46575b522ed4a4355628ba67ca4fb1 ^ 
0; 



wire Ibdf7ebe201cc10bc9e3809cf2240498e771574655b7f896bbfad6ee92aca8a23;
assign Ibdf7ebe201cc10bc9e3809cf2240498e771574655b7f896bbfad6ee92aca8a23 = 
        y_nr_in[3] ^ 
        y_nr_in[17] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[50] = 
Ibdf7ebe201cc10bc9e3809cf2240498e771574655b7f896bbfad6ee92aca8a23 ^ 
0; 



wire Ib60fade8c09d8680a36e5bf1a0284b796673a17e94a819251f2a71e15295fa3b;
assign Ib60fade8c09d8680a36e5bf1a0284b796673a17e94a819251f2a71e15295fa3b = 
        y_nr_in[0] ^ 
        y_nr_in[18] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[49] = 
Ib60fade8c09d8680a36e5bf1a0284b796673a17e94a819251f2a71e15295fa3b ^ 
0; 



wire I68ab23a12dceb8cda9709ed2a8e2988caa47f0fc29e1ff33f3b8940e4d5116ad;
assign I68ab23a12dceb8cda9709ed2a8e2988caa47f0fc29e1ff33f3b8940e4d5116ad = 
        y_nr_in[1] ^ 
        y_nr_in[19] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[48] = 
I68ab23a12dceb8cda9709ed2a8e2988caa47f0fc29e1ff33f3b8940e4d5116ad ^ 
0; 



wire I858df6bb38a70d9caf8b447cfe0dfbb9cb9bd24e9f42adc59d561e8e7425ef35;
assign I858df6bb38a70d9caf8b447cfe0dfbb9cb9bd24e9f42adc59d561e8e7425ef35 = 
        y_nr_in[11] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
0; 



wire I3cbddc8bfb69bb229bbc8084504f4d2d9b07f3cdfa924d0cce6b3c57a8ad8307;
assign I3cbddc8bfb69bb229bbc8084504f4d2d9b07f3cdfa924d0cce6b3c57a8ad8307 = 
        y_nr_in[36] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[47] = 
I858df6bb38a70d9caf8b447cfe0dfbb9cb9bd24e9f42adc59d561e8e7425ef35 ^ 
I3cbddc8bfb69bb229bbc8084504f4d2d9b07f3cdfa924d0cce6b3c57a8ad8307 ^ 
0; 



wire I89d0a135e12a1d3e58ab85368e7b060daafc1fc9debfd29b3faffb2b94fcc86f;
assign I89d0a135e12a1d3e58ab85368e7b060daafc1fc9debfd29b3faffb2b94fcc86f = 
        y_nr_in[8] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
0; 



wire I38239b6ab86f4ff40dff1abeb52aacc9694eba64eebab8322f0d15fca272c9d3;
assign I38239b6ab86f4ff40dff1abeb52aacc9694eba64eebab8322f0d15fca272c9d3 = 
        y_nr_in[37] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[46] = 
I89d0a135e12a1d3e58ab85368e7b060daafc1fc9debfd29b3faffb2b94fcc86f ^ 
I38239b6ab86f4ff40dff1abeb52aacc9694eba64eebab8322f0d15fca272c9d3 ^ 
0; 



wire Idcdd8b778353d44d370a1a3ebac9cda0d67cfe850715e86fdf4aa07c5711a951;
assign Idcdd8b778353d44d370a1a3ebac9cda0d67cfe850715e86fdf4aa07c5711a951 = 
        y_nr_in[9] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
0; 



wire If21d6269cf0a04b6ab675023508e3e7df981656e5426ac641504f414efc97789;
assign If21d6269cf0a04b6ab675023508e3e7df981656e5426ac641504f414efc97789 = 
        y_nr_in[38] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[45] = 
Idcdd8b778353d44d370a1a3ebac9cda0d67cfe850715e86fdf4aa07c5711a951 ^ 
If21d6269cf0a04b6ab675023508e3e7df981656e5426ac641504f414efc97789 ^ 
0; 



wire I4ec3b7ee477264f3d1c336bd00d2fabb40f0116218727e3619709e1296468c24;
assign I4ec3b7ee477264f3d1c336bd00d2fabb40f0116218727e3619709e1296468c24 = 
        y_nr_in[10] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
0; 



wire Ieceddce637e91b17dcdf72e43b0eeacc0af6b3c8983e8863316bf68711130abf;
assign Ieceddce637e91b17dcdf72e43b0eeacc0af6b3c8983e8863316bf68711130abf = 
        y_nr_in[39] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[44] = 
I4ec3b7ee477264f3d1c336bd00d2fabb40f0116218727e3619709e1296468c24 ^ 
Ieceddce637e91b17dcdf72e43b0eeacc0af6b3c8983e8863316bf68711130abf ^ 
0; 



wire I3e6bdfbaa1119c206b79fa1bd1482b00ec49e9faaf6fe9e6cc7a26d0e0cf5601;
assign I3e6bdfbaa1119c206b79fa1bd1482b00ec49e9faaf6fe9e6cc7a26d0e0cf5601 = 
        y_nr_in[6] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[43] = 
I3e6bdfbaa1119c206b79fa1bd1482b00ec49e9faaf6fe9e6cc7a26d0e0cf5601 ^ 
0; 



wire I14bcc7037579859fb0b78322d661a77583d6954f553bf1c312da3edfc4aea4d6;
assign I14bcc7037579859fb0b78322d661a77583d6954f553bf1c312da3edfc4aea4d6 = 
        y_nr_in[7] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[42] = 
I14bcc7037579859fb0b78322d661a77583d6954f553bf1c312da3edfc4aea4d6 ^ 
0; 



wire I1021f3960dc6d9dbead5d89ab46837450094ec1eb9995a54c3e035bc39b41e39;
assign I1021f3960dc6d9dbead5d89ab46837450094ec1eb9995a54c3e035bc39b41e39 = 
        y_nr_in[4] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[41] = 
I1021f3960dc6d9dbead5d89ab46837450094ec1eb9995a54c3e035bc39b41e39 ^ 
0; 



wire Iab07a22132333dc82dfd2bb37d146a4afe639be50119ec29071aef525973c414;
assign Iab07a22132333dc82dfd2bb37d146a4afe639be50119ec29071aef525973c414 = 
        y_nr_in[5] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[40] = 
Iab07a22132333dc82dfd2bb37d146a4afe639be50119ec29071aef525973c414 ^ 
0; 



wire I9a163a0141fb02d6e77ac5f98f95023777b1bdd2d0559a470adc41c4ea43577d;
assign I9a163a0141fb02d6e77ac5f98f95023777b1bdd2d0559a470adc41c4ea43577d = 
        y_nr_in[2] ^ 
        y_nr_in[20] ^ 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[39] = 
I9a163a0141fb02d6e77ac5f98f95023777b1bdd2d0559a470adc41c4ea43577d ^ 
0; 



wire I5a26e40c7eb43827255ff5b9e6899fdb0f953bdcb2713357a5e0df42354aaf6e;
assign I5a26e40c7eb43827255ff5b9e6899fdb0f953bdcb2713357a5e0df42354aaf6e = 
        y_nr_in[3] ^ 
        y_nr_in[21] ^ 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[38] = 
I5a26e40c7eb43827255ff5b9e6899fdb0f953bdcb2713357a5e0df42354aaf6e ^ 
0; 



wire I742b31b070d96174d7fa3e07d33c076cd5347558ac9f3748e8e295c62b9b6fb0;
assign I742b31b070d96174d7fa3e07d33c076cd5347558ac9f3748e8e295c62b9b6fb0 = 
        y_nr_in[0] ^ 
        y_nr_in[22] ^ 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[37] = 
I742b31b070d96174d7fa3e07d33c076cd5347558ac9f3748e8e295c62b9b6fb0 ^ 
0; 



wire I98e606527e6f6149476aaaad3058d09610eb3fce443d51b9f2ebb94eb0ba11d5;
assign I98e606527e6f6149476aaaad3058d09610eb3fce443d51b9f2ebb94eb0ba11d5 = 
        y_nr_in[1] ^ 
        y_nr_in[23] ^ 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[36] = 
I98e606527e6f6149476aaaad3058d09610eb3fce443d51b9f2ebb94eb0ba11d5 ^ 
0; 



wire Ifa6534e692c4719ff1d901c55ec571d49386ea8e467c38aa883ce5c083fe15b9;
assign Ifa6534e692c4719ff1d901c55ec571d49386ea8e467c38aa883ce5c083fe15b9 = 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
        y_nr_in[43] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[35] = 
Ifa6534e692c4719ff1d901c55ec571d49386ea8e467c38aa883ce5c083fe15b9 ^ 
0; 



wire I288a1aa23795bdff16b986b76e9a7129302260d57c547777325c08517ca9b20a;
assign I288a1aa23795bdff16b986b76e9a7129302260d57c547777325c08517ca9b20a = 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
        y_nr_in[40] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[34] = 
I288a1aa23795bdff16b986b76e9a7129302260d57c547777325c08517ca9b20a ^ 
0; 



wire I93810ca283430044c536db07dafa7f79a403cf6ff94f64a9c50460ded24a78ba;
assign I93810ca283430044c536db07dafa7f79a403cf6ff94f64a9c50460ded24a78ba = 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
        y_nr_in[41] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[33] = 
I93810ca283430044c536db07dafa7f79a403cf6ff94f64a9c50460ded24a78ba ^ 
0; 



wire I59ec86accc2b7589153960eec73dbd7768784a1f34484477ecea9c2c55c76049;
assign I59ec86accc2b7589153960eec73dbd7768784a1f34484477ecea9c2c55c76049 = 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
        y_nr_in[42] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[32] = 
I59ec86accc2b7589153960eec73dbd7768784a1f34484477ecea9c2c55c76049 ^ 
0; 



wire I195590f14ca7dabcf696e54d5aa57bc7a7575c819baa1806971d28891abe7284;
assign I195590f14ca7dabcf696e54d5aa57bc7a7575c819baa1806971d28891abe7284 = 
        y_nr_in[3] ^ 
        y_nr_in[49] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[31] = 
I195590f14ca7dabcf696e54d5aa57bc7a7575c819baa1806971d28891abe7284 ^ 
0; 



wire I11b5888b933b13672a1467f18527dfa8c32e0e507331d6fcffb9ccd38d4ce95b;
assign I11b5888b933b13672a1467f18527dfa8c32e0e507331d6fcffb9ccd38d4ce95b = 
        y_nr_in[0] ^ 
        y_nr_in[50] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[30] = 
I11b5888b933b13672a1467f18527dfa8c32e0e507331d6fcffb9ccd38d4ce95b ^ 
0; 



wire I9979b410519f8b7156eca8971de2f144c4c0768e53d3274f2ff10fa9c251cee6;
assign I9979b410519f8b7156eca8971de2f144c4c0768e53d3274f2ff10fa9c251cee6 = 
        y_nr_in[1] ^ 
        y_nr_in[51] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[29] = 
I9979b410519f8b7156eca8971de2f144c4c0768e53d3274f2ff10fa9c251cee6 ^ 
0; 



wire I6d4d8c9c5618d829ae0018df43f15d076f1ccc904a52a18e0389cb0c391339f4;
assign I6d4d8c9c5618d829ae0018df43f15d076f1ccc904a52a18e0389cb0c391339f4 = 
        y_nr_in[2] ^ 
        y_nr_in[48] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[28] = 
I6d4d8c9c5618d829ae0018df43f15d076f1ccc904a52a18e0389cb0c391339f4 ^ 
0; 



wire If296e9a72fef3ff98620606579b8af07856534777912ea92151d42f5be64b05d;
assign If296e9a72fef3ff98620606579b8af07856534777912ea92151d42f5be64b05d = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[27] = 
If296e9a72fef3ff98620606579b8af07856534777912ea92151d42f5be64b05d ^ 
0; 



wire I2af0bb5df1f0fe84b17e106c385543bd55c85e0365549990d04b33ab5f2e74fa;
assign I2af0bb5df1f0fe84b17e106c385543bd55c85e0365549990d04b33ab5f2e74fa = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[26] = 
I2af0bb5df1f0fe84b17e106c385543bd55c85e0365549990d04b33ab5f2e74fa ^ 
0; 



wire If632a83f77b0aa7549d123643fc2b4427d6391a72d838648dd03ab31352372f7;
assign If632a83f77b0aa7549d123643fc2b4427d6391a72d838648dd03ab31352372f7 = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[25] = 
If632a83f77b0aa7549d123643fc2b4427d6391a72d838648dd03ab31352372f7 ^ 
0; 



wire Ic8e0c1fab86c3fc2efbb461160d3db91df504461718a14701bb9c652661dadb6;
assign Ic8e0c1fab86c3fc2efbb461160d3db91df504461718a14701bb9c652661dadb6 = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[24] = 
Ic8e0c1fab86c3fc2efbb461160d3db91df504461718a14701bb9c652661dadb6 ^ 
0; 



wire Ib81aef819af7eaf50fdf170905ca5699723c458df23e7791d858966abe44da49;
assign Ib81aef819af7eaf50fdf170905ca5699723c458df23e7791d858966abe44da49 = 
        y_nr_in[0] ^ 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[23] = 
Ib81aef819af7eaf50fdf170905ca5699723c458df23e7791d858966abe44da49 ^ 
0; 



wire I704ac7d61669664b7f7a796f7e26155ae1f0f656a6de81d61aee29d14d302530;
assign I704ac7d61669664b7f7a796f7e26155ae1f0f656a6de81d61aee29d14d302530 = 
        y_nr_in[1] ^ 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[22] = 
I704ac7d61669664b7f7a796f7e26155ae1f0f656a6de81d61aee29d14d302530 ^ 
0; 



wire I9a3445c2c9c2e42f2041be87b3ea46e08a118a9d0d4dc6ebdd4ecc52c9d1cd15;
assign I9a3445c2c9c2e42f2041be87b3ea46e08a118a9d0d4dc6ebdd4ecc52c9d1cd15 = 
        y_nr_in[2] ^ 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[21] = 
I9a3445c2c9c2e42f2041be87b3ea46e08a118a9d0d4dc6ebdd4ecc52c9d1cd15 ^ 
0; 



wire I0827304f2332549c6da2e80ccf1fb5b7152bbfd2559afb0c5661d1298d90c659;
assign I0827304f2332549c6da2e80ccf1fb5b7152bbfd2559afb0c5661d1298d90c659 = 
        y_nr_in[3] ^ 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[20] = 
I0827304f2332549c6da2e80ccf1fb5b7152bbfd2559afb0c5661d1298d90c659 ^ 
0; 



wire I1f00da6ff425eed3e09c4bcfbbd7206baa0d744f27af21472d92d8bb292652bd;
assign I1f00da6ff425eed3e09c4bcfbbd7206baa0d744f27af21472d92d8bb292652bd = 
        y_nr_in[43] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[19] = 
I1f00da6ff425eed3e09c4bcfbbd7206baa0d744f27af21472d92d8bb292652bd ^ 
0; 



wire I0df5d59942ede8b6716c5c1d1818ed78f644a9071ce61109329bba43196318c1;
assign I0df5d59942ede8b6716c5c1d1818ed78f644a9071ce61109329bba43196318c1 = 
        y_nr_in[40] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[18] = 
I0df5d59942ede8b6716c5c1d1818ed78f644a9071ce61109329bba43196318c1 ^ 
0; 



wire I2d6be792841b5ee8a0774f54b95c77d16dd543bbe64f369c5b73d00e02a9e8ae;
assign I2d6be792841b5ee8a0774f54b95c77d16dd543bbe64f369c5b73d00e02a9e8ae = 
        y_nr_in[41] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[17] = 
I2d6be792841b5ee8a0774f54b95c77d16dd543bbe64f369c5b73d00e02a9e8ae ^ 
0; 



wire I51d939f878a58409a1ba113e3fef13e230ac7eca1814081d2b7c14fd7a4f0575;
assign I51d939f878a58409a1ba113e3fef13e230ac7eca1814081d2b7c14fd7a4f0575 = 
        y_nr_in[42] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[16] = 
I51d939f878a58409a1ba113e3fef13e230ac7eca1814081d2b7c14fd7a4f0575 ^ 
0; 



wire I8fe902ebd1fe8196d8f0e4d2a4d5c1b3232a2fa885024af241456ba02452ed41;
assign I8fe902ebd1fe8196d8f0e4d2a4d5c1b3232a2fa885024af241456ba02452ed41 = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[15] = 
I8fe902ebd1fe8196d8f0e4d2a4d5c1b3232a2fa885024af241456ba02452ed41 ^ 
0; 



wire I12ead1c5b4ad7a80282c7bf8a596b0b874da021e7dbdc0c5cf4318605b1f4db4;
assign I12ead1c5b4ad7a80282c7bf8a596b0b874da021e7dbdc0c5cf4318605b1f4db4 = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[14] = 
I12ead1c5b4ad7a80282c7bf8a596b0b874da021e7dbdc0c5cf4318605b1f4db4 ^ 
0; 



wire Ib49c30590196e02a7627c6582e18ce798c9c5205d2bd338d6fb162bbbd6ced82;
assign Ib49c30590196e02a7627c6582e18ce798c9c5205d2bd338d6fb162bbbd6ced82 = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[13] = 
Ib49c30590196e02a7627c6582e18ce798c9c5205d2bd338d6fb162bbbd6ced82 ^ 
0; 



wire I57294caecb5f3beed2193a3f9df63ffc1cf9943931d8493c19a8849dcbb8d3ef;
assign I57294caecb5f3beed2193a3f9df63ffc1cf9943931d8493c19a8849dcbb8d3ef = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[12] = 
I57294caecb5f3beed2193a3f9df63ffc1cf9943931d8493c19a8849dcbb8d3ef ^ 
0; 



wire I030aa23d83088b82f22244b4588a36ed10b1a6c67f1d278051f29bcebc358885;
assign I030aa23d83088b82f22244b4588a36ed10b1a6c67f1d278051f29bcebc358885 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[50] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[11] = 
I030aa23d83088b82f22244b4588a36ed10b1a6c67f1d278051f29bcebc358885 ^ 
0; 



wire I29f0260d83cd38f848de2e7ddbba4c28f003876cd1402cb2bedc9023cc3c78c4;
assign I29f0260d83cd38f848de2e7ddbba4c28f003876cd1402cb2bedc9023cc3c78c4 = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[51] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[10] = 
I29f0260d83cd38f848de2e7ddbba4c28f003876cd1402cb2bedc9023cc3c78c4 ^ 
0; 



wire I2132db60c0aa88eb27c8f004fdc471842f15122d18f4728df4322d5cdf565cdf;
assign I2132db60c0aa88eb27c8f004fdc471842f15122d18f4728df4322d5cdf565cdf = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[48] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[9] = 
I2132db60c0aa88eb27c8f004fdc471842f15122d18f4728df4322d5cdf565cdf ^ 
0; 



wire I1c007b005b9db6f68d869da323b7fda21f96c28446dffc2d43bda384042d8fc0;
assign I1c007b005b9db6f68d869da323b7fda21f96c28446dffc2d43bda384042d8fc0 = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[49] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[8] = 
I1c007b005b9db6f68d869da323b7fda21f96c28446dffc2d43bda384042d8fc0 ^ 
0; 



wire I5064f9ddff05e6df2591376d7d36499f80ea9f3e6be549d3ff52e99926a104c8;
assign I5064f9ddff05e6df2591376d7d36499f80ea9f3e6be549d3ff52e99926a104c8 = 
        y_nr_in[8] ^ 
        y_nr_in[43] ^ 
        y_nr_in[52] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[7] = 
I5064f9ddff05e6df2591376d7d36499f80ea9f3e6be549d3ff52e99926a104c8 ^ 
0; 



wire I87d977cdaf15f668b4205036e35be9f3c094da82f872551fd042574e219935cf;
assign I87d977cdaf15f668b4205036e35be9f3c094da82f872551fd042574e219935cf = 
        y_nr_in[9] ^ 
        y_nr_in[40] ^ 
        y_nr_in[53] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[6] = 
I87d977cdaf15f668b4205036e35be9f3c094da82f872551fd042574e219935cf ^ 
0; 



wire I4872eb6611eb72183b37df081976136b3c325f0cf01310feb4222628d7a1a105;
assign I4872eb6611eb72183b37df081976136b3c325f0cf01310feb4222628d7a1a105 = 
        y_nr_in[10] ^ 
        y_nr_in[41] ^ 
        y_nr_in[54] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[5] = 
I4872eb6611eb72183b37df081976136b3c325f0cf01310feb4222628d7a1a105 ^ 
0; 



wire Iccb824da507f3919bbf9fa2151dd363418877ac39d3ac57ebf5e596c23c312cf;
assign Iccb824da507f3919bbf9fa2151dd363418877ac39d3ac57ebf5e596c23c312cf = 
        y_nr_in[11] ^ 
        y_nr_in[42] ^ 
        y_nr_in[55] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[4] = 
Iccb824da507f3919bbf9fa2151dd363418877ac39d3ac57ebf5e596c23c312cf ^ 
0; 



wire Ia85f346fc9e3916dc0d6e486afa6f894d5125cca2984ed13de23f15b49ef26cd;
assign Ia85f346fc9e3916dc0d6e486afa6f894d5125cca2984ed13de23f15b49ef26cd = 
        y_nr_in[5] ^ 
        y_nr_in[21] ^ 
        y_nr_in[46] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[3] = 
Ia85f346fc9e3916dc0d6e486afa6f894d5125cca2984ed13de23f15b49ef26cd ^ 
0; 



wire I4b47082e58bc2efdc953ce47fd2f7e16b0e870dc6383ba90fd9f63cae7662a13;
assign I4b47082e58bc2efdc953ce47fd2f7e16b0e870dc6383ba90fd9f63cae7662a13 = 
        y_nr_in[6] ^ 
        y_nr_in[22] ^ 
        y_nr_in[47] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[2] = 
I4b47082e58bc2efdc953ce47fd2f7e16b0e870dc6383ba90fd9f63cae7662a13 ^ 
0; 



wire Icb4bb04fef3700255ae2029f363c33248ebe78dc94d53d303566a1e95a7d979c;
assign Icb4bb04fef3700255ae2029f363c33248ebe78dc94d53d303566a1e95a7d979c = 
        y_nr_in[7] ^ 
        y_nr_in[23] ^ 
        y_nr_in[44] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[1] = 
Icb4bb04fef3700255ae2029f363c33248ebe78dc94d53d303566a1e95a7d979c ^ 
0; 



wire If33d792729453c4e26ebc593398f9aa1b963b20b0cb22467be03a3c0e369a93d;
assign If33d792729453c4e26ebc593398f9aa1b963b20b0cb22467be03a3c0e369a93d = 
        y_nr_in[4] ^ 
        y_nr_in[20] ^ 
        y_nr_in[45] ^ 
0; 



assign Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c[0] = 
If33d792729453c4e26ebc593398f9aa1b963b20b0cb22467be03a3c0e369a93d ^ 
0; 



assign y_nr[m_int-1:0    ] = Ie92cd4bf91559fa3b7ff7e09054c786f5ead3b2e5930dda92caf0d4060cd714c [m_int-1       : 0          ]; //I65966f0faeeff2d783a9e9766d96bafb9ce7ea133ccabd263106f6d7ff1ddd14 Idec0f004eaa07c2a283ea326df8f00c2c3c60b002c9bb8d452b1dcff5ba795cb:m_int I8c6fb1e9e37a1aea1d308c785192e1a17d71cef08c7f50a68d2e0ab292b2e7f4 I83e01dda3eb5a450a0a4d3498dab1d7bc0b9e892edf23936a71188f7b595d815
assign y_nr[n_int-1:m_int] = y_nr_in[n_int-m_int-1 : 0          ]; //message Idec0f004eaa07c2a283ea326df8f00c2c3c60b002c9bb8d452b1dcff5ba795cb:n_int-m_int Iaee610558292023758a4229ddcf75f167c9904313a83cf795232ed7f7e2131c9 I83e01dda3eb5a450a0a4d3498dab1d7bc0b9e892edf23936a71188f7b595d815
