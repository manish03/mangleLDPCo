reg [flogtanh_WDTH -1:0] I51db5b688feb51ec24e6127d4c3dfdae, I869ad51812ced1ce31815a7ccaf5578d;
reg [flogtanh_WDTH -1:0] Ibc891c78cf9dbf2365d9c88acc400657, I6442979212fb9e03df3685a28065f02e;
reg [flogtanh_WDTH -1:0] I690dfdbfc7e73591927914aeb8cb121a, I5e2d92b7f01402ec98771a9026c756e5;
reg [flogtanh_WDTH -1:0] I531efe3d41d7bc16091c3c247cebaaf0, I3050b73b4bf3bb60e38178a3a372231f;
reg [flogtanh_WDTH -1:0] Icf7b3d66021580efed4e68c38d44ac48, I32f1d36a7d8d44da0bc6d3ad8d2a1153;
reg [flogtanh_WDTH -1:0] I93d13a86c9d185bf2c3cf5c34eeeb016, I7637d7cc7dc2189e17cce002a981082a;
reg [flogtanh_WDTH -1:0] I3ded617611b49004853f17e60013d498, I0cb1cf10cb15dd8c1066f460f67538c2;
reg [flogtanh_WDTH -1:0] Ia2414bf52998b14337d78da6aeaec255, Ifbe06c2706fb89aaa251789703159e25;
reg [flogtanh_WDTH -1:0] Ieac60a94c2a709b738af1f3465a59240, I8fe4558357f35c3e71ab801b22392c83;
reg [flogtanh_WDTH -1:0] I88349c865dbc4ddba373b69215a50400, Ic6a2f31a403a6389f0d7df052a5cfdec;
reg [flogtanh_WDTH -1:0] I72adcb5f4bd99318abd40c3b63287f93, I96b2c098a97cd3303228da6f6484e240;
reg [flogtanh_WDTH -1:0] I6cda0f5db099dbb900cd3d0a8f6dc245, I9d07ffc430043e95f348f4d05d3f6dbb;
reg [flogtanh_WDTH -1:0] I4b7867a55677b1a9264c6d1c3eac25e4, I4cd469fecb0f25820f04091a44c50b61;
reg [flogtanh_WDTH -1:0] I09a6bc8c6f42aa92f4b08511d5cd98b8, Ib7fe035c4d2cc2f25edc04489db7a532;
reg [flogtanh_WDTH -1:0] Ia64c991ab9c3fc3488a835de4fdb60b1, I923a9ae3ead074bc3abd711b3378060d;
reg [flogtanh_WDTH -1:0] I94cfcd3eeef047bb244a722337080b4d, I53c4fe7b76ec5282e86c2fb100bb6b18;
reg [flogtanh_WDTH -1:0] Ibebed3263875106ae630c0656211ee39, Ib1f88a9e7696e0798fbeedbbd1aaaf92;
reg [flogtanh_WDTH -1:0] I0439fd68942b4d70cdad2d56ee4b954c, Iabe16f9be9c25cd6e4c2b63984a7e09b;
reg [flogtanh_WDTH -1:0] If4c337b9bbfc2530377ac6db8f13014c, I606e85239115132c5e6281b7ed7ec81a;
reg [flogtanh_WDTH -1:0] I9b705704a3308d69156c7343fa4eb777, I4bddbe88c41a009f869df437614dfd3f;
reg [flogtanh_WDTH -1:0] I5849744db9fdcad905885f296a170c02, I5f13934441008d491b64e006c2704a7f;
reg [flogtanh_WDTH -1:0] I7cdf69d491d37935cef6eca36eb3fe81, I95fac6d42827444b8f030a140cf1ea13;
reg [flogtanh_WDTH -1:0] Idde15d5b821d09d8a406e09d1e4bda88, I33399cd8c4a4774d52f0ff4940f8321e;
reg [flogtanh_WDTH -1:0] I944a0b47e85dab69de22e950ba042e2a, I2abe8717ff4ddfa416d7b2cb47edf15d;
reg I5a0cb346d513664787453b72c079d980 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I869ad51812ced1ce31815a7ccaf5578d <= 'h0;
 I6442979212fb9e03df3685a28065f02e <= 'h0;
 I5e2d92b7f01402ec98771a9026c756e5 <= 'h0;
 I3050b73b4bf3bb60e38178a3a372231f <= 'h0;
 I32f1d36a7d8d44da0bc6d3ad8d2a1153 <= 'h0;
 I7637d7cc7dc2189e17cce002a981082a <= 'h0;
 I0cb1cf10cb15dd8c1066f460f67538c2 <= 'h0;
 Ifbe06c2706fb89aaa251789703159e25 <= 'h0;
 I8fe4558357f35c3e71ab801b22392c83 <= 'h0;
 Ic6a2f31a403a6389f0d7df052a5cfdec <= 'h0;
 I96b2c098a97cd3303228da6f6484e240 <= 'h0;
 I9d07ffc430043e95f348f4d05d3f6dbb <= 'h0;
 I4cd469fecb0f25820f04091a44c50b61 <= 'h0;
 Ib7fe035c4d2cc2f25edc04489db7a532 <= 'h0;
 I923a9ae3ead074bc3abd711b3378060d <= 'h0;
 I53c4fe7b76ec5282e86c2fb100bb6b18 <= 'h0;
 Ib1f88a9e7696e0798fbeedbbd1aaaf92 <= 'h0;
 Iabe16f9be9c25cd6e4c2b63984a7e09b <= 'h0;
 I606e85239115132c5e6281b7ed7ec81a <= 'h0;
 I4bddbe88c41a009f869df437614dfd3f <= 'h0;
 I5f13934441008d491b64e006c2704a7f <= 'h0;
 I95fac6d42827444b8f030a140cf1ea13 <= 'h0;
 I33399cd8c4a4774d52f0ff4940f8321e <= 'h0;
 I2abe8717ff4ddfa416d7b2cb47edf15d <= 'h0;
 I5a0cb346d513664787453b72c079d980 <= 'h0;
end
else
begin
 I869ad51812ced1ce31815a7ccaf5578d <=  I51db5b688feb51ec24e6127d4c3dfdae;
 I6442979212fb9e03df3685a28065f02e <=  Ibc891c78cf9dbf2365d9c88acc400657;
 I5e2d92b7f01402ec98771a9026c756e5 <=  I690dfdbfc7e73591927914aeb8cb121a;
 I3050b73b4bf3bb60e38178a3a372231f <=  I531efe3d41d7bc16091c3c247cebaaf0;
 I32f1d36a7d8d44da0bc6d3ad8d2a1153 <=  Icf7b3d66021580efed4e68c38d44ac48;
 I7637d7cc7dc2189e17cce002a981082a <=  I93d13a86c9d185bf2c3cf5c34eeeb016;
 I0cb1cf10cb15dd8c1066f460f67538c2 <=  I3ded617611b49004853f17e60013d498;
 Ifbe06c2706fb89aaa251789703159e25 <=  Ia2414bf52998b14337d78da6aeaec255;
 I8fe4558357f35c3e71ab801b22392c83 <=  Ieac60a94c2a709b738af1f3465a59240;
 Ic6a2f31a403a6389f0d7df052a5cfdec <=  I88349c865dbc4ddba373b69215a50400;
 I96b2c098a97cd3303228da6f6484e240 <=  I72adcb5f4bd99318abd40c3b63287f93;
 I9d07ffc430043e95f348f4d05d3f6dbb <=  I6cda0f5db099dbb900cd3d0a8f6dc245;
 I4cd469fecb0f25820f04091a44c50b61 <=  I4b7867a55677b1a9264c6d1c3eac25e4;
 Ib7fe035c4d2cc2f25edc04489db7a532 <=  I09a6bc8c6f42aa92f4b08511d5cd98b8;
 I923a9ae3ead074bc3abd711b3378060d <=  Ia64c991ab9c3fc3488a835de4fdb60b1;
 I53c4fe7b76ec5282e86c2fb100bb6b18 <=  I94cfcd3eeef047bb244a722337080b4d;
 Ib1f88a9e7696e0798fbeedbbd1aaaf92 <=  Ibebed3263875106ae630c0656211ee39;
 Iabe16f9be9c25cd6e4c2b63984a7e09b <=  I0439fd68942b4d70cdad2d56ee4b954c;
 I606e85239115132c5e6281b7ed7ec81a <=  If4c337b9bbfc2530377ac6db8f13014c;
 I4bddbe88c41a009f869df437614dfd3f <=  I9b705704a3308d69156c7343fa4eb777;
 I5f13934441008d491b64e006c2704a7f <=  I5849744db9fdcad905885f296a170c02;
 I95fac6d42827444b8f030a140cf1ea13 <=  I7cdf69d491d37935cef6eca36eb3fe81;
 I33399cd8c4a4774d52f0ff4940f8321e <=  Idde15d5b821d09d8a406e09d1e4bda88;
 I2abe8717ff4ddfa416d7b2cb47edf15d <=  I944a0b47e85dab69de22e950ba042e2a;
 I5a0cb346d513664787453b72c079d980 <=  Id11ca9ab1b4b30c21f7314a04c9c7fae;
end
