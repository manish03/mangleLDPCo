 reg  ['h3:0] [$clog2('h7000+1)-1:0] Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470 ;
