              I3f25e297b4ae3ff6c54ea0761a7741ab = 
          (!fgallag_sel[8]) ? 
                       I3d32661f72eecdf4328276db451f7f39: 
                       I5a79ce433bace8f19e5a49a5f0046bf1;
               I40768e536b89956ee6a20a300cf36fd7 =  0;
