reg [flogtanh_WDTH -1:0] flogtanh0x00005_0, flogtanh0x00005_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_1, flogtanh0x00005_1_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_2, flogtanh0x00005_2_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_3, flogtanh0x00005_3_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_4, flogtanh0x00005_4_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_5, flogtanh0x00005_5_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_6, flogtanh0x00005_6_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_7, flogtanh0x00005_7_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_8, flogtanh0x00005_8_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_9, flogtanh0x00005_9_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_10, flogtanh0x00005_10_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00005_11, flogtanh0x00005_11_q;
reg start_d_flogtanh0x00005_q ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 flogtanh0x00005_0_q <= 'h0;
 flogtanh0x00005_1_q <= 'h0;
 flogtanh0x00005_2_q <= 'h0;
 flogtanh0x00005_3_q <= 'h0;
 flogtanh0x00005_4_q <= 'h0;
 flogtanh0x00005_5_q <= 'h0;
 flogtanh0x00005_6_q <= 'h0;
 flogtanh0x00005_7_q <= 'h0;
 flogtanh0x00005_8_q <= 'h0;
 flogtanh0x00005_9_q <= 'h0;
 flogtanh0x00005_10_q <= 'h0;
 flogtanh0x00005_11_q <= 'h0;
 start_d_flogtanh0x00005_q <= 'h0;
end
else
begin
 flogtanh0x00005_0_q <=  flogtanh0x00005_0;
 flogtanh0x00005_1_q <=  flogtanh0x00005_1;
 flogtanh0x00005_2_q <=  flogtanh0x00005_2;
 flogtanh0x00005_3_q <=  flogtanh0x00005_3;
 flogtanh0x00005_4_q <=  flogtanh0x00005_4;
 flogtanh0x00005_5_q <=  flogtanh0x00005_5;
 flogtanh0x00005_6_q <=  flogtanh0x00005_6;
 flogtanh0x00005_7_q <=  flogtanh0x00005_7;
 flogtanh0x00005_8_q <=  flogtanh0x00005_8;
 flogtanh0x00005_9_q <=  flogtanh0x00005_9;
 flogtanh0x00005_10_q <=  flogtanh0x00005_10;
 flogtanh0x00005_11_q <=  flogtanh0x00005_11;
 start_d_flogtanh0x00005_q <=  start_d_flogtanh0x00004_q;
end
