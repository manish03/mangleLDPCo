              I84ab01f2ac31304c9525b8983d34300d = 
          (!fgallag_sel[1]) ? 
                       Ia6f93d7eab83c88b604f8a81a74c04e9: 
                       Ice05aa8a4d2a062da9785286081fd024;
              Iaf7ae8cb478fce9deaf537c13fa083cb = 
          (!fgallag_sel[1]) ? 
                       I6e41efdbe6eeb41b9c9b39e56f3d8b9c: 
                       Ibe53a3b8a9caa8643361263d463290c8;
              Idce9e18b46f498af68bbb108da7441bc = 
          (!fgallag_sel[1]) ? 
                       Ifbcddebb5f791d2df0b2e7aa94a81c22: 
                       I341146b894d9d94c2c803e6b6c464085;
              Ie3954c25e29ea2d7e1340a59d3d7165f = 
          (!fgallag_sel[1]) ? 
                       Iccfcaba2f6129c8201cb97323a8e740a: 
                       I850f7b404a1ab022498350d9ef0cbdc2;
              Iaa12f10c6588df5d8d8444c61b422c7c = 
          (!fgallag_sel[1]) ? 
                       Ie88f3ca2bc79208be9385225a7ad7268: 
                       If4137d66b193970e9ae89b8e1b00e8ca;
              I9851178cd4e84140f2c244f19c285e4a = 
          (!fgallag_sel[1]) ? 
                       I877047b00cef1f6a938ed9915215e203: 
                       Ic9e529e5e428a666bf6bcf2041969d1e;
              I463cc1b85874882aadc9fa0ed9eb7816 = 
          (!fgallag_sel[1]) ? 
                       I2e8ce46a773bcf5f2c3129441a267af4: 
                       Ie734c46bfea46055c73a2642b3f8a7da;
              I5249c4136a601a94d06d4955be304799 = 
          (!fgallag_sel[1]) ? 
                       Id980a518f6b9c84062f5bd7d6f57472f: 
                       I8901003e5fb9f89fddb0fa87dc5b2d05;
              I9ce88b0e18af39ed6dc46db59a2bb78b = 
          (!fgallag_sel[1]) ? 
                       Ia5402393b456807ca5fee0ecb219c7d9: 
                       I41d38680c5aca0364ef9c716cd4525e7;
              I3695c8773a6d76c02a9f8849ada96902 = 
          (!fgallag_sel[1]) ? 
                       I03ee8c787b49b08c0a5a503bd28fcca5: 
                       Id85bac587e9c200406f0aecafbaf3dd5;
              I4783f15f954421f7538cf39210bb44d5 = 
          (!fgallag_sel[1]) ? 
                       Ibb5dbc2fc80aca18dbaa13b7ecdb6c20: 
                       I9b5df9c23c9a2aaa14a99abd110075cb;
              Ia82244e3d80e219740368bab411242be = 
          (!fgallag_sel[1]) ? 
                       Ic00f5a4dfdbbf58316107417ccc6bb74: 
                       Ic208118fb71fea311016edcb1203407d;
              Ib42df9a31ffd2cfc4a63cf95cf89c4d7 = 
          (!fgallag_sel[1]) ? 
                       Ib3d96f215fc42ace8fddda8c64afbc05: 
                       Ie304d02670ae74fb93fb42328d43079e;
              I752d56e6caa726064dc20d4eeda763a9 = 
          (!fgallag_sel[1]) ? 
                       I1a875fdb7e3681839eeb5fdb8c6b47c3: 
                       I85c6964245f5e3423ddfcae7ae864429;
              Ie339fd09fbad7893452b9a2f92d45932 = 
          (!fgallag_sel[1]) ? 
                       Idd3396a16fde9c928bfd71f9b05b98bf: 
                       I3a124ec3bd01d433c39ecbfd0b153d74;
              Ifd15d58d88de80f2cfc98c7f66f8f88d = 
          (!fgallag_sel[1]) ? 
                       I7be57c1f60b38d43d0fe2c02175aeef5: 
                       I886a56b1cae34e1860e4cd2c28606a45;
              I994cd956aabc31d730d77d9b67bbc1db = 
          (!fgallag_sel[1]) ? 
                       I4dfc6b1e7b358ad6a32f6682e487d962: 
                       I4c60daf9c53a50f2a228ca9ad0d75115;
              Ie7086ba45d27b8fd48ad4dbbc1a6466b = 
          (!fgallag_sel[1]) ? 
                       I5fa487af5385cb6dcd0bac274a2b2261: 
                       If3024e217350078f9a06275cc31b6699;
              I8539ebc561f7f4d823623b1f11255213 = 
          (!fgallag_sel[1]) ? 
                       Ifb39ced2cc4424e46be38af68161181a: 
                       I17934cad1385024244ce8bd07b709db0;
              Iedbd35fd7ebaf3787a08b0551ffb324e = 
          (!fgallag_sel[1]) ? 
                       Ie43b90c9bb7dcb76f116c75615df246b: 
                       I7f095ecd42b65b1781e2290db664a73d;
              I23df575a91b34e0a642bf679a74a747c = 
          (!fgallag_sel[1]) ? 
                       I4d7c79dc1c72745d5750cac86454beb8: 
                       I00c66baa19546590a542100f8883d4ab;
              Icce0e60e3e31993ef47683a80567b1c4 = 
          (!fgallag_sel[1]) ? 
                       I97293ec9139e6e252c554d9f26619f06: 
                       I067a46089f564be32860d44b3c69af1a;
              I172b401633d8844fcabdd4b980f46c73 = 
          (!fgallag_sel[1]) ? 
                       Ib11764f9c254c7ddf0782d0cccae0067: 
                       Ic63385ac292f30c59ab2ad6f8b7d8903;
              I71ed80b7d77c2a35edcefe9ce7db28af = 
          (!fgallag_sel[1]) ? 
                       I5d3f02e43c3a9ab32c9769c1cf45ec6c: 
                       I968edb5f5a70a3d391db21db00dafe78;
              Ib1873b0070c00bfe5ed6fda941cfe95e = 
          (!fgallag_sel[1]) ? 
                       I59ad05479adc69422b7e06e4507a8f7a: 
                       I3755b61b6fb958538b1b906a4ad1103d;
              I6db83f8bbff7cde9c9db248c02fd9358 = 
          (!fgallag_sel[1]) ? 
                       I0ba5990e179758e1080a8407412a9a59: 
                       I7562a62ae85c4676605b60594722a950;
              If65d96ffe364426e1b90303ad323e7fb = 
          (!fgallag_sel[1]) ? 
                       I62c2ba2ded74107adfcbe43670718e65: 
                       Ie43871350b062263474a7e0dbca850ce;
              I8e6c7979ddefa5e27581107ca2495e3e = 
          (!fgallag_sel[1]) ? 
                       I12d1f6ac4ef39cb76907b09745b4f8ad: 
                       If9b05209071a1c16ecce1c28f886ee1d;
              I161c2f4e7657ff863ec2a319ee8d21d5 = 
          (!fgallag_sel[1]) ? 
                       Iebb87060282934e67cd1e7e8493fcf20: 
                       I22b235f6e6f0938fe2a026f91bfd72cf;
              Ic18bc04d9a02bccce383f311102a8b45 = 
          (!fgallag_sel[1]) ? 
                       I185299c78eca06f6174996089a2df4d5: 
                       I90f70f8385f7d8fc69fe21f42d96eeeb;
              I8a118ced20140ec0f90f1f82161bd2c1 = 
          (!fgallag_sel[1]) ? 
                       I5d03a9d2e8ca426a10005cf5a1689f4f: 
                       I1f30e3cf906aa5a09d71f23c5be461ba;
              I2b73e4b6134a9ca11b301452734741a1 = 
          (!fgallag_sel[1]) ? 
                       I13069dca0bc85e00a513e9fe7562b346: 
                       Ib69a5ff88f694a3cf18fa11fcccdd9c2;
              Ie432836bf5a95e8dbb6de2c29d9ab058 = 
          (!fgallag_sel[1]) ? 
                       If4b3a419df7ce8b8cd5f2b7a26e1a629: 
                       I03b2bc96c0edf4f4c27ab02d8beda293;
               I8a777efecfec25782e29fd4e8f270490 =  Iddd38c69253e1ba79f6762c9e69857ad ;
               I3ad4e40b398385b2c3a94cabd4736926 =  I0bb76633859552dc99f63b3c520037cc ;
               Ifcd756c806de58265e16199e27f64e22 =  Ia43aac10d65d1661b3d7f9968c829c21 ;
              Icac3b989b3d04d9c7a80d5eebcbb2027 = 
          (!fgallag_sel[1]) ? 
                       Ic9b31062ba9aedcda0f4c91e39fe1814: 
                       Ie5ff9375515964757ffe821812ed8e73;
              I806f4137adef04fa14f4c159fd47bb46 = 
          (!fgallag_sel[1]) ? 
                       I5152ee18b04c8d038ead4817bc68fa57: 
                       I606544d89b457531a204f0a9a061dc74;
              I6f6db1dfb50f19379683f16c549624b3 = 
          (!fgallag_sel[1]) ? 
                       If7bcb8673722495218ae395b5716c89a: 
                       I755d5c8837cace07fc3c0393a6ba2a43;
               Ib26efe2924ee3c384a8f8b0f7f63e0f4 =  I2051dc0ec4b2e1de6e3308c6e0ae74bd ;
              I0a45d8f9e12c5234855b972d39246589 = 
          (!fgallag_sel[1]) ? 
                       Id017562a43e853ec27712b3f8d449361: 
                       I7c408398d6b1e91c00962636fbf59b83;
              I7a9fe30fbe486c1fd6d92b334f04a97b = 
          (!fgallag_sel[1]) ? 
                       I53387cf352304840ccae53d5b5b153e7: 
                       I6d483d27683d84d2309d756d36f43ae9;
               Ia5bc1b93ee0908ca26a967bc4720e5c3 =  I1c44630f8f2d9bf2a5df81f22a67ed43 ;
              I6cd39d0d0d14283cd00870fa8697cbe2 = 
          (!fgallag_sel[1]) ? 
                       I591e5713ec07915309f4a588ea51a990: 
                       Ibab6e2a97bd19438998b97780bdae17d;
               Id33e3cde2a62f32d114a78300c2fdc1b =  Icb868f4e4f276036478f3977e8d831a3 ;
              I22f6c61d2512a383ecc57e2dac6e346a = 
          (!fgallag_sel[1]) ? 
                       I44049fcab453cba240bed48d89a664e5: 
                       I4c6d3af7a2d1adb1f60b61a523dd9bff;
               I00b3081cd7dd077a53bdd7781b98fe6c =  I70d83e5081cd2c9051f9c6b8652462d7 ;
               Ibdf94fc4ee66c4af146968bf34ae4c0c =  Ib9318ad9f3aa8b5fd8b8c59fe3bd1616 ;
               Idadb48591ec328a331bdcf45e9156485 =  Id399e2be28090c81e93743f1bfe00347 ;
               I6315c142854dc3c1893bcb08b46bc739 =  I23d474402240b1761c2f9d785cd2973b ;
              I362b966433fe2df6176a09951d0d88db = 
          (!fgallag_sel[1]) ? 
                       I116f8968c4a02e2a22a8ea4eb5dd3951: 
                       I1ebdf4675d0986c912c52af538ac358d;
               If210d0b145e2fd9cb2e1229c2c9c7a36 =  I92cd919b7b5b4ca8984668bfbdb43d3b ;
               Ia133b750fb093f377556735adb4e3097 =  Ie79b340519a003c4388b90a3d8fac445 ;
              I6d2fcf19c79a538ec57aff56b8579def = 
          (!fgallag_sel[1]) ? 
                       Id2a6a7580c31d450f8c78217e8997f7e: 
                       I74f0171925c0986fe140602b09a0caf2;
               If507c9ebcb1bc24a59ab4a00fc902d88 =  I5e9bef3789fd851fb793bea78beef829 ;
               I70be43895e7446395ee6f209431a4b0e =  I238a8e826a1d8f069455ae0163d508f2 ;
               Iec863324907434f27365ce30e0a3a636 =  Ib8a70644d197140114eacd4c9612dd77 ;
              Ifdd6e035d37dc6a726502ea875e19bf2 = 
          (!fgallag_sel[1]) ? 
                       I80d67b47c44a3b424d1ed4c8e357c265: 
                       Iaa9183f11cd736e6271b9e6259a807a7;
               I0bac49aa5c179287d028c0bbe2f26646 =  I1f2ac0b753cee68f5e984de8994f2f0d ;
               I676f1d8111d39181de6fb867fcc8aad9 =  I4c8185fc93a069b6fa81b3936de2b4b0 ;
               Ib6003647304cdf7e04f112ea1434d0c2 =  I8f8316a85f64267a15f99a0b47db5f08 ;
               I32f1ca64465d5ffd4c0abef6a0713795 =  I713819fe0cf6d54393d9cd5a32a37807 ;
               Iab2dbd174b3566d2eb0c32118a1d6ffc =  I8a99662ff2d2b8f153d6d9359b88eff5 ;
              I119a639a5c5243e5bbf6224fea9e0542 = 
          (!fgallag_sel[1]) ? 
                       I972077c6595b44e3113b0d7a925aa913: 
                       Idde043a5721004c3904eb2b55031e7c1;
               I51a744f6026f58a3ff9d47f7ad8441c7 =  Iebfd00d9a2a6e39e6fc73f95c4f29539 ;
               Ied88a6d77466adfacecc91792e092022 =  I62895b1265f950882fc5fb770dafd51d ;
               I531565b08841415ba9f98966030529f2 =  Icd6b85be80234c06eaeaf1347ebabb38 ;
               I35641e3719c76fbc8621771af415d10f =  Iea7a223f22fb02e29871f500b61fa205 ;
               I56baf72a394546e751edf096f5a87970 =  Ic767ff5ab4bfc377cf1b7bae10b42d3e ;
               I07ab92c9ad141c03101d587f00202c81 =  I41d92f30c38301789ac4155986c2a634 ;
               I0143dfa3c201c85bdcce5739dee11814 =  I1bf648fa37015e2997a689769881149c ;
              Ie9a0ea695884198a9fd7e5de0a9f73d0 = 
          (!fgallag_sel[1]) ? 
                       I74c408ce157c47049698b52949d1fd38: 
                       I3ed597f1774bf9274566cb5fc7dbbdc5;
               I0a066ff1810c068d1807dd5999880170 =  I8d111345e29debfc7addbb913d4e9054 ;
               I3d390c1d2a5df6decbc45bd682760b84 =  I68521e797f1f404e6a190855b1a322f1 ;
               I0b1c32f0732334693986eea6aaee2b12 =  I2adb86feb263103c1419d34eb9b8ae4e ;
               Ifb9c5b70184594cb9f7961cb99c0d62e =  I4db74afe0a9f15f643d8295051f762c0 ;
               I105a0656b51423653fd7428001efa81f =  Ifc1dfcb0afd77d1a01bbb54da77a5f70 ;
               Id9515c02ee595dc6ce4353decfbd2928 =  If878a4e87d963261e36cde448d6c3bbc ;
               Ib1d40c92e79f6562475204ba330c15e3 =  I8b553bf742d14f23835e62aeade33413 ;
               Ief1a527fee16c6cb996ca3363d4713d8 =  Ifc3d28213bc38fbcff2eb42ebc350c8a ;
               I5c7ed7d4a522cf1e94035b3475d07240 =  I5c42c7a5b8b8d73e5374eb00cf80f91b ;
               Ie59496301d7ef6565b69072f4530ceee =  I757c6c719d8455faea81fa0901a2c15e ;
               I2d2b69150858f521850b9d71ee17acbf =  I40fd0db59f8b8877f3f62b9b87e2892d ;
               I0556476f50843423945a3783fd5c9612 =  I07acde143b8be8c4ec4e562a66562b58 ;
               I34f9b6d4f00ab598a94274629c08e99c =  I13b47a7b710051dde6ab5cae17f216d4 ;
               I2f16d9a27f31109e57160fbc03a98853 =  Ica09fab419a2bd1a966956988b6507b3 ;
               Ib19a79508dff3510b087cb2c1df176f9 =  I354ec2d3605e41d982076dcb7e32d2c1 ;
               I48ac3afb4f8b31f9aadc59aaf1a28a44 =  I30084765c13a4c6a7514a16e3f45a9c2 ;
               Ia3bbc4519f9cd9651e10efaace317875 =  I7401e0464789f88be2b661eb055bbdef ;
               I51118baae7de42e5f69f1a78d1ceccad =  0;
