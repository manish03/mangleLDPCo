//`include "GF2_LDPC_fgallag_0x0000e_assign_inc.sv"
//always_comb begin
              I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00000] = 
          (!fgallag_sel['h0000e]) ? 
                       Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00000] : //%
                       Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00001] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00001] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00002] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00002] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00004] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00003] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00006] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00004] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00008] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00005] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000a] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00006] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000c] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00007] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000e] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00008] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00010] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00009] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00012] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000a] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00014] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000b] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00016] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000c] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00018] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000d] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001a] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000e] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001c] ;
//end
//always_comb begin // 
               I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000f] =  Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001e] ;
//end
