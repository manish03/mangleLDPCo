              Ib2aa0dad949a7608d49dfdec8811fead = 
          (!flogtanh_sel[2]) ? 
                       Iba870e87f87c875ff098cafadf28d262: 
                       Icca31b5b8e9f944b504a02ba62118cc7;
              Ia6b922271dbe47dd60eb4d0492fd5739 = 
          (!flogtanh_sel[2]) ? 
                       I43afe6aef28fcced58953c4b3a9b3eed: 
                       Ieed89d20b342594d04aa6adca4cf2edf;
              Idf881bd96e29e48e7efacbb467ff7c5c = 
          (!flogtanh_sel[2]) ? 
                       Ibc5eb7267931e83838a653795dc809b1: 
                       Iedd54575ec8e5a76566ae1313faedb7c;
              I20717481aece4914e0f7222ae35d1456 = 
          (!flogtanh_sel[2]) ? 
                       I7b3ee2f269cb1f90235f1af617e5c3d9: 
                       I7935f561c946b80813603b40e7652f91;
              Ifcfb5c6c620ff437f7830d0c6d939e62 = 
          (!flogtanh_sel[2]) ? 
                       I97c22b8b68524a584412c15361d761cc: 
                       I7d2a8ad5ee9f7a3e9d642735a85a9a23;
              I286aa151ea1dba5e7e6c4639e80b8cf2 = 
          (!flogtanh_sel[2]) ? 
                       I07057436f307eac4f43cd5cb9274f963: 
                       I2f4c421ebd4de08c8f660aa125eb06d3;
              Ia14165ce5e9de831dcd289ac0495e42e = 
          (!flogtanh_sel[2]) ? 
                       I760715bc18504dc4ef1f861035f6f8f7: 
                       If4e8fc4e2bbb39e7beb6db11b58d8232;
              Iad283604bd9143b0729e1d7d1f49dfbb = 
          (!flogtanh_sel[2]) ? 
                       I082a57b5a74e7e39bcf5d12acd15e272: 
                       Ief8973860cdc98a7e4cce37573e3acb9;
              If14b995d06822c80d9d714d4bbbcda58 = 
          (!flogtanh_sel[2]) ? 
                       If72bc16b595b4a2f27b2639e2b033e39: 
                       Ibc2aacfd2026e5970b2ae172c703784b;
              Iece268d0f9e7bdda5bcf50208cf24762 = 
          (!flogtanh_sel[2]) ? 
                       I71f0fb5ab1d8d8a20c53435e79081eef: 
                       Ic7937c4ac4365348de1d96ece551555c;
              I087bd6d6037f7ee9e82663387ac0f820 = 
          (!flogtanh_sel[2]) ? 
                       I7f4db8e60704ff9f4b74094d188e0dda: 
                       I34ad34e3ccac9eb915309c29568da011;
              I0c2fb3d39b747d63854302c08ec8b1c2 = 
          (!flogtanh_sel[2]) ? 
                       Ia006bebb09394969493a92514c8713b5: 
                       Ib2fbcacfe3daa5d49e950f5ebabf258f;
              Id3d9536b013c4766333f6d23066ead54 = 
          (!flogtanh_sel[2]) ? 
                       I98e3b2ac676d6e2555f2286631e0c43d: 
                       Iaaf05004e8c7866bb2ec1d46e76cd5a5;
              Ibc1ee835e7e2d5432583440c90304c56 = 
          (!flogtanh_sel[2]) ? 
                       Idbde787e711114043d18cd262802b234: 
                       I061dc14bf9bc7b97d69893ab5b084f00;
              I594ca16757d13f9bd17dae2114615a80 = 
          (!flogtanh_sel[2]) ? 
                       Iaa784a3cc93b4939eb183ccc94bb8089: 
                       Ifb75793136968aa2432e934f9e849695;
              Id7f43a01fda8433c8b72871f35ef7bdc = 
          (!flogtanh_sel[2]) ? 
                       I3f333a2b43e5db6062346394119bfbaf: 
                       I3b0f64d1ae335c61b01f2209bcdc8333;
              Id850fafd66d7cd6901821100a3290a23 = 
          (!flogtanh_sel[2]) ? 
                       Iccd3b8b6b6e2a4d60d81d4f367d971c7: 
                       Iae2e1facdac5fd4726d1a6b77849b2f6;
              I9a0a13f48f3e52b33be36fe03a9f2da3 = 
          (!flogtanh_sel[2]) ? 
                       Iac2dd16556eed4d7f826f2063d8979ff: 
                       I879638f9da54bd5a8a5ff78f7b011739;
              I77ad3e9b4bafb0b2a4e86f453c9c59a0 = 
          (!flogtanh_sel[2]) ? 
                       Ic4958fe74930007506b93064b9f87588: 
                       If1618b6028dfd675842dc0fa24485ddf;
              Ic3b0467ebe638a2bd44437784b22329e = 
          (!flogtanh_sel[2]) ? 
                       If22a928365940b767923b37527ec904f: 
                       I8586e464f05f813699f9d466970085dd;
              Id57e199202dd2b2fd585b7cbde5f2ad3 = 
          (!flogtanh_sel[2]) ? 
                       I3bc0dcbecfbefea5fb1d0b617d0efa78: 
                       I3ba79b98d30ac9111420c21e244bf338;
              I03ea04be646c4834304d4f82d3171243 = 
          (!flogtanh_sel[2]) ? 
                       Id0e2a5919dcda34c1fcd9230d79d402c: 
                       I203eedac26099a1b191c73411c443e3d;
              I8ac44624c0749e8e870c9dde42ffb8dd = 
          (!flogtanh_sel[2]) ? 
                       I31bce9c2121ec3e7de33fd80027cdf38: 
                       I13702c5d75b212144cc0a3f060887b46;
              I7852770263dd0c5503c75135d38058c4 = 
          (!flogtanh_sel[2]) ? 
                       I4e3c3bcf1ca00767b813fec32d679779: 
                       Iaabe6440ad8902891ba43f734d7c2935;
               Icf8a31b29e9f8918802c3bf5baa48fa5 =  I69dc2265888e6ff99b608329353fb5b8 ;
              I94a9a947dc58e38c7c3e13bf1bab6f51 = 
          (!flogtanh_sel[2]) ? 
                       Ic652a50c7dc405a941fe04abc2170434: 
                       Ic9b544f863bc0820276ac101c90d38f0;
              Ic92921fa31c014ee1c49384973b33176 = 
          (!flogtanh_sel[2]) ? 
                       I3d5ba70412e03b55a77463d256016a7f: 
                       I842efe9f673c4d17759b83e4b6e86a4b;
               Iabedd360b191a5862ad534eea51ab52e =  I23dfb343d3762798b72aec1aeb2f4b4d ;
              I4659f7245c85f3db58d6be3f97cb3cf0 = 
          (!flogtanh_sel[2]) ? 
                       I81ccdf38e45a3e285b02ef75c30b997d: 
                       I3bd029d3007a94b52c72423af9f0ae79;
               I164cbb304f4db6a716bd788036086266 =  I675db209cea9deaa18aaa4ace818d238 ;
               I8775c4f7dd528188506d94cc13862f93 =  Ifcd5afdf257eab5b1f6c7906290abdfd ;
              Ibb600c26f9f0972df669d2d04a96c7f6 = 
          (!flogtanh_sel[2]) ? 
                       Ie801d81c4251559ca6661da90df75c79: 
                       Ide9dd8e36e4508731c54d883e4a2e2ee;
               Ied0b82caf207f1992f7ec334a9fb423c =  Iaedb40c3bffbe0928b2b23275b85ddd4 ;
               I235cbb8f044d1ac3bf4f53c932b5a34b =  I7acb86a7e521fad3f1123b86e310b18a ;
               I1d25723c499c68dea49c4d762d80bcc3 =  I86df045ba01e5daeb569d9ea1a3263d7 ;
              I6309f136f930378ab3b8cf5a29cfafdf = 
          (!flogtanh_sel[2]) ? 
                       I0583dbd1d4e65defd1ba2fbe2bd87d0a: 
                       I1a7a8ed99d0d10bcefd5a51600d1ceb6;
               I4d5d1e9c151f5e4e18596916c57b891d =  Ic541d5047749fb2833bfa23bad86e2ae ;
               I134c07a35862ad54f8852c17a8bab5de =  I02cfa4d934a334809afc76213ef6cdff ;
               I5b663cc1d7cc3069f33b63799aa34796 =  I75c142058c4a21b970356e0575e2d025 ;
               Ia2ed52a8130a197b3a198aa454d980b0 =  I561431791c47fa1b7455126752aac55e ;
               I13acb2c915e11641c53157310e44892b =  I5004693a6347e9b31037639942d06504 ;
               I6a5212af01917f8e71e3e83bd9e8caf2 =  I73709d12931c354b73a1369cac5db3a9 ;
               I3fe2af1aa64d019af984fa86c1292ad9 =  I6e3a3dc54544c2601df65e24390247e4 ;
               Ic09f027112d6b05b07873fda8e85bea2 =  Ia7d3383c61357b1b2fa53a9f3728a3da ;
              If35467fdae216528f1dd248b2c19feba = 
          (!flogtanh_sel[2]) ? 
                       I1a296cef71412b570eaa40a564f146e2: 
                       Ib34c55a2554033229a576daae46633f1;
               I6681491d836b3bf63f771b708625f7b6 =  0;
