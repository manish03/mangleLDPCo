 reg  ['h3ff:0] [$clog2('h7000+1)-1:0] I230a233857da8a64905ea1b1de0d2509543fa79c4521eb44f066ab1d16a07322 ;
