 reg  ['h3ffff:0] [$clog2('h7000+1)-1:0] I92c63025ac2cd3f26f34ecb614257096b9bb60b5c9460c2f364ee04b9ed913df ;
