 reg  ['h7ff:0] [$clog2('h7000+1)-1:0] Ia940d1a12f2aecb1cf57d9d7b9e7b4aa ;
