 reg  ['h7:0] [$clog2('h7000+1)-1:0] Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7 ;
